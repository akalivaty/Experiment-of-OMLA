//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n578, new_n579,
    new_n580, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n651,
    new_n654, new_n655, new_n657, new_n658, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT69), .B1(new_n471), .B2(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n466), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n465), .A2(new_n468), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n468), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT70), .ZN(G162));
  OAI211_X1 g063(.A(G138), .B(new_n468), .C1(new_n463), .C2(new_n464), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n483), .A2(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n490), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G62), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n501), .B2(KEYINPUT72), .ZN(new_n505));
  OAI21_X1  g080(.A(G651), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n499), .A2(new_n500), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G88), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n511), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n515), .B1(new_n511), .B2(new_n514), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n506), .B1(new_n517), .B2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n524), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n521), .B(new_n526), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n510), .A2(G51), .B1(new_n512), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n512), .A2(new_n513), .A3(G89), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n521), .B1(new_n537), .B2(new_n526), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT74), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n526), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT73), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n541), .A2(new_n542), .A3(new_n533), .A4(new_n535), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(G168));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI21_X1  g120(.A(G543), .B1(new_n529), .B2(new_n530), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n531), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n528), .A2(new_n527), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G651), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n552), .B2(new_n553), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n548), .B1(new_n554), .B2(new_n556), .ZN(G171));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT76), .B(G43), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n531), .A2(new_n559), .B1(new_n546), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(G56), .B1(new_n528), .B2(new_n527), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n555), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n558), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n499), .B2(new_n500), .ZN(new_n567));
  INV_X1    g142(.A(new_n563), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n512), .A2(new_n513), .A3(G81), .ZN(new_n570));
  INV_X1    g145(.A(new_n560), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(new_n510), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n569), .A2(KEYINPUT77), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  NAND4_X1  g151(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT78), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT8), .ZN(new_n580));
  NAND4_X1  g155(.A1(G319), .A2(G483), .A3(G661), .A4(new_n580), .ZN(G188));
  OAI211_X1 g156(.A(G53), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n550), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n499), .A2(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n586), .A2(G651), .B1(new_n587), .B2(G91), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n583), .A2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  INV_X1    g165(.A(G168), .ZN(G286));
  NAND2_X1  g166(.A1(new_n587), .A2(G87), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n510), .A2(G49), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n596));
  OAI21_X1  g171(.A(G61), .B1(new_n528), .B2(new_n527), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  AOI211_X1 g173(.A(new_n596), .B(new_n555), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G86), .ZN(new_n600));
  INV_X1    g175(.A(G48), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n531), .A2(new_n600), .B1(new_n546), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n597), .A2(new_n598), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(new_n596), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT80), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G61), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n499), .B2(new_n500), .ZN(new_n609));
  INV_X1    g184(.A(new_n598), .ZN(new_n610));
  OAI211_X1 g185(.A(KEYINPUT79), .B(G651), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n587), .A2(G86), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n510), .A2(G48), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n615));
  AOI21_X1  g190(.A(KEYINPUT79), .B1(new_n604), .B2(G651), .ZN(new_n616));
  NOR3_X1   g191(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n607), .A2(new_n617), .ZN(G305));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n619));
  INV_X1    g194(.A(G72), .ZN(new_n620));
  INV_X1    g195(.A(G60), .ZN(new_n621));
  OAI221_X1 g196(.A(new_n619), .B1(new_n620), .B2(new_n507), .C1(new_n550), .C2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n499), .B2(new_n500), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n620), .A2(new_n507), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT81), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n622), .A2(G651), .A3(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G85), .ZN(new_n627));
  INV_X1    g202(.A(G47), .ZN(new_n628));
  OAI22_X1  g203(.A1(new_n531), .A2(new_n627), .B1(new_n546), .B2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(G290));
  XNOR2_X1  g206(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n632));
  INV_X1    g207(.A(G92), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n531), .B2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G66), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n499), .B2(new_n500), .ZN(new_n636));
  NAND2_X1  g211(.A1(G79), .A2(G543), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT83), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n639), .A2(G79), .A3(G543), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(G651), .B1(new_n636), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n643));
  NAND4_X1  g218(.A1(new_n643), .A2(G92), .A3(new_n512), .A4(new_n513), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n510), .A2(G54), .ZN(new_n645));
  NAND4_X1  g220(.A1(new_n634), .A2(new_n642), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G868), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(G171), .B2(new_n647), .ZN(G284));
  OAI21_X1  g224(.A(new_n648), .B1(G171), .B2(new_n647), .ZN(G321));
  NOR2_X1   g225(.A1(G299), .A2(G868), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(G168), .B2(G868), .ZN(G297));
  XNOR2_X1  g227(.A(G297), .B(KEYINPUT84), .ZN(G280));
  INV_X1    g228(.A(new_n646), .ZN(new_n654));
  INV_X1    g229(.A(G559), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n655), .B2(G860), .ZN(G148));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G868), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n575), .B2(G868), .ZN(G323));
  XNOR2_X1  g234(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g235(.A1(new_n472), .A2(new_n469), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT12), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT13), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(G2100), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n483), .A2(G123), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  OAI21_X1  g242(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(G111), .ZN(new_n671));
  AOI22_X1  g246(.A1(new_n668), .A2(new_n669), .B1(new_n671), .B2(G2105), .ZN(new_n672));
  AOI22_X1  g247(.A1(new_n466), .A2(G135), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n674), .A2(G2096), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n664), .A2(G2100), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(G2096), .ZN(new_n677));
  NAND4_X1  g252(.A1(new_n665), .A2(new_n675), .A3(new_n676), .A4(new_n677), .ZN(G156));
  XNOR2_X1  g253(.A(G2427), .B(G2438), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2430), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT15), .B(G2435), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(KEYINPUT14), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1341), .B(G1348), .Z(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G2451), .B(G2454), .Z(new_n689));
  XNOR2_X1  g264(.A(G2443), .B(G2446), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n691), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n692), .A2(G14), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n692), .A2(KEYINPUT88), .A3(G14), .A4(new_n693), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(G401));
  XOR2_X1   g273(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n699));
  XOR2_X1   g274(.A(G2084), .B(G2090), .Z(new_n700));
  XNOR2_X1  g275(.A(G2067), .B(G2678), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(KEYINPUT17), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n699), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G2096), .B(G2100), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT91), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G2072), .B(G2078), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT89), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n702), .B2(new_n699), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n708), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G227));
  XOR2_X1   g288(.A(G1991), .B(G1996), .Z(new_n714));
  XNOR2_X1  g289(.A(G1971), .B(G1976), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT19), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1961), .B(G1966), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  XOR2_X1   g293(.A(G1956), .B(G2474), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(new_n716), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  MUX2_X1   g297(.A(new_n716), .B(new_n721), .S(new_n722), .Z(new_n723));
  NOR2_X1   g298(.A1(new_n720), .A2(new_n716), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT20), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n723), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n727), .B1(new_n723), .B2(new_n726), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n714), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(new_n714), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n732), .A2(new_n733), .A3(new_n728), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(G1981), .B(G1986), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n731), .A2(new_n734), .A3(new_n736), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(G229));
  XNOR2_X1  g316(.A(KEYINPUT30), .B(G28), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  OR2_X1    g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n742), .A2(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n674), .B2(new_n743), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(G33), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n472), .A2(G127), .ZN(new_n749));
  AND2_X1   g324(.A1(G115), .A2(G2104), .ZN(new_n750));
  OAI21_X1  g325(.A(G2105), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n752));
  NAND2_X1  g327(.A1(G103), .A2(G2104), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G2105), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n466), .A2(G139), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n748), .B1(new_n758), .B2(new_n743), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n747), .B1(G2072), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  INV_X1    g336(.A(G16), .ZN(new_n762));
  NOR2_X1   g337(.A1(G171), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G5), .B2(new_n762), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n760), .B1(new_n761), .B2(new_n764), .C1(G2072), .C2(new_n759), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n743), .A2(G32), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n483), .A2(G129), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT100), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n469), .A2(G105), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT26), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n769), .B(new_n771), .C1(G141), .C2(new_n466), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n766), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(G164), .A2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G27), .B2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G2078), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n765), .A2(new_n776), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G286), .A2(new_n762), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT101), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(KEYINPUT101), .B1(G16), .B2(G21), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(G1966), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(G1966), .ZN(new_n791));
  INV_X1    g366(.A(G34), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(KEYINPUT24), .ZN(new_n793));
  AOI21_X1  g368(.A(G29), .B1(new_n792), .B2(KEYINPUT24), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(KEYINPUT99), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(KEYINPUT99), .B2(new_n794), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n480), .B2(new_n743), .ZN(new_n797));
  INV_X1    g372(.A(G2084), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n761), .B2(new_n764), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n784), .A2(new_n790), .A3(new_n791), .A4(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT102), .Z(new_n802));
  NAND2_X1  g377(.A1(G166), .A2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G16), .B2(G22), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(G305), .A2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT32), .B(G1981), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n762), .A2(G6), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n762), .A2(G23), .ZN(new_n812));
  INV_X1    g387(.A(G288), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n762), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT33), .B(G1976), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT96), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n804), .A2(new_n805), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n806), .A2(new_n811), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n809), .B1(new_n807), .B2(new_n810), .ZN(new_n820));
  OR3_X1    g395(.A1(new_n819), .A2(KEYINPUT34), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT34), .B1(new_n819), .B2(new_n820), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n743), .A2(G25), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n466), .A2(G131), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n483), .A2(G119), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT93), .B1(G95), .B2(G2105), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(KEYINPUT93), .A2(G95), .A3(G2105), .ZN(new_n829));
  OAI221_X1 g404(.A(G2104), .B1(G107), .B2(new_n468), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n823), .B1(new_n832), .B2(new_n743), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT35), .B(G1991), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT94), .Z(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n833), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(G16), .A2(G24), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n625), .A2(G651), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n629), .B1(new_n839), .B2(new_n622), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT95), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n838), .B1(new_n841), .B2(G16), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(G1986), .Z(new_n843));
  NAND4_X1  g418(.A1(new_n821), .A2(new_n822), .A3(new_n837), .A4(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT36), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n743), .A2(G35), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G162), .B2(new_n743), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT29), .B(G2090), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n762), .A2(G4), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n654), .B2(new_n762), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G1348), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n575), .A2(new_n762), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n762), .B2(G19), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT97), .B(G1341), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n743), .A2(G26), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT28), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n483), .A2(G128), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n483), .A2(KEYINPUT98), .A3(G128), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n865));
  INV_X1    g440(.A(G116), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n866), .B2(G2105), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n466), .B2(G140), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n859), .B1(new_n869), .B2(G29), .ZN(new_n870));
  INV_X1    g445(.A(G2067), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n854), .A2(new_n855), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n762), .A2(G20), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT23), .Z(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(G299), .B2(G16), .ZN(new_n876));
  INV_X1    g451(.A(G1956), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NOR4_X1   g453(.A1(new_n857), .A2(new_n872), .A3(new_n873), .A4(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n802), .A2(new_n845), .A3(new_n879), .ZN(G311));
  NAND3_X1  g455(.A1(new_n802), .A2(new_n845), .A3(new_n879), .ZN(G150));
  NAND2_X1  g456(.A1(G80), .A2(G543), .ZN(new_n882));
  INV_X1    g457(.A(G67), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n550), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G651), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n512), .A2(new_n513), .A3(G93), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n513), .A2(G55), .A3(G543), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT104), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT104), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(G860), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT37), .Z(new_n892));
  NOR2_X1   g467(.A1(new_n646), .A2(new_n655), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n574), .A2(new_n890), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n561), .A2(new_n564), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(new_n885), .C1(new_n889), .C2(new_n888), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n895), .B(new_n899), .Z(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n901), .A2(KEYINPUT39), .ZN(new_n902));
  INV_X1    g477(.A(G860), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n901), .B2(KEYINPUT39), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n892), .B1(new_n902), .B2(new_n904), .ZN(G145));
  NOR2_X1   g480(.A1(new_n773), .A2(new_n757), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n773), .A2(new_n757), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n466), .A2(G142), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n483), .A2(G130), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n468), .A2(G118), .ZN(new_n911));
  OAI21_X1  g486(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n909), .B(new_n910), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n662), .B(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n907), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n758), .B1(new_n768), .B2(new_n772), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n917), .B2(new_n906), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n869), .A2(new_n496), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n869), .A2(new_n496), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n832), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n922), .ZN(new_n924));
  INV_X1    g499(.A(new_n832), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n916), .A2(new_n918), .A3(new_n923), .A4(new_n926), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n674), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(new_n480), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n480), .ZN(new_n934));
  AOI21_X1  g509(.A(G162), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n934), .ZN(new_n936));
  INV_X1    g511(.A(G162), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n936), .A2(new_n932), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n935), .A2(new_n938), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(new_n928), .A3(new_n929), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g520(.A(new_n899), .B(new_n657), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n654), .B2(G299), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n949));
  INV_X1    g524(.A(G91), .ZN(new_n950));
  OAI22_X1  g525(.A1(new_n949), .A2(new_n555), .B1(new_n950), .B2(new_n531), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT9), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n582), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n954), .A2(KEYINPUT105), .A3(new_n646), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n654), .A2(G299), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n948), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n946), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT105), .B1(new_n954), .B2(new_n646), .ZN(new_n960));
  AND4_X1   g535(.A1(KEYINPUT105), .A2(new_n646), .A3(new_n583), .A4(new_n588), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n948), .A2(new_n955), .A3(KEYINPUT106), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n956), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT41), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n960), .A2(new_n961), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n654), .B2(G299), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n964), .A2(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n958), .B1(new_n968), .B2(new_n946), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  NAND2_X1  g545(.A1(G303), .A2(new_n840), .ZN(new_n971));
  INV_X1    g546(.A(G88), .ZN(new_n972));
  INV_X1    g547(.A(G50), .ZN(new_n973));
  OAI22_X1  g548(.A1(new_n531), .A2(new_n972), .B1(new_n546), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT71), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n516), .ZN(new_n976));
  NAND3_X1  g551(.A1(G290), .A2(new_n976), .A3(new_n506), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n979));
  INV_X1    g554(.A(new_n602), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n606), .A2(new_n980), .A3(KEYINPUT80), .A4(new_n611), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n979), .A2(G288), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G288), .B1(new_n979), .B2(new_n981), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n978), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n813), .B1(new_n607), .B2(new_n617), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n979), .A2(G288), .A3(new_n981), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n985), .A2(new_n986), .B1(new_n977), .B2(new_n971), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n989), .B(new_n958), .C1(new_n968), .C2(new_n946), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n970), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(new_n970), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g567(.A(G868), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n890), .A2(new_n647), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(G295));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n996));
  XNOR2_X1  g571(.A(G295), .B(new_n996), .ZN(G331));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n998));
  NAND2_X1  g573(.A1(G168), .A2(G301), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n539), .A2(new_n543), .A3(G171), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n899), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1000), .ZN(new_n1004));
  AOI21_X1  g579(.A(G171), .B1(new_n539), .B2(new_n543), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n896), .B(new_n898), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n999), .A2(new_n899), .A3(KEYINPUT108), .A4(new_n1000), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1003), .A2(new_n957), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1006), .A2(new_n1001), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1008), .B(new_n988), .C1(new_n968), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1010), .A2(new_n943), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1003), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n962), .A2(new_n963), .A3(new_n967), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n957), .A2(new_n965), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1006), .A2(new_n957), .A3(new_n1001), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n984), .B2(new_n987), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n978), .B1(new_n982), .B2(new_n983), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n985), .A2(new_n986), .A3(new_n977), .A4(new_n971), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(KEYINPUT109), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1011), .A2(KEYINPUT43), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1008), .B1(new_n968), .B2(new_n1009), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1028), .A2(new_n1024), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1010), .A2(new_n943), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n998), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT43), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1025), .A2(new_n1027), .A3(new_n943), .A4(new_n1010), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT44), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT110), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1024), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT43), .B1(new_n1011), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1030), .A2(new_n1040), .A3(new_n1027), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT44), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1027), .B1(new_n1011), .B2(new_n1037), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1030), .A2(new_n1040), .A3(KEYINPUT43), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n998), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1036), .A2(new_n1047), .ZN(G397));
  XOR2_X1   g623(.A(KEYINPUT111), .B(G1384), .Z(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT45), .B1(new_n496), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G125), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n465), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n474), .ZN(new_n1053));
  OAI21_X1  g628(.A(G2105), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT112), .B(G40), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1054), .A2(new_n470), .A3(new_n467), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1050), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1996), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n773), .B(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n869), .B(new_n871), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n832), .A2(new_n836), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n925), .A2(new_n835), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(G290), .B(G1986), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1059), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  INV_X1    g643(.A(G1384), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n496), .A2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1068), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n496), .A2(KEYINPUT115), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1057), .B1(new_n1070), .B2(KEYINPUT50), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n798), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT45), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1057), .B1(new_n1070), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n1069), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1966), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1077), .A2(G168), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G8), .ZN(new_n1085));
  AOI21_X1  g660(.A(G168), .B1(new_n1077), .B2(new_n1083), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT51), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1088), .A3(G8), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT62), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1070), .A2(new_n1057), .ZN(new_n1094));
  INV_X1    g669(.A(G8), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1976), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(G288), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1096), .B(new_n1098), .C1(new_n1097), .C2(G288), .ZN(new_n1099));
  INV_X1    g674(.A(G1981), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n603), .B2(new_n606), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n614), .A2(G1981), .A3(new_n616), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT49), .ZN(new_n1103));
  OR3_X1    g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n1096), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1058), .A2(new_n1069), .A3(new_n496), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(G8), .C1(new_n1097), .C2(G288), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT52), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1099), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G303), .A2(G8), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT55), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1057), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(KEYINPUT50), .B2(new_n1070), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT116), .B(G2090), .Z(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n1049), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n496), .A2(KEYINPUT113), .A3(KEYINPUT45), .A4(new_n1049), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(G1971), .B1(new_n1122), .B2(new_n1079), .ZN(new_n1123));
  OAI21_X1  g698(.A(G8), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1110), .B1(new_n1112), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1075), .A2(new_n1076), .A3(new_n1115), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT117), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1075), .A2(new_n1128), .A3(new_n1076), .A4(new_n1115), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1123), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1112), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(G8), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1122), .A2(new_n780), .A3(new_n1079), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1134), .A2(new_n1135), .B1(new_n1136), .B2(new_n761), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1135), .A2(G2078), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1079), .A2(new_n1080), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(G301), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1125), .A2(new_n1133), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1091), .A2(new_n1093), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1133), .A2(new_n1110), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1106), .A2(new_n1097), .A3(new_n813), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1144), .A2(new_n1102), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1096), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n1095), .B(G286), .C1(new_n1077), .C2(new_n1083), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1133), .A2(KEYINPUT63), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1132), .B1(new_n1131), .B2(G8), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT118), .B1(new_n1149), .B2(new_n1110), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1110), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1123), .B1(KEYINPUT117), .B2(new_n1126), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1095), .B1(new_n1153), .B2(new_n1129), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1151), .B(new_n1152), .C1(new_n1154), .C2(new_n1132), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1148), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1125), .A2(new_n1133), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n1157), .B2(new_n1147), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1142), .B(new_n1146), .C1(new_n1156), .C2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n476), .A2(G40), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n1162), .A2(new_n1050), .A3(KEYINPUT124), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT124), .B1(new_n1162), .B2(new_n1050), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1122), .A3(new_n1138), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1136), .A2(new_n761), .ZN(new_n1166));
  AND4_X1   g741(.A1(G301), .A2(new_n1161), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1160), .B1(new_n1140), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1161), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(G171), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1137), .A2(G301), .A3(new_n1139), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1170), .A2(new_n1171), .A3(KEYINPUT54), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1157), .A2(new_n1168), .A3(new_n1090), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1114), .A2(new_n877), .ZN(new_n1174));
  XNOR2_X1  g749(.A(KEYINPUT56), .B(G2072), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1122), .A2(new_n1079), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n954), .B(KEYINPUT57), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1174), .A2(new_n1178), .A3(new_n1176), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT61), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n646), .A2(KEYINPUT122), .ZN(new_n1183));
  INV_X1    g758(.A(G1348), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1136), .A2(new_n1184), .B1(new_n871), .B2(new_n1094), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1183), .B1(new_n1185), .B2(KEYINPUT60), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(KEYINPUT60), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n646), .A2(KEYINPUT122), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1185), .A2(KEYINPUT60), .A3(new_n1183), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1182), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1122), .A2(new_n1060), .A3(new_n1079), .ZN(new_n1192));
  XOR2_X1   g767(.A(KEYINPUT58), .B(G1341), .Z(new_n1193));
  NAND2_X1  g768(.A1(new_n1107), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT120), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1195), .A2(new_n1196), .A3(new_n575), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1196), .B1(new_n1195), .B2(new_n575), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT59), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1199), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT59), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1201), .A2(new_n1202), .A3(new_n1197), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1181), .A2(KEYINPUT121), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1181), .A2(KEYINPUT121), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1178), .B(KEYINPUT119), .Z(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1177), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1205), .A2(KEYINPUT61), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1191), .A2(new_n1204), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1185), .A2(new_n646), .ZN(new_n1211));
  AOI22_X1  g786(.A1(new_n1211), .A2(new_n1181), .B1(new_n1177), .B2(new_n1207), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1173), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1067), .B1(new_n1159), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1059), .A2(KEYINPUT46), .A3(new_n1060), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT126), .ZN(new_n1216));
  INV_X1    g791(.A(new_n773), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1062), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1216), .B1(new_n1059), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g794(.A(KEYINPUT46), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT125), .Z(new_n1221));
  AND3_X1   g796(.A1(new_n1219), .A2(KEYINPUT47), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g797(.A(KEYINPUT47), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1224));
  OAI22_X1  g799(.A1(new_n1224), .A2(new_n1063), .B1(G2067), .B2(new_n869), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1225), .A2(new_n1059), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1065), .A2(new_n1059), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT48), .ZN(new_n1228));
  NOR2_X1   g803(.A1(G290), .A2(G1986), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1059), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1227), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(new_n1230), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1232), .A2(KEYINPUT48), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1226), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  NOR3_X1   g809(.A1(new_n1222), .A2(new_n1223), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1214), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g811(.A1(new_n712), .A2(new_n461), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1238), .B1(new_n696), .B2(new_n697), .ZN(new_n1239));
  AND3_X1   g813(.A1(new_n944), .A2(new_n740), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g814(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1241));
  NAND2_X1  g815(.A1(new_n1240), .A2(new_n1241), .ZN(G225));
  XNOR2_X1  g816(.A(G225), .B(KEYINPUT127), .ZN(G308));
endmodule


