//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT67), .ZN(new_n211));
  AND2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n210), .A2(new_n211), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT68), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n214), .A2(new_n215), .B1(G77), .B2(G244), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(G116), .A2(G270), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT69), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n208), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G250), .ZN(new_n229));
  NOR2_X1   g0029(.A1(G257), .A2(G264), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n231), .A2(KEYINPUT0), .ZN(new_n232));
  INV_X1    g0032(.A(new_n201), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n235), .A2(G20), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n231), .A2(KEYINPUT0), .ZN(new_n239));
  NAND3_X1  g0039(.A1(new_n232), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  NOR2_X1   g0041(.A1(new_n226), .A2(new_n241), .ZN(G361));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  INV_X1    g0043(.A(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT2), .B(G226), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G250), .B(G257), .Z(new_n248));
  XNOR2_X1  g0048(.A(G264), .B(G270), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G358));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(G68), .B(G77), .Z(new_n255));
  XNOR2_X1  g0055(.A(G50), .B(G58), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n220), .ZN(new_n260));
  OAI21_X1  g0060(.A(G20), .B1(new_n260), .B2(new_n201), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G159), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G20), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT7), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT79), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(KEYINPUT79), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n271), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n269), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(KEYINPUT80), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT80), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n274), .A2(KEYINPUT79), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n283));
  AOI21_X1  g0083(.A(G33), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n284), .B2(new_n278), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n270), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n265), .B1(new_n286), .B2(new_n220), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT16), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n236), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n282), .A2(new_n283), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n274), .A2(new_n271), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(new_n269), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n220), .B1(new_n295), .B2(KEYINPUT7), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT7), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n293), .A2(new_n297), .A3(new_n269), .A4(new_n294), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n264), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n292), .B1(new_n299), .B2(KEYINPUT16), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n259), .A2(KEYINPUT8), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT71), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n259), .A2(KEYINPUT8), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G1), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G20), .ZN(new_n310));
  INV_X1    g0110(.A(G13), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n292), .A2(new_n310), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n289), .A2(new_n300), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n309), .B1(G41), .B2(G45), .ZN(new_n318));
  INV_X1    g0118(.A(G274), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G41), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(G1), .A3(G13), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n318), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G232), .ZN(new_n326));
  INV_X1    g0126(.A(G87), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n271), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G223), .A2(G1698), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n293), .B2(new_n294), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(G226), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n328), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT70), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n323), .A2(KEYINPUT70), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n321), .B(new_n326), .C1(new_n334), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n338), .ZN(new_n342));
  AOI211_X1 g0142(.A(new_n329), .B(new_n332), .C1(new_n293), .C2(new_n294), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(new_n328), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n344), .A2(G179), .A3(new_n321), .A4(new_n326), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n317), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(KEYINPUT18), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n314), .A2(new_n316), .ZN(new_n350));
  INV_X1    g0150(.A(new_n270), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT80), .B1(new_n276), .B2(new_n279), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n284), .A2(new_n281), .A3(new_n278), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G68), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT16), .B1(new_n355), .B2(new_n265), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n295), .A2(KEYINPUT7), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(G68), .A3(new_n298), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n265), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n291), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n350), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n341), .A2(new_n345), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(KEYINPUT18), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT82), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n363), .A2(KEYINPUT81), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n363), .B2(KEYINPUT81), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n349), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT18), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n317), .A2(new_n346), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT81), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT82), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n363), .A2(KEYINPUT81), .A3(new_n364), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n348), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G200), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n340), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G190), .B2(new_n340), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT83), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n375), .B(KEYINPUT83), .C1(G190), .C2(new_n340), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n317), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT17), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n367), .A2(new_n373), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n271), .A2(G20), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n307), .A2(new_n384), .B1(G150), .B2(new_n262), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n203), .A2(G20), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n292), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n202), .B2(new_n312), .ZN(new_n388));
  INV_X1    g0188(.A(new_n315), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G50), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT74), .B1(new_n392), .B2(KEYINPUT9), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n294), .A2(new_n277), .ZN(new_n394));
  NOR2_X1   g0194(.A1(G222), .A2(G1698), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n331), .A2(G223), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n342), .B(new_n397), .C1(G77), .C2(new_n394), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n321), .C1(new_n219), .C2(new_n324), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G200), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n399), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n392), .B2(KEYINPUT9), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT74), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT9), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n391), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n393), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT10), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n402), .B2(KEYINPUT75), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n393), .A2(new_n403), .A3(new_n409), .A4(new_n406), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G169), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n399), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n391), .B(new_n415), .C1(G179), .C2(new_n399), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n383), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT15), .B(G87), .Z(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n384), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT72), .ZN(new_n422));
  INV_X1    g0222(.A(G77), .ZN(new_n423));
  INV_X1    g0223(.A(new_n262), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n302), .A2(new_n304), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n422), .B1(new_n269), .B2(new_n423), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n291), .B1(new_n423), .B2(new_n312), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n315), .A2(new_n423), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT73), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(G232), .A2(G1698), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n331), .A2(G238), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n394), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n342), .B(new_n433), .C1(G107), .C2(new_n394), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n325), .A2(G244), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n321), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n414), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n436), .A2(G179), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n430), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT13), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n219), .A2(new_n331), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n442), .B1(G232), .B2(new_n331), .C1(new_n266), .C2(new_n267), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G97), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n320), .B1(new_n445), .B2(new_n342), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n324), .A2(new_n221), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n441), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n444), .A2(new_n443), .B1(new_n337), .B2(new_n338), .ZN(new_n450));
  NOR4_X1   g0250(.A1(new_n450), .A2(KEYINPUT13), .A3(new_n447), .A4(new_n320), .ZN(new_n451));
  OAI21_X1  g0251(.A(G169), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT14), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n294), .A2(new_n277), .B1(new_n244), .B2(G1698), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n454), .A2(new_n442), .B1(G33), .B2(G97), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n321), .B(new_n448), .C1(new_n339), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT13), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n446), .A2(new_n441), .A3(new_n448), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT14), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(G169), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT77), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n451), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n458), .A2(KEYINPUT77), .ZN(new_n465));
  AOI211_X1 g0265(.A(KEYINPUT76), .B(new_n441), .C1(new_n446), .C2(new_n448), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT76), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n456), .B2(KEYINPUT13), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G179), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT78), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n464), .A2(new_n465), .ZN(new_n472));
  INV_X1    g0272(.A(new_n468), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n449), .A2(new_n467), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n472), .A2(new_n475), .A3(new_n476), .A4(G179), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n462), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n384), .A2(G77), .ZN(new_n479));
  OAI221_X1 g0279(.A(new_n479), .B1(new_n269), .B2(G68), .C1(new_n202), .C2(new_n424), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n291), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT11), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n389), .A2(G68), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n312), .A2(new_n220), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT12), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(G200), .B2(new_n459), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n401), .B2(new_n469), .ZN(new_n490));
  INV_X1    g0290(.A(new_n430), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n436), .A2(new_n401), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n436), .A2(G200), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n488), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n293), .A2(new_n294), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G264), .A3(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT88), .ZN(new_n499));
  AOI21_X1  g0299(.A(G1698), .B1(new_n293), .B2(new_n294), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(G257), .B1(G303), .B2(new_n268), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT88), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n497), .A2(new_n502), .A3(G264), .A4(G1698), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n499), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n342), .ZN(new_n505));
  XNOR2_X1  g0305(.A(KEYINPUT5), .B(G41), .ZN(new_n506));
  INV_X1    g0306(.A(G45), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G1), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n335), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(G274), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n509), .A2(G270), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n414), .B1(new_n505), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT84), .B(G116), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n312), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n309), .A2(G33), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n313), .A2(G116), .A3(new_n292), .A4(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(KEYINPUT84), .A2(G116), .ZN(new_n518));
  NOR2_X1   g0318(.A1(KEYINPUT84), .A2(G116), .ZN(new_n519));
  OAI21_X1  g0319(.A(G20), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n269), .C1(G33), .C2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n291), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n515), .B(new_n517), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n524), .B(new_n525), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT89), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n515), .A4(new_n517), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n513), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT21), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n505), .A2(new_n512), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n470), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n533), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n513), .A2(KEYINPUT21), .A3(new_n533), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n533), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n537), .A2(new_n401), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(G200), .B2(new_n537), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G107), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(KEYINPUT6), .A3(G97), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n522), .A2(new_n546), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n550), .B2(KEYINPUT6), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n286), .B2(new_n546), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n291), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n313), .A2(G97), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n313), .A2(new_n292), .A3(new_n516), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n522), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n554), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n331), .A2(G244), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n561), .A2(new_n562), .B1(new_n229), .B2(new_n331), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n394), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n293), .B2(new_n294), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n521), .B(new_n564), .C1(new_n565), .C2(KEYINPUT4), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(new_n342), .B1(G257), .B2(new_n509), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n511), .A2(new_n506), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n414), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n470), .A3(new_n568), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n560), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(G200), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n555), .B1(new_n553), .B2(new_n291), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n567), .A2(G190), .A3(new_n568), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n559), .A4(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n313), .A2(new_n420), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n497), .A2(new_n269), .A3(G68), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT85), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n384), .A2(new_n581), .A3(G97), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n549), .A2(new_n327), .B1(new_n444), .B2(new_n269), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(new_n581), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n497), .A2(KEYINPUT85), .A3(new_n269), .A4(G68), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n577), .B1(new_n586), .B2(new_n291), .ZN(new_n587));
  INV_X1    g0387(.A(new_n420), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n557), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n589), .B(KEYINPUT86), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G238), .A2(G1698), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n331), .A2(G244), .ZN(new_n593));
  AOI211_X1 g0393(.A(new_n592), .B(new_n593), .C1(new_n293), .C2(new_n294), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n514), .A2(new_n271), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n342), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n323), .B(G250), .C1(G1), .C2(new_n507), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n510), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n414), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n596), .A2(new_n510), .A3(new_n597), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n470), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n591), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n557), .A2(new_n327), .ZN(new_n603));
  AOI211_X1 g0403(.A(new_n577), .B(new_n603), .C1(new_n586), .C2(new_n291), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n598), .A2(G200), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n596), .A2(G190), .A3(new_n510), .A4(new_n597), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n572), .A2(new_n576), .A3(new_n602), .A4(new_n607), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n608), .A2(KEYINPUT87), .ZN(new_n609));
  AOI211_X1 g0409(.A(G20), .B(new_n327), .C1(new_n293), .C2(new_n294), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT22), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT90), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n497), .A2(new_n269), .A3(G87), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT90), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(KEYINPUT22), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n394), .A2(new_n611), .A3(new_n269), .A4(G87), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT24), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT23), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n269), .B2(G107), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n546), .A2(KEYINPUT23), .A3(G20), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n595), .A2(new_n269), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n618), .B1(new_n617), .B2(new_n622), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n291), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n557), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT25), .B1(new_n312), .B2(new_n546), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n312), .A2(KEYINPUT25), .A3(new_n546), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n626), .A2(G107), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n509), .A2(G264), .ZN(new_n631));
  INV_X1    g0431(.A(G294), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n271), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(G250), .A2(G1698), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n293), .B2(new_n294), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n331), .A2(G257), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n568), .B(new_n631), .C1(new_n637), .C2(new_n339), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n374), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(G190), .B2(new_n638), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n625), .A2(new_n630), .A3(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n638), .A2(KEYINPUT91), .A3(G169), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT91), .B1(new_n638), .B2(G169), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n638), .A2(new_n470), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n625), .B2(new_n630), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n608), .A2(KEYINPUT87), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n545), .A2(new_n609), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  NOR4_X1   g0449(.A1(new_n419), .A2(new_n440), .A3(new_n496), .A4(new_n649), .ZN(G372));
  NOR3_X1   g0450(.A1(new_n419), .A2(new_n496), .A3(new_n440), .ZN(new_n651));
  INV_X1    g0451(.A(new_n602), .ZN(new_n652));
  INV_X1    g0452(.A(new_n645), .ZN(new_n653));
  INV_X1    g0453(.A(new_n624), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n292), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n630), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n513), .A2(KEYINPUT21), .A3(new_n533), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT21), .B1(new_n513), .B2(new_n533), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n661), .A3(new_n539), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n641), .A2(new_n608), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n652), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n587), .A2(new_n590), .B1(new_n600), .B2(new_n470), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n605), .A2(new_n606), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n599), .A2(new_n665), .B1(new_n666), .B2(new_n604), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n572), .A2(KEYINPUT92), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT92), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n560), .A2(new_n570), .A3(new_n669), .A4(new_n571), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n602), .A2(new_n607), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n572), .ZN(new_n675));
  XOR2_X1   g0475(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n664), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n651), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n440), .A2(new_n490), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n488), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT17), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n380), .B(new_n683), .ZN(new_n684));
  OAI22_X1  g0484(.A1(new_n682), .A2(new_n684), .B1(new_n348), .B2(new_n369), .ZN(new_n685));
  INV_X1    g0485(.A(new_n413), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n417), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n680), .A2(new_n687), .ZN(G369));
  NOR2_X1   g0488(.A1(new_n311), .A2(G20), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n309), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n656), .B2(new_n657), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n647), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n695), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n658), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n545), .B1(new_n542), .B2(new_n698), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n541), .A2(new_n533), .A3(new_n695), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(KEYINPUT94), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT94), .ZN(new_n705));
  AOI211_X1 g0505(.A(new_n705), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n699), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n695), .B1(new_n661), .B2(new_n539), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n647), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n646), .A2(new_n698), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n711), .ZN(G399));
  NOR2_X1   g0512(.A1(new_n228), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n549), .A2(new_n327), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n234), .B2(new_n714), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n569), .A2(new_n638), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT95), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n470), .A3(new_n537), .A4(new_n598), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n638), .B1(KEYINPUT96), .B2(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n726), .A2(new_n567), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n538), .A3(new_n600), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(KEYINPUT96), .B2(new_n725), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n725), .A2(KEYINPUT96), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n727), .A2(new_n538), .A3(new_n600), .A4(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n724), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n695), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n733), .B(KEYINPUT31), .C1(new_n649), .C2(new_n695), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n733), .A2(KEYINPUT31), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n572), .A2(new_n576), .A3(new_n602), .A4(new_n607), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n625), .A2(new_n630), .A3(new_n640), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n739), .B(new_n740), .C1(new_n541), .C2(new_n646), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT26), .A4(new_n670), .ZN(new_n742));
  INV_X1    g0542(.A(new_n676), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n674), .B2(new_n572), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n745), .A3(new_n602), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n698), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n695), .B1(new_n664), .B2(new_n678), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  MUX2_X1   g0549(.A(new_n747), .B(new_n748), .S(new_n749), .Z(new_n750));
  NOR2_X1   g0550(.A1(new_n738), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n720), .B1(new_n751), .B2(G1), .ZN(G364));
  AOI21_X1  g0552(.A(new_n309), .B1(new_n689), .B2(G45), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n714), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n470), .A2(new_n374), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n269), .A2(G190), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n758), .A2(KEYINPUT99), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(KEYINPUT99), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n757), .A2(G179), .A3(new_n374), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n762), .A2(new_n220), .B1(new_n767), .B2(new_n423), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n757), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G159), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n269), .A2(new_n401), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n374), .A2(G179), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G87), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n776), .A2(new_n757), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n268), .B1(new_n781), .B2(G107), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n775), .A2(G179), .A3(new_n374), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n775), .A2(new_n756), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n783), .A2(new_n259), .B1(new_n784), .B2(new_n202), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n269), .B1(new_n769), .B2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n785), .B1(G97), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n774), .A2(new_n779), .A3(new_n782), .A4(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  NOR2_X1   g0590(.A1(new_n762), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n767), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n783), .A2(new_n794), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n791), .A2(new_n793), .A3(new_n394), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n787), .A2(G294), .ZN(new_n797));
  INV_X1    g0597(.A(new_n784), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G326), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G283), .A2(new_n781), .B1(new_n771), .B2(G329), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n796), .A2(new_n797), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G303), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n777), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n789), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n236), .B1(G20), .B2(new_n414), .ZN(new_n805));
  NOR3_X1   g0605(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n805), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n228), .A2(new_n497), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n235), .A2(new_n507), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n810), .B(new_n811), .C1(new_n507), .C2(new_n257), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n228), .A2(new_n268), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G355), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(G116), .C2(new_n227), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n804), .A2(new_n805), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n701), .A2(new_n702), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n755), .B(new_n816), .C1(new_n817), .C2(new_n807), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(G330), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n705), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n703), .A2(KEYINPUT94), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(G330), .C2(new_n817), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n818), .B1(new_n822), .B2(new_n755), .ZN(G396));
  NAND2_X1  g0623(.A1(new_n440), .A2(KEYINPUT102), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT102), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n439), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n827), .B(new_n495), .C1(new_n491), .C2(new_n698), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G13), .A2(G33), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n440), .A2(new_n695), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT100), .B(G283), .Z(new_n832));
  AOI22_X1  g0632(.A1(new_n761), .A2(new_n832), .B1(G97), .B2(new_n787), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n780), .A2(new_n327), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n784), .A2(new_n802), .B1(new_n770), .B2(new_n792), .ZN(new_n835));
  INV_X1    g0635(.A(new_n783), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n834), .B(new_n835), .C1(G294), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n514), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n766), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n394), .B1(new_n778), .B2(G107), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n833), .A2(new_n837), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n761), .A2(G150), .B1(new_n766), .B2(G159), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n784), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G143), .B2(new_n836), .ZN(new_n845));
  XNOR2_X1  g0645(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n780), .A2(new_n220), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G50), .B2(new_n778), .ZN(new_n849));
  INV_X1    g0649(.A(new_n497), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G132), .B2(new_n771), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n847), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n786), .A2(new_n259), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n841), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n805), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n805), .A2(new_n829), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n423), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n831), .A2(new_n755), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT104), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n737), .B(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n494), .B1(new_n824), .B2(new_n826), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n541), .A2(new_n646), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n572), .A2(new_n576), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n740), .A3(new_n667), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n602), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n671), .A2(new_n672), .B1(new_n675), .B2(new_n676), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n698), .B(new_n861), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT103), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n679), .A2(KEYINPUT103), .A3(new_n698), .A4(new_n861), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n828), .A2(new_n830), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n748), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n860), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n754), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n859), .B2(new_n737), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n858), .B1(new_n875), .B2(new_n876), .ZN(G384));
  OAI211_X1 g0677(.A(G20), .B(new_n237), .C1(new_n551), .C2(KEYINPUT35), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n715), .B(new_n878), .C1(KEYINPUT35), .C2(new_n551), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  OAI21_X1  g0680(.A(G77), .B1(new_n259), .B2(new_n220), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n234), .A2(new_n881), .B1(G50), .B2(new_n220), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(G1), .A3(new_n311), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n299), .A2(KEYINPUT16), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n350), .B1(new_n360), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n693), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n382), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n885), .B1(new_n362), .B2(new_n886), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n380), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  INV_X1    g0691(.A(new_n347), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n361), .A2(new_n886), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n892), .A2(new_n380), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n894), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n348), .A2(new_n369), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n899), .B1(new_n684), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n892), .A2(new_n380), .A3(new_n894), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n895), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT39), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n888), .B2(new_n897), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n906), .B(new_n896), .C1(new_n382), .C2(new_n887), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(KEYINPUT39), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n488), .A2(new_n695), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n900), .A2(new_n693), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n827), .A2(new_n695), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n871), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n486), .B2(new_n695), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n486), .A2(new_n919), .A3(new_n695), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n490), .B(new_n921), .C1(new_n478), .C2(new_n487), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n920), .A2(new_n922), .B1(new_n488), .B2(new_n698), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n918), .B(new_n923), .C1(new_n910), .C2(new_n909), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n914), .A2(new_n915), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n750), .A2(new_n651), .A3(KEYINPUT106), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT106), .B1(new_n750), .B2(new_n651), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n687), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n925), .B(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n734), .A2(new_n872), .A3(new_n735), .A4(new_n923), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n901), .B2(new_n904), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n896), .B1(new_n382), .B2(new_n887), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(KEYINPUT38), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT40), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(KEYINPUT107), .A2(KEYINPUT40), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n930), .A2(new_n935), .B1(new_n910), .B2(new_n909), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT107), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n934), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(G330), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n651), .A2(new_n736), .A3(G330), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n651), .A3(new_n736), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n929), .A2(new_n944), .B1(new_n309), .B2(new_n689), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT108), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n929), .A2(new_n944), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n880), .B(new_n883), .C1(new_n946), .C2(new_n947), .ZN(G367));
  AOI21_X1  g0748(.A(KEYINPUT46), .B1(new_n778), .B2(new_n838), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n780), .A2(new_n522), .B1(new_n786), .B2(new_n546), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n949), .A2(new_n497), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G317), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n951), .B1(new_n952), .B2(new_n770), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n761), .A2(G294), .B1(G303), .B2(new_n836), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(new_n792), .C2(new_n784), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n953), .B(new_n956), .C1(new_n766), .C2(new_n832), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n777), .A2(new_n259), .B1(new_n770), .B2(new_n843), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT113), .Z(new_n959));
  INV_X1    g0759(.A(G159), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n959), .B1(new_n202), .B2(new_n767), .C1(new_n960), .C2(new_n762), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n780), .A2(new_n423), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n268), .B1(new_n798), .B2(G143), .ZN(new_n963));
  INV_X1    g0763(.A(G150), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n963), .B1(new_n220), .B2(new_n786), .C1(new_n964), .C2(new_n783), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n961), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n957), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT47), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n805), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n604), .A2(new_n698), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n674), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n652), .A2(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n808), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n810), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n809), .B1(new_n227), .B2(new_n588), .C1(new_n974), .C2(new_n250), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n969), .A2(new_n755), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n753), .B(KEYINPUT111), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n751), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n820), .A2(new_n821), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(KEYINPUT110), .A3(new_n699), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT110), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n707), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT109), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n560), .A2(new_n695), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n863), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n572), .B2(new_n698), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n984), .B(KEYINPUT44), .C1(new_n711), .C2(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n984), .A2(KEYINPUT44), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n984), .A2(KEYINPUT44), .ZN(new_n990));
  OR4_X1    g0790(.A1(new_n711), .A2(new_n989), .A3(new_n987), .A4(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n709), .A2(new_n710), .A3(new_n987), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n981), .A2(new_n983), .A3(new_n988), .A4(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n988), .A3(new_n994), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(new_n982), .A3(new_n707), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n709), .B1(new_n699), .B2(new_n708), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n980), .B(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n979), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n713), .B(KEYINPUT41), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n978), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT112), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n709), .A2(new_n986), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT42), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n572), .B1(new_n986), .B2(new_n658), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n698), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n971), .A2(new_n972), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1008), .A2(new_n1010), .B1(KEYINPUT43), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n980), .A2(new_n699), .A3(new_n987), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1005), .A2(new_n1006), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1006), .B1(new_n1005), .B2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n976), .B1(new_n1017), .B2(new_n1018), .ZN(G387));
  NAND2_X1  g0819(.A1(new_n1001), .A2(new_n977), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1001), .A2(new_n751), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n713), .B1(new_n1001), .B2(new_n751), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n761), .A2(G311), .B1(new_n766), .B2(G303), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n952), .B2(new_n783), .C1(new_n794), .C2(new_n784), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT48), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n632), .B2(new_n777), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n787), .B2(new_n832), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT49), .Z(new_n1028));
  NAND2_X1  g0828(.A1(new_n771), .A2(G326), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n497), .B1(new_n838), .B2(new_n781), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n767), .A2(new_n220), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n770), .A2(new_n964), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n777), .A2(new_n423), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n783), .A2(new_n202), .B1(new_n780), .B2(new_n522), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n308), .B2(new_n762), .C1(new_n588), .C2(new_n786), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n497), .B1(new_n960), .B2(new_n784), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1031), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT114), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n805), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n247), .A2(new_n507), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1042), .A2(new_n810), .B1(new_n716), .B2(new_n813), .ZN(new_n1043));
  AOI21_X1  g0843(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n425), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n202), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n717), .B(new_n1044), .C1(new_n1046), .C2(KEYINPUT50), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT50), .B2(new_n1046), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1043), .A2(new_n1048), .B1(G107), .B2(new_n227), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n809), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1041), .A2(new_n755), .A3(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n699), .A2(new_n807), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .C1(new_n1051), .C2(new_n1052), .ZN(G393));
  OR2_X1    g0853(.A1(new_n1021), .A2(new_n999), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1021), .A2(new_n999), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n713), .A3(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n987), .A2(new_n807), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n783), .A2(new_n960), .B1(new_n784), .B2(new_n964), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT51), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n786), .A2(new_n423), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n850), .A2(new_n834), .A3(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n761), .A2(G50), .B1(new_n766), .B2(new_n1045), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1059), .B(new_n1061), .C1(new_n1062), .C2(KEYINPUT115), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n220), .B2(new_n777), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(G143), .C2(new_n771), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n394), .B1(new_n778), .B2(new_n832), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n836), .A2(G311), .B1(new_n798), .B2(G317), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1067), .B1(new_n546), .B2(new_n780), .C1(new_n1068), .C2(KEYINPUT52), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n761), .A2(G303), .B1(new_n838), .B2(new_n787), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(KEYINPUT52), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n794), .C2(new_n770), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1069), .B(new_n1072), .C1(G294), .C2(new_n766), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n805), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n809), .B1(new_n522), .B2(new_n227), .C1(new_n974), .C2(new_n254), .ZN(new_n1075));
  AND4_X1   g0875(.A1(new_n755), .A2(new_n1057), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n999), .B2(new_n977), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1056), .A2(new_n1077), .ZN(G390));
  INV_X1    g0878(.A(KEYINPUT116), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n734), .A2(new_n872), .A3(new_n735), .A4(G330), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n478), .A2(new_n487), .A3(new_n698), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n922), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n920), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n908), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n888), .A2(new_n897), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n906), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n913), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n916), .B1(new_n869), .B2(new_n870), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n1084), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n746), .A2(new_n698), .A3(new_n861), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1084), .B1(new_n1095), .B2(new_n917), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n933), .A2(new_n1096), .A3(new_n913), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1079), .B(new_n1085), .C1(new_n1094), .C2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1079), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1100));
  AOI211_X1 g0900(.A(KEYINPUT116), .B(new_n1097), .C1(new_n1090), .C2(new_n1093), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1099), .B1(new_n1102), .B2(new_n1085), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1103), .A2(new_n978), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n798), .A2(G283), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n767), .B2(new_n522), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n848), .B(new_n1106), .C1(G294), .C2(new_n771), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n761), .A2(G107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n394), .B(new_n1060), .C1(G87), .C2(new_n778), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n836), .A2(G116), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT117), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n767), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n762), .A2(new_n843), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n964), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n786), .A2(new_n960), .ZN(new_n1117));
  INV_X1    g0917(.A(G132), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n783), .A2(new_n1118), .B1(new_n780), .B2(new_n202), .ZN(new_n1119));
  NOR4_X1   g0919(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n268), .B1(new_n798), .B2(G128), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n771), .A2(G125), .ZN(new_n1122));
  OAI21_X1  g0922(.A(KEYINPUT53), .B1(new_n777), .B2(new_n964), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1111), .B1(new_n1114), .B2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT118), .Z(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n805), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n829), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n755), .B(new_n1127), .C1(new_n912), .C2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n308), .B2(new_n856), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1104), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n687), .B(new_n941), .C1(new_n926), .C2(new_n927), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1085), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1134), .A2(new_n917), .A3(new_n1095), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1135), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n918), .B1(new_n1137), .B2(new_n1085), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n913), .B1(new_n918), .B2(new_n923), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1098), .B1(new_n1141), .B2(new_n912), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT116), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1094), .A2(new_n1079), .A3(new_n1098), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n1085), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1100), .A2(new_n1134), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1140), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(new_n714), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1103), .A2(new_n1140), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1131), .A2(new_n1150), .ZN(G378));
  NAND2_X1  g0951(.A1(new_n391), .A2(new_n886), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n418), .B(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n939), .A2(new_n1156), .A3(G330), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n939), .B2(G330), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n925), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n940), .A2(new_n1155), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n925), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n939), .A2(new_n1156), .A3(G330), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1147), .B2(new_n1132), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n714), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1164), .B(KEYINPUT57), .C1(new_n1147), .C2(new_n1132), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT120), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1133), .B1(new_n1103), .B2(new_n1140), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1171), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n1164), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1167), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(G41), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n293), .A2(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n762), .A2(new_n522), .B1(new_n220), .B2(new_n786), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n420), .C2(new_n766), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1034), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n781), .A2(G58), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n771), .A2(G283), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1178), .A2(new_n294), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G107), .B2(new_n836), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1177), .B(new_n1182), .C1(new_n715), .C2(new_n784), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1183), .A2(new_n1184), .B1(new_n202), .B2(new_n1175), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT119), .Z(new_n1186));
  OAI22_X1  g0986(.A1(new_n1113), .A2(new_n777), .B1(new_n964), .B2(new_n786), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G137), .B2(new_n766), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n798), .A2(G125), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n761), .A2(G132), .B1(G128), .B2(new_n836), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n781), .A2(G159), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G41), .B1(new_n771), .B2(G124), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1192), .A2(new_n271), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1183), .A2(new_n1184), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n805), .B1(new_n1186), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1155), .A2(new_n829), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n856), .A2(new_n202), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1199), .A2(new_n755), .A3(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1164), .A2(new_n977), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1173), .A2(new_n1202), .ZN(G375));
  NAND3_X1  g1003(.A1(new_n1132), .A2(new_n1138), .A3(new_n1136), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1140), .A2(new_n1003), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1084), .A2(new_n829), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n766), .A2(G107), .B1(G294), .B2(new_n798), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n761), .A2(new_n838), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n394), .B1(new_n836), .B2(G283), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n771), .A2(G303), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n588), .A2(new_n786), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n777), .A2(new_n522), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1211), .A2(new_n962), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n762), .A2(new_n1113), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n766), .A2(G150), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n784), .A2(new_n1118), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT121), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n787), .A2(G50), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G159), .A2(new_n778), .B1(new_n781), .B2(G58), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1216), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n771), .A2(G128), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n497), .B1(new_n843), .B2(new_n783), .C1(new_n1217), .C2(KEYINPUT121), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1215), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n805), .B1(new_n1214), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n856), .A2(new_n220), .ZN(new_n1226));
  AND4_X1   g1026(.A1(new_n755), .A2(new_n1206), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1139), .B2(new_n977), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1205), .A2(new_n1228), .ZN(G381));
  AND2_X1   g1029(.A1(new_n1131), .A2(new_n1150), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1173), .A2(new_n1230), .A3(new_n1202), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1231), .A2(G384), .A3(G387), .A4(G381), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(G393), .A2(G390), .A3(G396), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(G407));
  OAI211_X1 g1034(.A(G407), .B(G213), .C1(G343), .C2(new_n1231), .ZN(G409));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1204), .A2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1132), .A2(KEYINPUT60), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1237), .A2(new_n713), .A3(new_n1140), .A4(new_n1238), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1239), .A2(G384), .A3(new_n1228), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G384), .B1(new_n1239), .B2(new_n1228), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(G213), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(G343), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(G2897), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT124), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(KEYINPUT123), .A2(G2897), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(KEYINPUT123), .A2(G2897), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1249), .A2(new_n1245), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1247), .B1(new_n1242), .B2(new_n1252), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1240), .A2(new_n1241), .A3(KEYINPUT124), .A4(new_n1251), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1230), .B1(new_n1173), .B2(new_n1202), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1202), .B1(new_n1165), .B2(new_n1004), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(G378), .A2(new_n1257), .B1(new_n1244), .B2(G343), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1246), .B(new_n1255), .C1(new_n1256), .C2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1256), .A2(new_n1258), .A3(new_n1243), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT63), .B1(new_n1262), .B2(KEYINPUT122), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G375), .A2(G378), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1258), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(new_n1242), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT122), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(G393), .B(G396), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G390), .ZN(new_n1272));
  AND2_X1   g1072(.A1(G387), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n976), .B(G390), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1271), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT125), .ZN(new_n1277));
  AND3_X1   g1077(.A1(G387), .A2(new_n1277), .A3(new_n1272), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(G387), .B2(new_n1272), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1270), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT126), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1274), .B(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1276), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1261), .A2(new_n1263), .A3(new_n1269), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1258), .B1(G375), .B2(G378), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1287), .B2(new_n1242), .ZN(new_n1288));
  NOR4_X1   g1088(.A1(new_n1256), .A2(new_n1258), .A3(KEYINPUT62), .A4(new_n1243), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1285), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1284), .B1(new_n1290), .B2(new_n1283), .ZN(G405));
  NAND2_X1  g1091(.A1(new_n1242), .A2(KEYINPUT127), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1283), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1276), .B(new_n1292), .C1(new_n1280), .C2(new_n1282), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OR2_X1    g1096(.A1(new_n1242), .A2(KEYINPUT127), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1264), .A2(new_n1231), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1298), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1294), .A2(new_n1300), .A3(new_n1295), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(G402));
endmodule


