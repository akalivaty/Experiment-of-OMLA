//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n443, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT65), .B(G108), .ZN(new_n443));
  INV_X1    g018(.A(new_n443), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G235), .A2(G238), .A3(G237), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(new_n458), .B2(G567), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n462), .A2(G137), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G101), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT68), .B1(new_n466), .B2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(new_n463), .A3(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n463), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n462), .A2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n472), .A2(new_n474), .A3(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(G124), .B2(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n463), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n462), .A2(G126), .A3(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n472), .A2(new_n474), .A3(G138), .A4(new_n463), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n462), .A2(new_n503), .A3(G138), .A4(new_n463), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n496), .A2(KEYINPUT70), .A3(new_n497), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n500), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT71), .A3(G62), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(new_n512), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n514), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(G88), .B1(G50), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n521), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT72), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n531), .B(new_n533), .C1(new_n534), .C2(new_n523), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(G51), .B2(new_n526), .ZN(G168));
  AOI22_X1  g111(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n523), .A2(new_n540), .B1(new_n525), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n517), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT73), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n524), .A2(G81), .B1(G43), .B2(new_n526), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n526), .A2(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n523), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n517), .B(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n559), .A2(new_n562), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  OAI21_X1  g145(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n526), .A2(G49), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT77), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n561), .A2(new_n574), .A3(G87), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n574), .B1(new_n561), .B2(G87), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n571), .B(new_n573), .C1(new_n575), .C2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n561), .A2(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n517), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(G48), .A2(new_n526), .B1(new_n581), .B2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n538), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n523), .A2(new_n586), .B1(new_n525), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n561), .A2(G92), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n564), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n561), .A2(new_n598), .A3(G92), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n593), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G168), .B2(new_n604), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(G168), .B2(new_n604), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n601), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n467), .A2(new_n469), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n462), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n486), .A2(G123), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n621));
  INV_X1    g196(.A(G135), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n621), .C1(new_n622), .C2(new_n483), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT15), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2435), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XOR2_X1   g205(.A(G2443), .B(G2446), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G1341), .B(G1348), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G14), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(G401));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT78), .Z(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(KEYINPUT17), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n645), .C1(new_n641), .C2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n642), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n648), .A2(new_n640), .A3(new_n644), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n641), .A2(new_n646), .A3(new_n644), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n647), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2096), .B(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT80), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n656), .A2(new_n657), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT79), .B(KEYINPUT20), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n659), .A2(new_n661), .A3(new_n664), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  INV_X1    g247(.A(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1986), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n671), .B(new_n675), .Z(G229));
  NOR2_X1   g251(.A1(G16), .A2(G23), .ZN(new_n677));
  INV_X1    g252(.A(G288), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(G16), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT33), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G166), .B2(new_n682), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(G1971), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(G6), .ZN(new_n686));
  INV_X1    g261(.A(G305), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n682), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n681), .A2(new_n685), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT81), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT34), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n462), .A2(new_n463), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G131), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n486), .A2(G119), .ZN(new_n696));
  OR2_X1    g271(.A1(G95), .A2(G2105), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  MUX2_X1   g274(.A(G25), .B(new_n699), .S(G29), .Z(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT35), .B(G1991), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n682), .A2(G24), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n589), .B2(new_n682), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1986), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n693), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT82), .B(KEYINPUT36), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n694), .A2(G141), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n486), .A2(G129), .B1(new_n614), .B2(G105), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G32), .B(new_n715), .S(G29), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT27), .B(G1996), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n708), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n693), .A2(new_n719), .A3(new_n706), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G27), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G164), .B2(new_n721), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT91), .B(G2078), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n726));
  NAND2_X1  g301(.A1(G168), .A2(G16), .ZN(new_n727));
  OR2_X1    g302(.A1(G16), .A2(G21), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n726), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1966), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n721), .A2(G33), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(new_n463), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n694), .A2(KEYINPUT83), .A3(G139), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT83), .ZN(new_n736));
  INV_X1    g311(.A(G139), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n483), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT25), .Z(new_n740));
  NAND3_X1  g315(.A1(new_n735), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT84), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(KEYINPUT84), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n734), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n732), .B1(new_n744), .B2(new_n721), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n725), .B(new_n731), .C1(G2072), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI22_X1  g325(.A1(G160), .A2(G29), .B1(KEYINPUT85), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(KEYINPUT85), .B2(new_n750), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT86), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G2084), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT87), .Z(new_n755));
  INV_X1    g330(.A(KEYINPUT28), .ZN(new_n756));
  INV_X1    g331(.A(G26), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G29), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n486), .A2(G128), .ZN(new_n760));
  INV_X1    g335(.A(G140), .ZN(new_n761));
  OAI21_X1  g336(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n463), .A2(G116), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n760), .B1(new_n761), .B2(new_n483), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n758), .B1(new_n765), .B2(new_n756), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT30), .B(G28), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n766), .A2(G2067), .B1(new_n721), .B2(new_n767), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n768), .B1(G2067), .B2(new_n766), .C1(new_n753), .C2(G2084), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n755), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G5), .B2(G16), .ZN(new_n772));
  OR3_X1    g347(.A1(new_n771), .A2(G5), .A3(G16), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n772), .B(new_n773), .C1(G301), .C2(new_n682), .ZN(new_n774));
  INV_X1    g349(.A(G1961), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n746), .A2(new_n770), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT31), .B(G11), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G35), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G162), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2090), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n601), .A2(new_n682), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G4), .B2(new_n682), .ZN(new_n786));
  INV_X1    g361(.A(G1348), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n782), .A2(new_n783), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n784), .B(new_n790), .C1(new_n787), .C2(new_n786), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n682), .A2(G19), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n551), .B2(new_n682), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1341), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT94), .B(KEYINPUT23), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n682), .A2(G20), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G299), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n682), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1956), .ZN(new_n800));
  AOI211_X1 g375(.A(new_n794), .B(new_n800), .C1(new_n788), .C2(new_n789), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n791), .B(new_n801), .C1(new_n775), .C2(new_n774), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n777), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n709), .A2(new_n718), .A3(new_n720), .A4(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n745), .A2(G2072), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n623), .A2(new_n721), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(G311));
  AND3_X1   g383(.A1(new_n709), .A2(new_n720), .A3(new_n803), .ZN(new_n809));
  INV_X1    g384(.A(new_n807), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n809), .A2(new_n805), .A3(new_n810), .A4(new_n718), .ZN(G150));
  AOI22_X1  g386(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n538), .ZN(new_n813));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  INV_X1    g389(.A(G55), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n523), .A2(new_n814), .B1(new_n525), .B2(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NOR2_X1   g394(.A1(new_n600), .A2(new_n608), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n817), .A2(KEYINPUT95), .ZN(new_n823));
  OR3_X1    g398(.A1(new_n813), .A2(new_n816), .A3(KEYINPUT95), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n551), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n550), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n822), .B(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n819), .B1(new_n830), .B2(G860), .ZN(G145));
  NAND2_X1  g406(.A1(new_n486), .A2(G130), .ZN(new_n832));
  INV_X1    g407(.A(G142), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n463), .A2(G118), .ZN(new_n835));
  OAI221_X1 g410(.A(new_n832), .B1(new_n833), .B2(new_n483), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n616), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n699), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT96), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n744), .B(new_n715), .ZN(new_n841));
  AOI22_X1  g416(.A1(G126), .A2(new_n486), .B1(new_n491), .B2(new_n495), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n505), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n764), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n841), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n479), .B(new_n623), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(G162), .Z(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n845), .A2(KEYINPUT98), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n845), .A2(KEYINPUT98), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n853), .A3(new_n838), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n848), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT99), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n848), .A2(KEYINPUT99), .A3(new_n851), .A4(new_n854), .ZN(new_n858));
  AOI21_X1  g433(.A(G37), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n848), .B1(new_n845), .B2(new_n840), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n850), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g438(.A(G305), .B(G303), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT101), .ZN(new_n865));
  XNOR2_X1  g440(.A(G288), .B(new_n589), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n610), .B(KEYINPUT100), .Z(new_n868));
  AND2_X1   g443(.A1(new_n868), .A2(new_n829), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n829), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n601), .A2(G299), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n600), .A2(new_n798), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n874), .B1(new_n869), .B2(new_n870), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n867), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(new_n867), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n880), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n886), .A3(G868), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT102), .B1(new_n817), .B2(new_n604), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(new_n887), .ZN(G295));
  AOI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n887), .ZN(G331));
  NAND2_X1  g467(.A1(new_n826), .A2(new_n550), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n551), .A2(new_n823), .A3(new_n824), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n893), .A2(new_n894), .A3(G301), .ZN(new_n895));
  AOI21_X1  g470(.A(G301), .B1(new_n893), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(G286), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(G171), .B1(new_n825), .B2(new_n827), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n894), .A3(G301), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(G168), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n876), .A2(new_n901), .A3(KEYINPUT103), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT103), .B1(new_n876), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n897), .A2(new_n900), .A3(new_n874), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n867), .A4(new_n906), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n895), .A2(new_n896), .A3(G286), .ZN(new_n908));
  AOI21_X1  g483(.A(G168), .B1(new_n898), .B2(new_n899), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n874), .A2(new_n875), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT41), .B1(new_n872), .B2(new_n873), .ZN(new_n911));
  OAI22_X1  g486(.A1(new_n908), .A2(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n876), .A2(new_n901), .A3(KEYINPUT103), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n914), .A2(new_n867), .A3(new_n906), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT104), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n906), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n885), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n907), .A2(new_n917), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n912), .A2(new_n906), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n885), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n907), .A2(new_n917), .A3(new_n918), .A4(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(new_n922), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT105), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n921), .A2(new_n932), .A3(KEYINPUT43), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n928), .B1(new_n935), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g511(.A(G40), .ZN(new_n937));
  NOR4_X1   g512(.A1(new_n477), .A2(new_n464), .A3(new_n937), .A4(new_n470), .ZN(new_n938));
  AOI21_X1  g513(.A(G1384), .B1(new_n842), .B2(new_n505), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n507), .A2(new_n940), .A3(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n938), .B(KEYINPUT113), .C1(new_n939), .C2(new_n940), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(KEYINPUT116), .B(G1956), .Z(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT57), .ZN(new_n950));
  NAND2_X1  g525(.A1(G299), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n567), .A2(new_n562), .A3(new_n559), .A4(KEYINPUT57), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n471), .A2(G40), .A3(new_n478), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n507), .A2(new_n944), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n939), .A2(KEYINPUT45), .ZN(new_n958));
  XNOR2_X1  g533(.A(KEYINPUT56), .B(G2072), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n949), .A2(new_n953), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n949), .A2(new_n960), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n953), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n949), .A2(KEYINPUT119), .A3(new_n960), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT120), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n965), .A2(KEYINPUT120), .A3(new_n966), .A4(new_n967), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n955), .A2(new_n956), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n938), .A4(new_n958), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT121), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT58), .B(G1341), .Z(new_n977));
  INV_X1    g552(.A(new_n939), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(new_n954), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT118), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n978), .A2(KEYINPUT118), .A3(new_n954), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT121), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n957), .A2(new_n984), .A3(new_n974), .A4(new_n958), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n976), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n551), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT59), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT59), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n989), .A3(new_n551), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n961), .A2(KEYINPUT117), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n949), .A2(new_n993), .A3(new_n960), .A4(new_n953), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n963), .A2(new_n966), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n991), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT123), .B1(new_n972), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n962), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n949), .A2(KEYINPUT119), .A3(new_n960), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT119), .B1(new_n949), .B2(new_n960), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT120), .B1(new_n1004), .B2(new_n966), .ZN(new_n1005));
  INV_X1    g580(.A(new_n971), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1001), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT123), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n988), .A2(new_n990), .B1(new_n996), .B2(new_n997), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n981), .A2(G2067), .A3(new_n982), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n939), .A2(new_n940), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n938), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1011), .B1(new_n787), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1015), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n600), .B1(new_n1015), .B2(KEYINPUT60), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n1016), .A2(new_n1017), .B1(KEYINPUT60), .B2(new_n1015), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1000), .A2(new_n1010), .A3(new_n1018), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n1005), .A2(new_n1006), .B1(new_n600), .B2(new_n1015), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(new_n992), .A3(new_n994), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT124), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n678), .A2(G1976), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n979), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  OR3_X1    g603(.A1(new_n1024), .A2(KEYINPUT52), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G305), .A2(G1981), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n524), .A2(G86), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n673), .B1(new_n582), .B2(new_n1033), .ZN(new_n1034));
  OR3_X1    g609(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1032), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1026), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1029), .A2(new_n1030), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G303), .A2(G8), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT107), .B(G1971), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT106), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n957), .A2(new_n1045), .A3(new_n958), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n957), .B2(new_n958), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n947), .A2(G2090), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1049), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1048), .B1(G2090), .B2(new_n1014), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1042), .B(KEYINPUT109), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(G8), .A3(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1046), .A2(new_n1047), .A3(G2078), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1058), .A2(KEYINPUT53), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n954), .B1(new_n978), .B2(new_n956), .ZN(new_n1060));
  INV_X1    g635(.A(G2078), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n1061), .A4(new_n958), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1014), .A2(new_n775), .ZN(new_n1063));
  XOR2_X1   g638(.A(G171), .B(KEYINPUT54), .Z(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1059), .A2(new_n1062), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  AND4_X1   g641(.A1(new_n1039), .A2(new_n1054), .A3(new_n1057), .A4(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT115), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n507), .A2(new_n1070), .A3(KEYINPUT45), .A4(new_n944), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n1061), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1059), .B(new_n1063), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1064), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G168), .A2(new_n1025), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT126), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1069), .A2(new_n1060), .A3(new_n1071), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  INV_X1    g657(.A(G2084), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1012), .A2(new_n1083), .A3(new_n938), .A4(new_n1013), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1082), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1078), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT125), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1025), .B1(new_n1090), .B2(new_n1085), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT51), .B(new_n1088), .C1(new_n1091), .C2(new_n1078), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1025), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1078), .A2(KEYINPUT51), .A3(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1092), .A2(KEYINPUT127), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT127), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1067), .B(new_n1075), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1019), .A2(new_n1099), .A3(new_n1021), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1023), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1037), .A2(new_n1027), .A3(new_n678), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1031), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT111), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1026), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1038), .B(KEYINPUT110), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n1057), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT112), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1106), .B(KEYINPUT112), .C1(new_n1107), .C2(new_n1057), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1054), .A2(new_n1039), .A3(new_n1057), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1093), .A2(G168), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1107), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1055), .A2(G8), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1118), .B2(new_n1042), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1117), .A2(new_n1057), .A3(new_n1113), .A4(new_n1119), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1110), .A2(new_n1111), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  AOI21_X1  g698(.A(G301), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT62), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1112), .A3(new_n1074), .A4(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1101), .A2(new_n1121), .A3(new_n1126), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n939), .A2(new_n954), .A3(KEYINPUT45), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n764), .B(G2067), .Z(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n715), .B(G1996), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n699), .A2(new_n701), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n699), .A2(new_n701), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1986), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1137), .B1(new_n1138), .B2(new_n589), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G290), .A2(G1986), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1128), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1127), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1128), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n764), .A2(G2067), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1128), .B1(new_n1130), .B2(new_n715), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1128), .A2(KEYINPUT46), .A3(new_n974), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT46), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1143), .B2(G1996), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT47), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n1136), .A2(new_n1128), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1140), .A2(new_n1128), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT48), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1146), .B(new_n1152), .C1(new_n1153), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1142), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g732(.A(G229), .ZN(new_n1159));
  OAI21_X1  g733(.A(new_n654), .B1(new_n637), .B2(new_n638), .ZN(new_n1160));
  AOI21_X1  g734(.A(new_n1160), .B1(new_n859), .B2(new_n861), .ZN(new_n1161));
  NAND4_X1  g735(.A1(new_n934), .A2(G319), .A3(new_n1159), .A4(new_n1161), .ZN(G225));
  INV_X1    g736(.A(G225), .ZN(G308));
endmodule


