//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT93), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT92), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n191), .B2(new_n193), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n195), .A2(new_n196), .A3(G134), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n192), .A2(G143), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n190), .A2(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT92), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n198), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n189), .B1(new_n197), .B2(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT68), .A2(G116), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT68), .A2(G116), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(G122), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G122), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n207), .A2(G107), .A3(new_n209), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(KEYINPUT14), .A3(G107), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(G134), .B1(new_n195), .B2(new_n196), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n201), .A2(new_n198), .A3(new_n202), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT93), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n207), .A2(KEYINPUT14), .A3(G107), .A4(new_n209), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n204), .A2(new_n215), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  XOR2_X1   g034(.A(KEYINPUT91), .B(KEYINPUT13), .Z(new_n221));
  AOI21_X1  g035(.A(new_n198), .B1(new_n221), .B2(new_n199), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n191), .A2(new_n193), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(new_n221), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n224), .A2(new_n217), .A3(new_n212), .A4(new_n213), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT9), .B(G234), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n227), .A2(new_n228), .A3(G953), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n220), .A2(new_n225), .A3(new_n229), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(KEYINPUT94), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G902), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT94), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n226), .A2(new_n235), .A3(new_n230), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G478), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(G475), .A2(G902), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT16), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT76), .A2(G125), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT76), .A2(G125), .ZN(new_n248));
  OAI21_X1  g062(.A(G140), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OR2_X1    g063(.A1(G125), .A2(G140), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n247), .A2(new_n248), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n252), .A2(KEYINPUT16), .A3(G140), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n245), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G140), .ZN(new_n255));
  OR2_X1    g069(.A1(KEYINPUT76), .A2(G125), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT76), .A2(G125), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n250), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT16), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n257), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(new_n246), .A3(new_n255), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(G146), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(G237), .A2(G953), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n264), .A2(G143), .A3(G214), .ZN(new_n265));
  AOI21_X1  g079(.A(G143), .B1(new_n264), .B2(G214), .ZN(new_n266));
  OAI21_X1  g080(.A(G131), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT17), .ZN(new_n268));
  INV_X1    g082(.A(G237), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G214), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n190), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n264), .A2(G143), .A3(G214), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n267), .A2(new_n268), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n274), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT17), .A3(G131), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n254), .A2(new_n263), .A3(new_n276), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT18), .A2(G131), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n272), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT90), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT90), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n272), .A2(new_n283), .A3(new_n274), .A4(new_n280), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT77), .ZN(new_n286));
  NAND2_X1  g100(.A1(G125), .A2(G140), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n250), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n250), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n245), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n249), .A2(G146), .A3(new_n250), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n277), .A2(KEYINPUT18), .A3(G131), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n285), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(G113), .B(G122), .ZN(new_n295));
  INV_X1    g109(.A(G104), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n295), .B(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n279), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT19), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n288), .B2(new_n289), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n249), .A2(KEYINPUT19), .A3(new_n250), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n245), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n267), .A2(new_n275), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n263), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n297), .B1(new_n304), .B2(new_n294), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n244), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT20), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT20), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n308), .B(new_n244), .C1(new_n298), .C2(new_n305), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n297), .B1(new_n279), .B2(new_n294), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n234), .B1(new_n298), .B2(new_n310), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n307), .A2(new_n309), .B1(G475), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n242), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n233), .A2(new_n234), .A3(new_n236), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n270), .A2(G952), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G234), .B2(G237), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT21), .B(G898), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(G234), .A2(G237), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(G902), .A3(G953), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n317), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT96), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n243), .A2(new_n312), .A3(new_n314), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n245), .A2(G143), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n190), .A2(G146), .ZN(new_n326));
  AND4_X1   g140(.A1(KEYINPUT0), .A2(new_n325), .A3(new_n326), .A4(G128), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n245), .B2(G143), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n190), .A2(KEYINPUT65), .A3(G146), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT64), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(G143), .B2(new_n245), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n329), .B(new_n330), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  XOR2_X1   g148(.A(KEYINPUT0), .B(G128), .Z(new_n335));
  AOI211_X1 g149(.A(new_n252), .B(new_n327), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n192), .B1(new_n325), .B2(KEYINPUT1), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n325), .A2(new_n326), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n340), .A2(KEYINPUT1), .A3(new_n192), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n261), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT7), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n270), .A2(G224), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI22_X1  g160(.A1(new_n336), .A2(new_n343), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n327), .B1(new_n334), .B2(new_n335), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n261), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n346), .A2(new_n344), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n329), .A2(new_n330), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT64), .B1(new_n190), .B2(G146), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n331), .A2(new_n245), .A3(G143), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n337), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(new_n341), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n349), .B(new_n350), .C1(new_n356), .C2(new_n261), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(new_n296), .B2(G107), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n211), .A3(G104), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n296), .A2(G107), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G101), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n365), .A2(KEYINPUT4), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(KEYINPUT4), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(KEYINPUT79), .ZN(new_n370));
  INV_X1    g184(.A(G101), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n359), .A2(new_n361), .A3(new_n371), .A4(new_n362), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n363), .A2(new_n373), .A3(G101), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(KEYINPUT4), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  OR2_X1    g189(.A1(KEYINPUT67), .A2(G119), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT67), .A2(G119), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(G116), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n205), .A2(G119), .A3(new_n206), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT2), .B(G113), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n381), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n378), .A3(new_n379), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n369), .A2(new_n375), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n211), .A2(G104), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n296), .A2(G107), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n372), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n390), .A2(new_n384), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n376), .A2(new_n392), .A3(G116), .A4(new_n377), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n393), .A2(G113), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT5), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n394), .A2(KEYINPUT87), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT87), .B1(new_n394), .B2(new_n395), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n391), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G122), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n386), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n358), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n399), .B(KEYINPUT8), .Z(new_n402));
  OAI21_X1  g216(.A(new_n384), .B1(new_n396), .B2(new_n397), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n372), .A2(new_n389), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n395), .B1(new_n394), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n394), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT88), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n391), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n402), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n234), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT89), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n386), .A2(new_n398), .ZN(new_n414));
  INV_X1    g228(.A(new_n399), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n400), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n418), .A3(new_n415), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n336), .A2(new_n343), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(new_n346), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT89), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(new_n234), .C1(new_n401), .C2(new_n411), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n413), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G210), .B1(G237), .B2(G902), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n413), .A2(new_n422), .A3(new_n426), .A4(new_n424), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n188), .B(new_n324), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G221), .B1(new_n227), .B2(G902), .ZN(new_n431));
  XNOR2_X1  g245(.A(G110), .B(G140), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n270), .A2(G227), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT12), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n339), .A2(new_n342), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(new_n390), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(KEYINPUT1), .C1(new_n190), .C2(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G128), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n438), .B1(new_n325), .B2(KEYINPUT1), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n340), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(KEYINPUT82), .B(new_n340), .C1(new_n440), .C2(new_n441), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n342), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n437), .B1(new_n390), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT11), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n198), .B2(G137), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n198), .A2(G137), .ZN(new_n450));
  INV_X1    g264(.A(G137), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT11), .A3(G134), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(KEYINPUT66), .A3(G131), .ZN(new_n454));
  NAND2_X1  g268(.A1(KEYINPUT66), .A2(G131), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n449), .A2(new_n452), .A3(new_n455), .A4(new_n450), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n435), .B1(new_n447), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n446), .A2(new_n390), .ZN(new_n460));
  OAI211_X1 g274(.A(KEYINPUT12), .B(new_n457), .C1(new_n460), .C2(new_n437), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n446), .A2(new_n390), .ZN(new_n462));
  XOR2_X1   g276(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n390), .B(KEYINPUT10), .C1(new_n355), .C2(new_n341), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n436), .A2(KEYINPUT84), .A3(KEYINPUT10), .A4(new_n390), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n369), .A2(new_n375), .A3(new_n348), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n464), .A2(new_n469), .A3(new_n458), .A4(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n372), .A2(KEYINPUT4), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(KEYINPUT79), .B2(new_n364), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n368), .B1(new_n475), .B2(new_n374), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n348), .A2(new_n476), .B1(new_n467), .B2(new_n468), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n477), .A2(KEYINPUT85), .A3(new_n458), .A4(new_n464), .ZN(new_n478));
  AOI221_X4 g292(.A(new_n434), .B1(new_n459), .B2(new_n461), .C1(new_n473), .C2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n434), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n473), .A2(new_n478), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(new_n464), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n457), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT86), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n473), .A2(new_n478), .B1(new_n459), .B2(new_n461), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT86), .B1(new_n486), .B2(new_n480), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI211_X1 g302(.A(G469), .B(G902), .C1(new_n485), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G469), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n480), .A3(new_n483), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n480), .B2(new_n486), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n490), .B1(new_n492), .B2(new_n234), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n430), .B(new_n431), .C1(new_n489), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT97), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT72), .ZN(new_n496));
  INV_X1    g310(.A(new_n385), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n348), .A2(new_n457), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n451), .A2(G134), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n273), .B1(new_n198), .B2(G137), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n453), .A2(new_n273), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT69), .ZN(new_n502));
  OAI22_X1  g316(.A1(new_n355), .A2(new_n341), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n453), .A2(new_n273), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n499), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(KEYINPUT69), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n497), .B(new_n498), .C1(new_n503), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT28), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n498), .B1(new_n356), .B2(new_n501), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n385), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(KEYINPUT69), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n501), .A2(new_n502), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n436), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n497), .A4(new_n498), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n510), .B1(new_n519), .B2(KEYINPUT28), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n264), .A2(G210), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT27), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(G101), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(KEYINPUT30), .B(new_n498), .C1(new_n503), .C2(new_n507), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT70), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT70), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n516), .A2(new_n529), .A3(KEYINPUT30), .A4(new_n498), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n436), .A2(new_n506), .B1(new_n348), .B2(new_n457), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n385), .B1(new_n532), .B2(KEYINPUT30), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n511), .A2(new_n518), .A3(new_n525), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT31), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT31), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n533), .B1(new_n528), .B2(new_n530), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n511), .A2(new_n518), .A3(new_n525), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n521), .A2(new_n526), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G472), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n234), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n496), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT31), .B1(new_n535), .B2(new_n536), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n539), .A2(new_n540), .A3(new_n538), .ZN(new_n547));
  OAI22_X1  g361(.A1(new_n546), .A2(new_n547), .B1(new_n520), .B2(new_n525), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n548), .A2(KEYINPUT72), .A3(new_n543), .A4(new_n234), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT32), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n548), .A2(KEYINPUT32), .A3(new_n543), .A4(new_n234), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT29), .B1(new_n520), .B2(new_n525), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n511), .A2(new_n518), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n554), .B(new_n526), .C1(new_n539), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n526), .B1(new_n539), .B2(new_n555), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT73), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n516), .A2(new_n498), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n511), .B(new_n518), .C1(new_n497), .C2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n510), .B1(new_n561), .B2(KEYINPUT28), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n525), .A2(KEYINPUT29), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G472), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n551), .A2(new_n552), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n228), .B1(G234), .B2(new_n234), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT78), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT22), .B(G137), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n254), .A2(new_n263), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n376), .A2(G128), .A3(new_n377), .ZN(new_n575));
  INV_X1    g389(.A(G119), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n575), .B1(new_n576), .B2(G128), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT24), .B(G110), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(G128), .B1(new_n376), .B2(new_n377), .ZN(new_n584));
  AOI22_X1  g398(.A1(KEYINPUT74), .A2(new_n584), .B1(new_n575), .B2(KEYINPUT23), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n376), .A2(new_n377), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n192), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n576), .A2(G128), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT23), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT75), .B1(new_n593), .B2(G110), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n585), .A2(new_n589), .B1(KEYINPUT23), .B2(new_n591), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n596));
  INV_X1    g410(.A(G110), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n583), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n263), .A2(new_n290), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n595), .A2(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n577), .A2(new_n579), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n573), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n593), .A2(KEYINPUT75), .A3(G110), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n582), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n573), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n608), .A2(new_n603), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n234), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT25), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n599), .A2(new_n604), .A3(new_n573), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n609), .B1(new_n608), .B2(new_n603), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(KEYINPUT25), .A3(new_n234), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n569), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n616), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n568), .A2(G902), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n567), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n431), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT86), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n481), .A2(new_n483), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n434), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n459), .A2(new_n461), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n481), .A2(new_n480), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n627), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n490), .B(new_n234), .C1(new_n632), .C2(new_n487), .ZN(new_n633));
  INV_X1    g447(.A(new_n493), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n626), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n636), .A3(new_n430), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n495), .A2(new_n625), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G101), .ZN(G3));
  OAI21_X1  g453(.A(G472), .B1(new_n542), .B2(G902), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(KEYINPUT98), .B(G472), .C1(new_n542), .C2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n545), .A2(new_n549), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n623), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n648), .A2(new_n635), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n429), .A2(KEYINPUT99), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n188), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n428), .A2(KEYINPUT99), .A3(new_n429), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT33), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n233), .A2(new_n654), .A3(new_n236), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n231), .A2(KEYINPUT33), .A3(new_n232), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(G478), .A3(new_n234), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n237), .A2(new_n238), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n312), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n653), .A2(new_n323), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n649), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  NAND2_X1  g477(.A1(new_n307), .A2(new_n309), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT100), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n243), .A2(new_n314), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n311), .A2(G475), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(new_n651), .A3(new_n323), .A4(new_n652), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n649), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G107), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  AOI21_X1  g490(.A(KEYINPUT25), .B1(new_n616), .B2(new_n234), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n612), .B(G902), .C1(new_n614), .C2(new_n615), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n568), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n599), .A2(new_n604), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n620), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n679), .A2(KEYINPUT102), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT102), .B1(new_n679), .B2(new_n683), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n686), .A2(new_n645), .A3(new_n644), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n495), .A2(new_n637), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT37), .B(G110), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G12));
  OAI21_X1  g504(.A(new_n317), .B1(G900), .B2(new_n321), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n668), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n665), .A2(new_n667), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n635), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n567), .A2(new_n653), .A3(new_n686), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n192), .ZN(G30));
  XNOR2_X1  g511(.A(new_n691), .B(KEYINPUT39), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n635), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n539), .A2(new_n555), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n526), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n234), .B1(new_n561), .B2(new_n525), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n551), .A2(new_n552), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n679), .A3(new_n683), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n428), .A2(new_n429), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT38), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n667), .A2(new_n312), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n710), .A2(new_n187), .A3(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n700), .A2(new_n701), .A3(new_n708), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT103), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n190), .ZN(G45));
  NAND2_X1  g529(.A1(new_n659), .A2(new_n691), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n635), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(new_n695), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  AOI22_X1  g534(.A1(new_n473), .A2(new_n478), .B1(new_n457), .B2(new_n482), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n631), .B1(new_n480), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n487), .B1(new_n722), .B2(KEYINPUT86), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n723), .B2(G902), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n431), .A3(new_n633), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n624), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n660), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  AOI21_X1  g543(.A(KEYINPUT104), .B1(new_n726), .B2(new_n672), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n624), .A2(new_n725), .A3(new_n671), .A4(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n733), .B(G116), .Z(G18));
  INV_X1    g548(.A(new_n324), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n567), .A2(new_n735), .A3(new_n686), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n651), .A2(new_n652), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n725), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT105), .B(G119), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G21));
  NAND3_X1  g555(.A1(new_n651), .A2(new_n652), .A3(new_n711), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  OAI22_X1  g557(.A1(new_n546), .A2(new_n547), .B1(new_n562), .B2(new_n525), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n543), .A3(new_n234), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n623), .A2(new_n323), .A3(new_n640), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT106), .B1(new_n747), .B2(new_n725), .ZN(new_n748));
  INV_X1    g562(.A(new_n725), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n743), .A4(new_n746), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NAND2_X1  g567(.A1(new_n724), .A2(new_n633), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n679), .A2(new_n683), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n640), .A2(new_n717), .A3(new_n756), .A4(new_n745), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n755), .A2(new_n757), .A3(new_n431), .A4(new_n653), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G125), .ZN(G27));
  OAI21_X1  g573(.A(new_n550), .B1(new_n542), .B2(new_n544), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n552), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n543), .B1(new_n559), .B2(new_n564), .ZN(new_n762));
  OAI211_X1 g576(.A(KEYINPUT107), .B(new_n623), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n566), .A2(new_n552), .A3(new_n760), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT107), .B1(new_n765), .B2(new_n623), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n709), .A2(new_n188), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n635), .A2(new_n717), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT42), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n625), .A2(new_n635), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  NAND4_X1  g588(.A1(new_n625), .A2(new_n635), .A3(new_n693), .A4(new_n768), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  INV_X1    g590(.A(KEYINPUT46), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n490), .B1(new_n492), .B2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n491), .B(KEYINPUT45), .C1(new_n480), .C2(new_n486), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(KEYINPUT108), .A3(new_n780), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n490), .A2(new_n234), .ZN(new_n786));
  OAI211_X1 g600(.A(KEYINPUT109), .B(new_n777), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n783), .B2(new_n784), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n788), .B1(new_n789), .B2(KEYINPUT46), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n489), .B1(new_n789), .B2(KEYINPUT46), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n787), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n792), .A2(new_n431), .A3(new_n698), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n657), .A2(new_n658), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n312), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT43), .Z(new_n796));
  AND3_X1   g610(.A1(new_n796), .A2(new_n646), .A3(new_n756), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n797), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT110), .B1(new_n797), .B2(KEYINPUT44), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(KEYINPUT44), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n799), .A2(new_n768), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n793), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  NAND3_X1  g617(.A1(new_n768), .A2(new_n647), .A3(new_n717), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n567), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n431), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT47), .B1(new_n792), .B2(new_n431), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  XOR2_X1   g623(.A(new_n754), .B(KEYINPUT49), .Z(new_n810));
  NAND3_X1  g624(.A1(new_n623), .A2(new_n431), .A3(new_n187), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n710), .A2(new_n706), .A3(new_n795), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n726), .A2(new_n660), .B1(new_n736), .B2(new_n738), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n814), .B(new_n752), .C1(new_n730), .C2(new_n732), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n665), .A2(new_n666), .A3(new_n692), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n567), .A2(new_n686), .A3(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n635), .B(new_n768), .C1(new_n817), .C2(new_n757), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n770), .A2(new_n772), .A3(new_n818), .A4(new_n775), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n653), .A2(new_n431), .A3(new_n633), .A4(new_n724), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n756), .A2(new_n640), .A3(new_n745), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n717), .ZN(new_n823));
  OAI22_X1  g637(.A1(new_n695), .A2(new_n694), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n758), .B(KEYINPUT113), .C1(new_n695), .C2(new_n694), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n691), .B(KEYINPUT114), .Z(new_n829));
  NAND3_X1  g643(.A1(new_n743), .A2(new_n635), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n828), .B1(new_n831), .B2(new_n708), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n826), .A2(new_n827), .A3(new_n832), .A4(new_n719), .ZN(new_n833));
  OAI22_X1  g647(.A1(new_n830), .A2(new_n707), .B1(new_n718), .B2(new_n695), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n828), .B1(new_n834), .B2(new_n824), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n188), .B1(new_n428), .B2(new_n429), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n323), .A3(new_n659), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT111), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n837), .A2(new_n840), .A3(new_n323), .A4(new_n659), .ZN(new_n841));
  INV_X1    g655(.A(new_n312), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n667), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n837), .A2(new_n323), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n839), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n648), .A2(new_n845), .A3(new_n635), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n638), .A2(new_n688), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n638), .A2(new_n688), .A3(new_n846), .A4(KEYINPUT112), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n820), .A2(new_n836), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(KEYINPUT115), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n824), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n831), .A2(new_n708), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n719), .A3(KEYINPUT52), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n835), .ZN(new_n858));
  XOR2_X1   g672(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n820), .A2(new_n851), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT115), .B1(new_n852), .B2(new_n853), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT54), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n749), .A2(new_n768), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n706), .A2(new_n647), .A3(new_n317), .ZN(new_n866));
  INV_X1    g680(.A(new_n659), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n796), .A2(new_n316), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n640), .A2(new_n745), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n869), .A2(new_n647), .A3(new_n870), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n315), .B(new_n868), .C1(new_n738), .C2(new_n871), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n767), .A2(new_n865), .A3(KEYINPUT48), .A4(new_n869), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT48), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n865), .A2(new_n869), .ZN(new_n875));
  INV_X1    g689(.A(new_n767), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n872), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n865), .A2(new_n866), .A3(new_n842), .A4(new_n794), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n875), .A2(new_n822), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n710), .A2(new_n187), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n749), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT50), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n871), .A2(KEYINPUT50), .A3(new_n749), .A4(new_n881), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n879), .B(new_n880), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n754), .A2(new_n431), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n806), .A2(new_n807), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n871), .A2(new_n768), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT51), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n886), .B(new_n892), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n878), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n820), .A2(new_n851), .A3(new_n858), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n859), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n820), .A2(new_n836), .A3(new_n851), .A4(KEYINPUT53), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n864), .A2(new_n894), .A3(KEYINPUT117), .A4(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(G952), .A2(G953), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n899), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n852), .A2(new_n853), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n861), .A3(new_n854), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n907), .B2(KEYINPUT54), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT117), .B1(new_n908), .B2(new_n894), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n813), .B1(new_n902), .B2(new_n909), .ZN(G75));
  NAND2_X1  g724(.A1(new_n417), .A2(new_n419), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n421), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT55), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n234), .B1(new_n896), .B2(new_n898), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(G210), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n270), .A2(G952), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n916), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n916), .A2(new_n923), .ZN(new_n926));
  INV_X1    g740(.A(new_n921), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT119), .B1(new_n928), .B2(new_n918), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n925), .A2(new_n929), .ZN(G51));
  NAND2_X1  g744(.A1(new_n896), .A2(new_n898), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n897), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n786), .B(KEYINPUT120), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT57), .ZN(new_n934));
  OAI22_X1  g748(.A1(new_n932), .A2(new_n934), .B1(new_n632), .B2(new_n487), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n915), .A2(new_n785), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n921), .B1(new_n935), .B2(new_n938), .ZN(G54));
  NAND3_X1  g753(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n298), .A2(new_n305), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n927), .B1(new_n940), .B2(new_n943), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n940), .B2(new_n943), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G60));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT59), .Z(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n655), .A2(new_n656), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n927), .B1(new_n932), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n655), .A2(new_n656), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n864), .A2(new_n899), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n950), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n953), .B2(new_n955), .ZN(G63));
  XNOR2_X1  g770(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n228), .A2(new_n234), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n931), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n921), .B1(new_n960), .B2(new_n619), .ZN(new_n961));
  AND4_X1   g775(.A1(KEYINPUT124), .A2(new_n931), .A3(new_n682), .A4(new_n959), .ZN(new_n962));
  INV_X1    g776(.A(new_n959), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n896), .B2(new_n898), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT124), .B1(new_n964), .B2(new_n682), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n961), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n962), .B2(new_n965), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI221_X1 g784(.A(new_n961), .B1(new_n967), .B2(KEYINPUT61), .C1(new_n962), .C2(new_n965), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(G66));
  NAND3_X1  g786(.A1(new_n319), .A2(G224), .A3(G953), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n815), .B1(new_n849), .B2(new_n850), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n975), .B2(G953), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n911), .B1(G898), .B2(new_n270), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT126), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n976), .B(new_n978), .ZN(G69));
  AND2_X1   g793(.A1(new_n826), .A2(new_n719), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n773), .A2(new_n980), .A3(new_n775), .A4(new_n827), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n793), .A2(new_n743), .A3(new_n876), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n981), .A2(new_n802), .A3(new_n982), .A4(new_n808), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(G953), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n531), .B1(KEYINPUT30), .B2(new_n532), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n300), .A2(new_n301), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(G900), .A2(G953), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n980), .A2(new_n827), .ZN(new_n992));
  OR3_X1    g806(.A1(new_n714), .A2(new_n992), .A3(KEYINPUT62), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT62), .B1(new_n714), .B2(new_n992), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n843), .A2(new_n659), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n997), .A2(KEYINPUT127), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n768), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  OR4_X1    g814(.A1(new_n624), .A2(new_n699), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n808), .A2(new_n802), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(G953), .B1(new_n995), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n991), .B1(new_n1003), .B2(new_n987), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n270), .B1(G227), .B2(G900), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1005), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n991), .B(new_n1007), .C1(new_n1003), .C2(new_n987), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(G72));
  AND3_X1   g823(.A1(new_n995), .A2(new_n974), .A3(new_n1002), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n703), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n539), .A2(new_n540), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n558), .A2(new_n556), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n907), .B(new_n1012), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1012), .B1(new_n983), .B2(new_n975), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n539), .A2(new_n555), .A3(new_n525), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n921), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1014), .A2(new_n1017), .A3(new_n1020), .ZN(G57));
endmodule


