//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  XOR2_X1   g008(.A(new_n208), .B(new_n209), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT69), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(KEYINPUT69), .A3(new_n209), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT78), .B(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT2), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  INV_X1    g018(.A(G155gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(new_n217), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n223), .B(KEYINPUT77), .Z(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT76), .B(G141gat), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  OAI221_X1 g025(.A(new_n218), .B1(new_n219), .B2(new_n221), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n229));
  INV_X1    g028(.A(new_n219), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n221), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G141gat), .B(G148gat), .ZN(new_n232));
  OAI221_X1 g031(.A(new_n231), .B1(new_n229), .B2(new_n230), .C1(KEYINPUT2), .C2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n227), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT71), .B(KEYINPUT29), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n214), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT84), .ZN(new_n238));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n212), .A2(new_n213), .ZN(new_n240));
  INV_X1    g039(.A(new_n234), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n235), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT84), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n233), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n240), .B2(KEYINPUT29), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n228), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n240), .A2(new_n247), .A3(KEYINPUT29), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n210), .A2(new_n235), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n246), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n242), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n239), .B(KEYINPUT82), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G78gat), .B(G106gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT31), .B(G50gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT85), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n202), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n261), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n265), .B1(new_n252), .B2(new_n257), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n266), .A2(KEYINPUT85), .A3(G22gat), .ZN(new_n267));
  OAI22_X1  g066(.A1(new_n264), .A2(new_n267), .B1(new_n258), .B2(new_n261), .ZN(new_n268));
  XNOR2_X1  g067(.A(G15gat), .B(G43gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(G71gat), .B(G99gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n273));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(KEYINPUT23), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(KEYINPUT23), .B2(new_n276), .ZN(new_n278));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n273), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n284), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n274), .A2(KEYINPUT25), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288));
  INV_X1    g087(.A(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n287), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(KEYINPUT65), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n286), .B(new_n292), .C1(new_n293), .C2(new_n288), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n275), .B1(KEYINPUT26), .B2(new_n291), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n293), .B2(KEYINPUT26), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT27), .B(G183gat), .Z(new_n298));
  OR3_X1    g097(.A1(new_n298), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT28), .B1(new_n298), .B2(G190gat), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n279), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(G113gat), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(G120gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n304), .B1(new_n307), .B2(KEYINPUT66), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(KEYINPUT66), .B2(new_n307), .ZN(new_n309));
  XOR2_X1   g108(.A(G127gat), .B(G134gat), .Z(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(KEYINPUT1), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n306), .A2(new_n304), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n310), .B1(new_n313), .B2(KEYINPUT1), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n302), .B(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(G227gat), .A2(G233gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n272), .B1(new_n318), .B2(KEYINPUT32), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT67), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT33), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  AOI211_X1 g121(.A(KEYINPUT67), .B(KEYINPUT33), .C1(new_n316), .C2(new_n317), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n319), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n318), .B(KEYINPUT32), .C1(new_n321), .C2(new_n272), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT34), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n316), .A2(new_n317), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT34), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n329), .A3(new_n325), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n262), .A2(new_n263), .A3(new_n202), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n258), .A2(new_n261), .ZN(new_n333));
  OAI21_X1  g132(.A(G22gat), .B1(new_n266), .B2(KEYINPUT85), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n330), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n317), .B2(new_n316), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n268), .A2(new_n331), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n302), .B(KEYINPUT70), .Z(new_n339));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n302), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n340), .B1(new_n343), .B2(KEYINPUT29), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n345), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n214), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n339), .A2(new_n340), .A3(new_n236), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n341), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n240), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G92gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT73), .B(G64gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(KEYINPUT30), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n214), .B1(new_n350), .B2(new_n351), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n214), .B2(new_n348), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n358), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n362), .B2(new_n358), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n354), .A2(KEYINPUT74), .A3(new_n359), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT35), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373));
  INV_X1    g172(.A(G85gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n227), .A2(new_n233), .A3(new_n314), .A4(new_n312), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT4), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n315), .A3(new_n234), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n385));
  NAND2_X1  g184(.A1(new_n246), .A2(new_n315), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n379), .ZN(new_n387));
  INV_X1    g186(.A(new_n381), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n380), .A2(new_n381), .A3(new_n383), .A4(new_n385), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n378), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT80), .B1(new_n384), .B2(new_n389), .ZN(new_n393));
  OAI211_X1 g192(.A(KEYINPUT6), .B(new_n377), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n377), .B1(new_n392), .B2(new_n393), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT87), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n392), .A2(new_n393), .ZN(new_n398));
  INV_X1    g197(.A(new_n377), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT6), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n395), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  OR3_X1    g200(.A1(new_n338), .A2(new_n372), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n396), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n394), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n370), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n403), .B1(new_n370), .B2(new_n405), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n406), .A2(new_n407), .A3(new_n338), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n408), .B2(new_n371), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n268), .A2(new_n335), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n406), .B2(new_n407), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT37), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n359), .B1(new_n354), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n350), .A2(new_n214), .A3(new_n351), .ZN(new_n414));
  OAI211_X1 g213(.A(KEYINPUT37), .B(new_n414), .C1(new_n348), .C2(new_n214), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(KEYINPUT38), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n413), .B(new_n418), .C1(new_n416), .C2(new_n415), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n413), .B1(new_n412), .B2(new_n354), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT38), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n401), .A2(new_n419), .A3(new_n368), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n368), .A2(new_n369), .ZN(new_n423));
  INV_X1    g222(.A(new_n364), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT86), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n380), .A2(new_n383), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(new_n388), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n426), .A3(new_n388), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n386), .A2(new_n381), .A3(new_n379), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n429), .A2(KEYINPUT39), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n430), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(new_n428), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n432), .B(new_n399), .C1(KEYINPUT39), .C2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT40), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n425), .A2(new_n397), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n410), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n337), .A2(new_n331), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT36), .B1(new_n440), .B2(KEYINPUT68), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT68), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n442), .B(new_n443), .C1(new_n337), .C2(new_n331), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n411), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n409), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G113gat), .B(G141gat), .ZN(new_n448));
  INV_X1    g247(.A(G197gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT11), .B(G169gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  XOR2_X1   g251(.A(new_n452), .B(KEYINPUT12), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT93), .ZN(new_n455));
  XOR2_X1   g254(.A(G15gat), .B(G22gat), .Z(new_n456));
  INV_X1    g255(.A(G1gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G15gat), .B(G22gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT16), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(G1gat), .ZN(new_n461));
  INV_X1    g260(.A(G8gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n458), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n466), .B(G8gat), .C1(new_n465), .C2(new_n461), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT92), .ZN(new_n468));
  INV_X1    g267(.A(new_n461), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n462), .B1(new_n469), .B2(KEYINPUT91), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n466), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n464), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G43gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G50gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT15), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G43gat), .B(G50gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g280(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT90), .ZN(new_n484));
  AND2_X1   g283(.A1(G29gat), .A2(G36gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n479), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(KEYINPUT15), .B(new_n478), .C1(new_n483), .C2(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n455), .B1(new_n473), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n472), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n471), .B1(new_n470), .B2(new_n466), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n463), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT93), .A3(new_n490), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n490), .B(KEYINPUT17), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n492), .A2(new_n496), .B1(new_n473), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT18), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n454), .B1(new_n500), .B2(KEYINPUT95), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n492), .A2(new_n496), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n473), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n496), .A3(KEYINPUT94), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n473), .A2(new_n491), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n499), .B(KEYINPUT13), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n498), .A2(KEYINPUT18), .A3(new_n499), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n501), .A2(new_n506), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT95), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n453), .B1(new_n506), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n502), .A2(new_n507), .B1(new_n473), .B2(new_n491), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n512), .B1(new_n519), .B2(new_n509), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n506), .A2(new_n515), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G176gat), .B(G204gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT105), .ZN(new_n526));
  XNOR2_X1  g325(.A(G120gat), .B(G148gat), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  INV_X1    g327(.A(KEYINPUT96), .ZN(new_n529));
  XOR2_X1   g328(.A(G57gat), .B(G64gat), .Z(new_n530));
  XNOR2_X1  g329(.A(G71gat), .B(G78gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT9), .ZN(new_n532));
  INV_X1    g331(.A(G71gat), .ZN(new_n533));
  INV_X1    g332(.A(G78gat), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n531), .B1(new_n530), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n529), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n530), .A2(new_n535), .ZN(new_n539));
  INV_X1    g338(.A(new_n531), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT96), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G99gat), .B(G106gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT100), .ZN(new_n547));
  OR3_X1    g346(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT99), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n547), .B1(new_n546), .B2(KEYINPUT7), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n546), .A2(new_n552), .A3(KEYINPUT7), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n548), .A2(new_n550), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT101), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(KEYINPUT101), .A2(G99gat), .A3(G106gat), .ZN(new_n560));
  AOI211_X1 g359(.A(KEYINPUT102), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT102), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(new_n558), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(KEYINPUT8), .A3(new_n560), .ZN(new_n564));
  INV_X1    g363(.A(new_n555), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n545), .B(new_n554), .C1(new_n561), .C2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n554), .B1(new_n561), .B2(new_n566), .ZN(new_n568));
  INV_X1    g367(.A(new_n545), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n544), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n536), .A2(new_n537), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n567), .ZN(new_n574));
  OAI22_X1  g373(.A1(new_n571), .A2(KEYINPUT103), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT103), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n570), .A2(new_n576), .A3(new_n572), .A4(new_n567), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n538), .A2(new_n543), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n574), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT103), .B1(new_n574), .B2(new_n582), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n574), .A2(new_n573), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n583), .B(new_n577), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT104), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT104), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n575), .A2(new_n589), .A3(new_n583), .A4(new_n577), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n584), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n581), .B1(new_n591), .B2(new_n580), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT106), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n528), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n593), .A3(new_n528), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n524), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G127gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n220), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  INV_X1    g403(.A(G183gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n205), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n602), .B(G155gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n607), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n473), .B1(new_n613), .B2(new_n582), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n612), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n497), .A2(new_n574), .ZN(new_n618));
  NAND3_X1  g417(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n618), .B(new_n619), .C1(new_n491), .C2(new_n574), .ZN(new_n620));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621));
  AND2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT98), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(new_n622), .B2(new_n623), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n447), .A2(new_n598), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n405), .B(KEYINPUT107), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g437(.A1(new_n634), .A2(new_n425), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT42), .B1(new_n639), .B2(new_n462), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT16), .B(G8gat), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  MUX2_X1   g441(.A(KEYINPUT42), .B(new_n640), .S(new_n642), .Z(G1325gat));
  INV_X1    g442(.A(new_n440), .ZN(new_n644));
  AOI21_X1  g443(.A(G15gat), .B1(new_n634), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n445), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n646), .A2(G15gat), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n634), .B2(new_n647), .ZN(G1326gat));
  NAND2_X1  g447(.A1(new_n634), .A2(new_n410), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT108), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT43), .B(G22gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  INV_X1    g451(.A(new_n632), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n409), .B2(new_n446), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n598), .A2(new_n617), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n657), .A2(G29gat), .A3(new_n635), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT45), .Z(new_n659));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n447), .B2(new_n632), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n632), .B(KEYINPUT109), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI211_X1 g462(.A(KEYINPUT44), .B(new_n663), .C1(new_n409), .C2(new_n446), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n656), .ZN(new_n666));
  OAI21_X1  g465(.A(G29gat), .B1(new_n666), .B2(new_n635), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n659), .A2(new_n667), .ZN(G1328gat));
  OAI21_X1  g467(.A(G36gat), .B1(new_n666), .B2(new_n370), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n657), .A2(G36gat), .A3(new_n370), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT46), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(G1329gat));
  NOR3_X1   g471(.A1(new_n657), .A2(G43gat), .A3(new_n440), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n646), .B(new_n656), .C1(new_n661), .C2(new_n664), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(G43gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g475(.A1(new_n665), .A2(G50gat), .A3(new_n410), .A4(new_n656), .ZN(new_n677));
  INV_X1    g476(.A(G50gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n657), .B2(new_n438), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n677), .A2(KEYINPUT48), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT48), .B1(new_n677), .B2(new_n679), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(G1331gat));
  INV_X1    g481(.A(new_n597), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n617), .A2(new_n523), .A3(new_n632), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n683), .B(new_n685), .C1(new_n409), .C2(new_n446), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n636), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT110), .B(G57gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1332gat));
  AOI21_X1  g488(.A(new_n370), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT111), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(KEYINPUT111), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n694), .B(new_n696), .ZN(G1333gat));
  AOI21_X1  g496(.A(new_n533), .B1(new_n686), .B2(new_n646), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n440), .A2(G71gat), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n686), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n410), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G78gat), .ZN(G1335gat));
  INV_X1    g502(.A(new_n617), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n523), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n654), .B2(KEYINPUT112), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n707), .B(new_n653), .C1(new_n409), .C2(new_n446), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT51), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n411), .A2(new_n439), .A3(new_n445), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n338), .A2(new_n372), .A3(new_n401), .ZN(new_n711));
  INV_X1    g510(.A(new_n405), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT81), .B1(new_n425), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n338), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n370), .A2(new_n405), .A3(new_n403), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n711), .B1(new_n716), .B2(KEYINPUT35), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n632), .B1(new_n710), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n707), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n654), .A2(KEYINPUT112), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n705), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n709), .A2(new_n597), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n374), .A3(new_n636), .ZN(new_n724));
  INV_X1    g523(.A(new_n665), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n705), .A2(new_n597), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n725), .A2(new_n635), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n374), .B2(new_n727), .ZN(G1336gat));
  NOR2_X1   g527(.A1(new_n370), .A2(G92gat), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n709), .A2(new_n722), .A3(new_n597), .A4(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n726), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n425), .B(new_n731), .C1(new_n661), .C2(new_n664), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G92gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n730), .B(new_n733), .C1(new_n736), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1337gat));
  INV_X1    g539(.A(G99gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n723), .A2(new_n741), .A3(new_n644), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n725), .A2(new_n445), .A3(new_n726), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(G1338gat));
  NOR2_X1   g543(.A1(new_n438), .A2(G106gat), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n709), .A2(new_n722), .A3(new_n597), .A4(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n410), .B(new_n731), .C1(new_n661), .C2(new_n664), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G106gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n750), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n746), .A2(new_n752), .A3(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1339gat));
  NAND2_X1  g553(.A1(new_n684), .A2(new_n683), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT115), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n588), .A2(new_n590), .ZN(new_n757));
  INV_X1    g556(.A(new_n584), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n760), .A3(new_n579), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT54), .B1(new_n591), .B2(new_n580), .ZN(new_n762));
  AOI211_X1 g561(.A(new_n579), .B(new_n584), .C1(new_n588), .C2(new_n590), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n761), .B(new_n528), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n579), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n591), .A2(new_n580), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n767), .A2(KEYINPUT54), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n528), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n580), .B1(new_n757), .B2(new_n758), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n760), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(KEYINPUT55), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n767), .A2(new_n581), .A3(new_n770), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n766), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n521), .A2(new_n520), .ZN(new_n776));
  INV_X1    g575(.A(new_n452), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n511), .A2(new_n513), .B1(new_n499), .B2(new_n498), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n776), .A2(new_n453), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n662), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n523), .A3(new_n773), .A4(new_n774), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n597), .A2(new_n779), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n662), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n617), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n756), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n636), .A3(new_n714), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n425), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(new_n305), .A3(new_n523), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n787), .A2(new_n425), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G113gat), .B1(new_n793), .B2(new_n524), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(G1340gat));
  NAND3_X1  g594(.A1(new_n790), .A2(new_n303), .A3(new_n597), .ZN(new_n796));
  OAI21_X1  g595(.A(G120gat), .B1(new_n793), .B2(new_n683), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1341gat));
  AOI21_X1  g597(.A(G127gat), .B1(new_n790), .B2(new_n704), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n617), .A2(new_n601), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n792), .B2(new_n800), .ZN(G1342gat));
  NOR2_X1   g600(.A1(new_n425), .A2(new_n653), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(G134gat), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT56), .B1(new_n789), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n787), .A2(new_n788), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n787), .A2(new_n788), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n804), .ZN(new_n811));
  OAI21_X1  g610(.A(G134gat), .B1(new_n793), .B2(new_n653), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n806), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n806), .A2(new_n811), .A3(KEYINPUT117), .A4(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1343gat));
  NAND2_X1  g616(.A1(new_n786), .A2(new_n410), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n646), .A2(new_n635), .A3(new_n425), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OR3_X1    g620(.A1(new_n821), .A2(G141gat), .A3(new_n524), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n820), .B1(new_n818), .B2(KEYINPUT57), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n782), .A2(new_n783), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n632), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n782), .A2(new_n783), .A3(KEYINPUT118), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n704), .B1(new_n830), .B2(new_n780), .ZN(new_n831));
  INV_X1    g630(.A(new_n756), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n410), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n825), .B1(KEYINPUT57), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n225), .B1(new_n834), .B2(new_n523), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n821), .A2(G141gat), .A3(new_n524), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n824), .B(KEYINPUT58), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT58), .B1(new_n836), .B2(KEYINPUT119), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n834), .A2(new_n523), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n838), .B(new_n822), .C1(new_n839), .C2(new_n225), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(G1344gat));
  INV_X1    g640(.A(new_n821), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n222), .A3(new_n597), .ZN(new_n843));
  AOI211_X1 g642(.A(KEYINPUT59), .B(new_n222), .C1(new_n834), .C2(new_n597), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n775), .A2(new_n632), .A3(new_n779), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n828), .B2(new_n829), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n617), .B1(new_n847), .B2(KEYINPUT120), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n782), .A2(KEYINPUT118), .A3(new_n783), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT118), .B1(new_n782), .B2(new_n783), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n849), .A2(new_n850), .A3(new_n632), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(new_n846), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n755), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n438), .A2(KEYINPUT57), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n818), .A2(KEYINPUT57), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n856), .A2(new_n597), .A3(new_n820), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n845), .B1(new_n858), .B2(G148gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(new_n859), .ZN(G1345gat));
  AOI21_X1  g659(.A(new_n215), .B1(new_n842), .B2(new_n704), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n617), .A2(new_n216), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n834), .B2(new_n862), .ZN(G1346gat));
  AND2_X1   g662(.A1(new_n834), .A2(new_n662), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n445), .A2(new_n217), .A3(new_n636), .A4(new_n802), .ZN(new_n865));
  OAI22_X1  g664(.A1(new_n864), .A2(new_n217), .B1(new_n818), .B2(new_n865), .ZN(G1347gat));
  AOI21_X1  g665(.A(new_n636), .B1(new_n756), .B2(new_n785), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n338), .A2(new_n370), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(KEYINPUT122), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(KEYINPUT122), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873), .B2(new_n524), .ZN(new_n874));
  XOR2_X1   g673(.A(new_n868), .B(KEYINPUT121), .Z(new_n875));
  AND2_X1   g674(.A1(new_n867), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n289), .A3(new_n523), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n876), .B2(new_n597), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n683), .A2(new_n290), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n872), .B2(new_n880), .ZN(G1349gat));
  AOI21_X1  g680(.A(new_n605), .B1(new_n872), .B2(new_n704), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n617), .A2(new_n298), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n876), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT123), .Z(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n886), .B(KEYINPUT123), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT60), .B1(new_n882), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1350gat));
  INV_X1    g690(.A(G190gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n892), .A3(new_n662), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n872), .A2(new_n632), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(G190gat), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT61), .B(new_n892), .C1(new_n872), .C2(new_n632), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(G1351gat));
  NAND3_X1  g697(.A1(new_n445), .A2(new_n635), .A3(new_n425), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n818), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n449), .A3(new_n523), .ZN(new_n901));
  INV_X1    g700(.A(new_n855), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n852), .B1(new_n851), .B2(new_n846), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n847), .A2(KEYINPUT120), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n904), .A3(new_n617), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n905), .B2(new_n755), .ZN(new_n906));
  INV_X1    g705(.A(new_n857), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n906), .A2(new_n907), .A3(new_n899), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(new_n523), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n901), .B1(new_n909), .B2(new_n449), .ZN(G1352gat));
  XOR2_X1   g709(.A(KEYINPUT124), .B(G204gat), .Z(new_n911));
  AND2_X1   g710(.A1(new_n597), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n900), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT125), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT62), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT62), .B1(new_n914), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR4_X1   g718(.A1(new_n906), .A2(new_n907), .A3(new_n683), .A4(new_n899), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n911), .B2(new_n920), .ZN(G1353gat));
  INV_X1    g720(.A(new_n899), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n856), .A2(new_n704), .A3(new_n857), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT126), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(G211gat), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n923), .A2(new_n929), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n925), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n900), .A2(new_n205), .A3(new_n704), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1354gat));
  AOI21_X1  g732(.A(G218gat), .B1(new_n900), .B2(new_n662), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n632), .A2(G218gat), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT127), .Z(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n908), .B2(new_n936), .ZN(G1355gat));
endmodule


