//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT66), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT67), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(G101), .A2(new_n472), .B1(new_n473), .B2(G137), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n467), .A2(new_n475), .A3(G2105), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(new_n470), .B2(G112), .ZN(new_n478));
  INV_X1    g053(.A(G100), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(new_n470), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT68), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n465), .A2(new_n470), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n473), .A2(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .A3(G138), .ZN(new_n488));
  NAND2_X1  g063(.A1(G102), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n487), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT4), .B1(new_n491), .B2(new_n470), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n473), .A2(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(G543), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT5), .B1(new_n495), .B2(KEYINPUT69), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT69), .B1(new_n495), .B2(KEYINPUT70), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(KEYINPUT69), .B(KEYINPUT5), .C1(new_n495), .C2(KEYINPUT70), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(G543), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n502), .A2(G88), .B1(G50), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n498), .A2(new_n499), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  AOI22_X1  g089(.A1(new_n500), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n515), .A2(new_n509), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n518), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n516), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G168));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(G543), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n529), .B2(G543), .ZN(new_n530));
  OAI211_X1 g105(.A(G64), .B(new_n499), .C1(new_n528), .C2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n532), .B1(new_n531), .B2(new_n533), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n520), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n501), .B2(new_n539), .ZN(new_n540));
  NOR3_X1   g115(.A1(new_n537), .A2(KEYINPUT73), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n531), .A2(new_n533), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT72), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(G651), .A3(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n502), .A2(G90), .B1(new_n520), .B2(G52), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n541), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND3_X1  g125(.A1(new_n498), .A2(G56), .A3(new_n499), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n518), .B1(new_n500), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n519), .ZN(new_n556));
  OAI21_X1  g131(.A(G43), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT74), .B(G81), .Z(new_n558));
  NAND4_X1  g133(.A1(new_n498), .A2(new_n558), .A3(new_n499), .A4(new_n500), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n554), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  NAND3_X1  g142(.A1(new_n498), .A2(G65), .A3(new_n499), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n536), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n501), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g149(.A(G53), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n576), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n500), .A2(KEYINPUT75), .A3(G53), .A4(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT9), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n571), .A2(new_n574), .A3(new_n578), .A4(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n524), .A2(KEYINPUT76), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n516), .A2(new_n521), .A3(new_n584), .A4(new_n523), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(G286));
  NAND2_X1  g161(.A1(new_n506), .A2(G49), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n498), .A2(G87), .A3(new_n499), .A4(new_n500), .ZN(new_n588));
  AOI21_X1  g163(.A(G74), .B1(new_n498), .B2(new_n499), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(new_n536), .ZN(G288));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n509), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n502), .A2(G86), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n506), .A2(G48), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n520), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n501), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n498), .A2(G60), .A3(new_n499), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n536), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n509), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n498), .A2(G92), .A3(new_n499), .A4(new_n500), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(KEYINPUT10), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(KEYINPUT10), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G171), .B2(new_n614), .ZN(G284));
  OAI21_X1  g191(.A(new_n615), .B1(G171), .B2(new_n614), .ZN(G321));
  NAND2_X1  g192(.A1(G299), .A2(new_n614), .ZN(new_n618));
  INV_X1    g193(.A(G286), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n614), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n614), .ZN(G280));
  INV_X1    g196(.A(new_n613), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n560), .A2(new_n614), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n613), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g203(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT78), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n472), .A2(new_n487), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n482), .A2(G123), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n473), .A2(G135), .ZN(new_n639));
  OR2_X1    g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n640), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n482), .A2(KEYINPUT80), .A3(G123), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n638), .A2(new_n639), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n635), .A2(new_n644), .ZN(G156));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2438), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2430), .Z(new_n648));
  OAI21_X1  g223(.A(KEYINPUT14), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT81), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  AOI21_X1  g246(.A(KEYINPUT18), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n669), .B(new_n672), .Z(G227));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n675), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n677), .A2(new_n679), .A3(new_n681), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n684), .B(new_n685), .C1(new_n683), .C2(new_n682), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT82), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(G160), .A2(G29), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT24), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G34), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT94), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(G34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(KEYINPUT94), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G2084), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n705), .A2(KEYINPUT23), .A3(G20), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT23), .ZN(new_n707));
  INV_X1    g282(.A(G20), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n581), .A2(new_n578), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n710), .A2(new_n570), .A3(new_n573), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n706), .B(new_n709), .C1(new_n711), .C2(new_n705), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1956), .ZN(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  NAND2_X1  g289(.A1(G168), .A2(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G16), .B2(G21), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n704), .B(new_n713), .C1(new_n714), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n561), .A2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G16), .B2(G19), .ZN(new_n719));
  INV_X1    g294(.A(G1341), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n622), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G4), .B2(G16), .ZN(new_n723));
  INV_X1    g298(.A(G1348), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G5), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G171), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n721), .B(new_n725), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT84), .ZN(new_n732));
  INV_X1    g307(.A(G24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G16), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(G16), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G290), .B2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(new_n736), .B2(new_n732), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G1986), .ZN(new_n738));
  INV_X1    g313(.A(G1986), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n739), .B(new_n734), .C1(new_n736), .C2(new_n732), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n482), .A2(G119), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n473), .A2(G131), .ZN(new_n742));
  NOR2_X1   g317(.A1(G95), .A2(G2105), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(new_n470), .B2(G107), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT83), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n695), .A2(G25), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n745), .A2(G29), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT35), .B(G1991), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n749), .B(new_n750), .Z(new_n751));
  NAND3_X1  g326(.A1(new_n738), .A2(new_n740), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n753));
  NOR2_X1   g328(.A1(G16), .A2(G23), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT85), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G288), .B2(new_n705), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT86), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT33), .B(G1976), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n705), .A2(G6), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G305), .B2(G16), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT32), .B(G1981), .Z(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n705), .A2(G22), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G303), .B2(G16), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT87), .B(G1971), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT88), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n762), .A2(new_n763), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n764), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n753), .B1(new_n760), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n772), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n774), .A2(KEYINPUT34), .A3(new_n759), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n752), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI211_X1 g353(.A(KEYINPUT36), .B(new_n752), .C1(new_n773), .C2(new_n775), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n717), .B(new_n731), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n473), .A2(G141), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT95), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n472), .A2(G105), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT26), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n482), .A2(G129), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n782), .A2(new_n783), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G29), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G29), .B2(G32), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT27), .B(G1996), .ZN(new_n792));
  AND3_X1   g367(.A1(new_n791), .A2(KEYINPUT97), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(KEYINPUT97), .B1(new_n791), .B2(new_n792), .ZN(new_n794));
  NOR2_X1   g369(.A1(G164), .A2(new_n695), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n695), .A2(G27), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT99), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(KEYINPUT99), .B2(new_n796), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2078), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n793), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n719), .A2(new_n720), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n702), .A2(new_n703), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT98), .Z(new_n803));
  NOR4_X1   g378(.A1(new_n780), .A2(new_n800), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n487), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n470), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT93), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G139), .B2(new_n473), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT25), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G33), .B(new_n811), .S(G29), .Z(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G2072), .Z(new_n813));
  XOR2_X1   g388(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n695), .A2(G26), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n482), .A2(G128), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT89), .ZN(new_n818));
  NOR2_X1   g393(.A1(G104), .A2(G2105), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT90), .Z(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(new_n470), .B2(G116), .ZN(new_n821));
  INV_X1    g396(.A(G140), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n487), .A2(new_n470), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n816), .B1(new_n826), .B2(new_n695), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT92), .B(G2067), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT30), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(G28), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(G28), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n831), .A2(new_n832), .A3(new_n695), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n829), .B(new_n833), .C1(new_n695), .C2(new_n643), .ZN(new_n834));
  INV_X1    g409(.A(G2090), .ZN(new_n835));
  INV_X1    g410(.A(G35), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT100), .B1(new_n836), .B2(G29), .ZN(new_n837));
  OR3_X1    g412(.A1(new_n836), .A2(KEYINPUT100), .A3(G29), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n837), .B(new_n838), .C1(G162), .C2(new_n695), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT29), .Z(new_n840));
  AOI21_X1  g415(.A(new_n834), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n791), .A2(new_n792), .ZN(new_n842));
  INV_X1    g417(.A(G11), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT31), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI221_X1 g420(.A(new_n845), .B1(KEYINPUT31), .B2(new_n843), .C1(new_n724), .C2(new_n723), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n804), .A2(new_n813), .A3(new_n841), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n840), .A2(new_n835), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n716), .A2(new_n714), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G311));
  AND3_X1   g426(.A1(new_n804), .A2(new_n841), .A3(new_n847), .ZN(new_n852));
  INV_X1    g427(.A(new_n849), .ZN(new_n853));
  INV_X1    g428(.A(new_n850), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n813), .ZN(G150));
  OAI211_X1 g430(.A(G67), .B(new_n499), .C1(new_n528), .C2(new_n530), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G651), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n502), .A2(G93), .B1(new_n520), .B2(G55), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(KEYINPUT101), .A3(G651), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT103), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n622), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT38), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT39), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n864), .A2(KEYINPUT102), .A3(new_n560), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n557), .A2(new_n559), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n536), .B1(new_n551), .B2(new_n552), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT102), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT101), .B1(new_n858), .B2(G651), .ZN(new_n875));
  AOI211_X1 g450(.A(new_n860), .B(new_n536), .C1(new_n856), .C2(new_n857), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n554), .A2(new_n878), .A3(new_n557), .A4(new_n559), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n874), .A2(new_n877), .A3(new_n879), .A4(new_n862), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n870), .B(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n867), .B1(new_n882), .B2(G860), .ZN(G145));
  XNOR2_X1  g458(.A(G160), .B(new_n485), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n643), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n632), .B(new_n745), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n482), .A2(G130), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n473), .A2(G142), .ZN(new_n888));
  NOR2_X1   g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(new_n470), .B2(G118), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n886), .B(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n811), .A2(G164), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n462), .A2(new_n464), .A3(G126), .ZN(new_n894));
  NAND2_X1  g469(.A1(G114), .A2(G2104), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n470), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT4), .ZN(new_n897));
  INV_X1    g472(.A(G138), .ZN(new_n898));
  OAI22_X1  g473(.A1(new_n896), .A2(new_n897), .B1(new_n898), .B2(new_n823), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n488), .A2(new_n489), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n470), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n808), .B2(new_n810), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n893), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n787), .B(KEYINPUT96), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n825), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n826), .A3(new_n906), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n892), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n885), .B1(new_n912), .B2(KEYINPUT104), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n911), .A3(new_n892), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n913), .B1(new_n916), .B2(KEYINPUT104), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n915), .A3(new_n885), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g496(.A1(new_n864), .A2(new_n614), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n881), .B(KEYINPUT105), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(new_n626), .ZN(new_n924));
  NAND4_X1  g499(.A1(G299), .A2(new_n609), .A3(new_n611), .A4(new_n612), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n613), .A2(new_n711), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n924), .A2(KEYINPUT106), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT107), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n613), .A2(new_n931), .A3(new_n711), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n929), .B1(new_n933), .B2(KEYINPUT41), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT106), .B1(new_n924), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n924), .A2(new_n927), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n928), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G288), .B1(new_n507), .B2(new_n512), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n507), .A2(new_n512), .A3(G288), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(G305), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G305), .ZN(new_n943));
  INV_X1    g518(.A(new_n941), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n943), .B1(new_n944), .B2(new_n939), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n945), .A3(new_n604), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n604), .B1(new_n942), .B2(new_n945), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT42), .ZN(new_n949));
  INV_X1    g524(.A(new_n948), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n946), .A3(KEYINPUT108), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n947), .B2(new_n948), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n949), .B1(new_n954), .B2(KEYINPUT42), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n938), .B(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n922), .B1(new_n956), .B2(new_n614), .ZN(G295));
  OAI21_X1  g532(.A(new_n922), .B1(new_n956), .B2(new_n614), .ZN(G331));
  NOR3_X1   g533(.A1(new_n541), .A2(new_n548), .A3(new_n524), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT73), .B1(new_n537), .B2(new_n540), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n546), .A2(new_n542), .A3(new_n547), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n960), .A2(new_n961), .B1(new_n583), .B2(new_n585), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n881), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n964));
  OAI21_X1  g539(.A(G286), .B1(new_n541), .B2(new_n548), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n871), .A2(new_n880), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n960), .A2(G168), .A3(new_n961), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n963), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n966), .A2(new_n965), .A3(KEYINPUT109), .A4(new_n967), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n970), .A3(new_n934), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n963), .A2(new_n927), .A3(new_n968), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n954), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n918), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n954), .B1(new_n971), .B2(new_n972), .ZN(new_n975));
  OR3_X1    g550(.A1(new_n974), .A2(KEYINPUT43), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n969), .A2(new_n970), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n930), .A2(KEYINPUT41), .A3(new_n932), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n968), .B2(new_n963), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n927), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(KEYINPUT41), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n954), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT43), .B1(new_n982), .B2(new_n974), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n976), .A2(KEYINPUT44), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n974), .B2(new_n975), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n982), .A2(new_n974), .A3(KEYINPUT43), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n986), .A2(new_n988), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n985), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI211_X1 g568(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n989), .C2(new_n990), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n984), .B1(new_n993), .B2(new_n994), .ZN(G397));
  INV_X1    g570(.A(KEYINPUT126), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(G164), .B2(G1384), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n899), .B2(new_n901), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT45), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n469), .A2(new_n474), .A3(G40), .A4(new_n476), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n714), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1000), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT50), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1000), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1007), .A2(new_n703), .A3(new_n1003), .A4(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n997), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT115), .B(G8), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G168), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT51), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1015), .A2(KEYINPUT51), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT124), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT124), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1000), .A2(new_n1022), .ZN(new_n1023));
  AOI211_X1 g598(.A(G1384), .B(new_n1008), .C1(new_n899), .C2(new_n901), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n1002), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1025), .A2(new_n703), .B1(new_n1004), .B2(new_n714), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1021), .B(new_n1018), .C1(new_n1026), .C2(new_n1014), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1016), .A2(new_n1020), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1017), .A2(new_n524), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1031));
  INV_X1    g606(.A(G1971), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1004), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1004), .A2(KEYINPUT112), .A3(new_n1032), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1007), .A2(new_n1003), .A3(new_n1010), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1035), .B(new_n1036), .C1(G2090), .C2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1039), .A2(KEYINPUT114), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(G166), .B2(new_n997), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(KEYINPUT114), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1038), .A2(G8), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1006), .A2(new_n1002), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(new_n1014), .ZN(new_n1047));
  INV_X1    g622(.A(G288), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT116), .B(G1976), .Z(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT117), .B1(new_n1048), .B2(G1976), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1047), .B(new_n1052), .C1(KEYINPUT52), .C2(new_n1050), .ZN(new_n1055));
  OR2_X1    g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G305), .A2(G1981), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT49), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT49), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1054), .A2(new_n1055), .B1(new_n1060), .B2(new_n1047), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1044), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1000), .A2(new_n1022), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1003), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1000), .A2(new_n1009), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1064), .A2(G2090), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1032), .B2(new_n1004), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1067), .B2(new_n1014), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1045), .A2(new_n1061), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1037), .A2(new_n728), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1004), .B2(G2078), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n999), .A2(new_n1001), .ZN(new_n1074));
  INV_X1    g649(.A(G2078), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(KEYINPUT53), .A3(new_n1075), .A4(new_n1003), .ZN(new_n1076));
  AOI21_X1  g651(.A(G301), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1028), .A2(new_n1078), .A3(new_n1029), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1031), .A2(new_n1069), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1017), .A2(new_n619), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1038), .A2(G8), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1062), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(KEYINPUT63), .A3(new_n1045), .A4(new_n1061), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1081), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1045), .A2(new_n1061), .A3(new_n1068), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1061), .A2(G8), .A3(new_n1044), .A4(new_n1038), .ZN(new_n1090));
  AOI21_X1  g665(.A(G1976), .B1(new_n1060), .B2(new_n1047), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1048), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1056), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1047), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1080), .A2(new_n1089), .A3(new_n1090), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G2067), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1037), .A2(new_n724), .B1(new_n1097), .B2(new_n1046), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n613), .ZN(new_n1099));
  NAND2_X1  g674(.A1(G299), .A2(KEYINPUT118), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n570), .A2(new_n573), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n581), .A2(new_n578), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(KEYINPUT57), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1103), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1107));
  NOR4_X1   g682(.A1(new_n710), .A2(new_n570), .A3(new_n573), .A4(KEYINPUT118), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT119), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1105), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G1956), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1099), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1116), .A2(new_n1105), .A3(new_n1109), .A4(new_n1118), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT120), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1120), .A2(KEYINPUT120), .A3(new_n1122), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1118), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1002), .B1(new_n1022), .B2(new_n1000), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1956), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1110), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1130), .A3(new_n1121), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1119), .A2(KEYINPUT122), .A3(new_n1110), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1131), .A2(KEYINPUT123), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1113), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1112), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1119), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1121), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1098), .A2(new_n613), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT60), .B1(new_n1143), .B2(new_n1099), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT58), .B(G1341), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1004), .A2(G1996), .B1(new_n1046), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n561), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(KEYINPUT121), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1147), .B(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1098), .A2(new_n1151), .A3(new_n622), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1142), .A2(new_n1144), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1123), .B(new_n1124), .C1(new_n1138), .C2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n474), .A2(KEYINPUT53), .A3(new_n1075), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1074), .A2(G40), .A3(new_n468), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1073), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(G171), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1073), .A2(G301), .A3(new_n1076), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1160), .A2(KEYINPUT54), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1069), .A2(new_n1030), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1157), .A2(G171), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n1077), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1154), .A2(new_n1163), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n999), .A2(new_n1002), .ZN(new_n1169));
  INV_X1    g744(.A(G1996), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n789), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n905), .A2(G1996), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n825), .B(new_n1097), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n745), .A2(new_n750), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n745), .A2(new_n750), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(G290), .A2(G1986), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n604), .A2(new_n739), .ZN(new_n1181));
  OR3_X1    g756(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1096), .A2(new_n1168), .B1(new_n1169), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1169), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1180), .A2(new_n1169), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT48), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1169), .B1(new_n1174), .B2(new_n905), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT46), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1169), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(G1996), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1169), .A2(KEYINPUT46), .A3(new_n1170), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1188), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT47), .ZN(new_n1194));
  AOI22_X1  g769(.A1(new_n1175), .A2(new_n1178), .B1(new_n1097), .B2(new_n826), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1195), .A2(new_n1190), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1187), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n996), .B1(new_n1183), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1182), .A2(new_n1169), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1168), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1199), .B1(new_n1200), .B2(new_n1095), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1197), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1201), .A2(KEYINPUT126), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1198), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g779(.A(G227), .ZN(new_n1206));
  NOR2_X1   g780(.A1(G229), .A2(new_n458), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n660), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1208), .A2(KEYINPUT127), .ZN(new_n1209));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n1210));
  NAND4_X1  g784(.A1(new_n660), .A2(new_n1210), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1211));
  NAND4_X1  g785(.A1(new_n920), .A2(new_n991), .A3(new_n1209), .A4(new_n1211), .ZN(G225));
  INV_X1    g786(.A(G225), .ZN(G308));
endmodule


