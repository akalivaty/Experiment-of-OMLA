//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n641, new_n642, new_n643, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n463), .B1(new_n471), .B2(G2105), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G137), .A3(new_n462), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G137), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n473), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NOR3_X1   g061(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G112), .B2(new_n462), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n476), .A2(G136), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n473), .A2(G126), .A3(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n473), .A2(new_n462), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n497), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n476), .B(new_n500), .C1(new_n496), .C2(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n495), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT71), .B1(new_n506), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT6), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(new_n510), .B1(new_n506), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n511), .A2(G88), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n511), .A2(G50), .A3(G543), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n514), .B2(new_n515), .ZN(new_n520));
  AND2_X1   g095(.A1(G75), .A2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(G651), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n517), .A2(new_n518), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  AOI21_X1  g099(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n528), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n525), .A2(G63), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n507), .A2(new_n510), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n506), .A2(G651), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n531), .A2(G89), .A3(new_n532), .A4(new_n516), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n531), .A2(G51), .A3(G543), .A4(new_n532), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n509), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT72), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n511), .A2(G52), .A3(G543), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n531), .A2(new_n532), .A3(new_n516), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n539), .A2(new_n543), .ZN(G171));
  NAND3_X1  g119(.A1(new_n511), .A2(G81), .A3(new_n516), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n531), .A2(G43), .A3(G543), .A4(new_n532), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n514), .B2(new_n515), .ZN(new_n548));
  AND2_X1   g123(.A1(G68), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n554));
  XOR2_X1   g129(.A(new_n554), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  AND2_X1   g133(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  AND3_X1   g135(.A1(KEYINPUT75), .A2(G53), .A3(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n560), .B1(new_n511), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(G53), .A2(G543), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n559), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n565), .A2(new_n531), .A3(new_n532), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT76), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n531), .A2(new_n532), .A3(new_n561), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(new_n559), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n511), .A2(new_n565), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n542), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n515), .ZN(new_n576));
  NOR2_X1   g151(.A1(KEYINPUT5), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  NOR3_X1   g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT77), .B1(new_n514), .B2(new_n515), .ZN(new_n580));
  OAI21_X1  g155(.A(G65), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n575), .B1(new_n583), .B2(G651), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n573), .A2(KEYINPUT78), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT78), .B1(new_n573), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(G299));
  INV_X1    g162(.A(G171), .ZN(G301));
  NAND2_X1  g163(.A1(new_n516), .A2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(G74), .A2(G651), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n589), .A2(KEYINPUT79), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n592), .B(G651), .C1(new_n516), .C2(G74), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n511), .A2(G87), .A3(new_n516), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n511), .A2(G49), .A3(G543), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n514), .B2(new_n515), .ZN(new_n599));
  AND2_X1   g174(.A1(G73), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n531), .A2(G48), .A3(G543), .A4(new_n532), .ZN(new_n602));
  INV_X1    g177(.A(G86), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(new_n602), .C1(new_n542), .C2(new_n603), .ZN(G305));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n514), .B2(new_n515), .ZN(new_n606));
  AND2_X1   g181(.A1(G72), .A2(G543), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n531), .A2(G47), .A3(G543), .A4(new_n532), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n608), .B(new_n609), .C1(new_n542), .C2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n511), .A2(G92), .A3(new_n516), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n578), .B1(new_n576), .B2(new_n577), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n514), .A2(KEYINPUT77), .A3(new_n515), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(G651), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n511), .A2(G54), .A3(G543), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n622), .A2(KEYINPUT80), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(KEYINPUT80), .B1(new_n622), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n615), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT81), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n613), .B(KEYINPUT10), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n629));
  OAI21_X1  g204(.A(G66), .B1(new_n579), .B2(new_n580), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n509), .B1(new_n630), .B2(new_n620), .ZN(new_n631));
  INV_X1    g206(.A(new_n623), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n622), .A2(KEYINPUT80), .A3(new_n623), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n628), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n627), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n612), .B1(new_n638), .B2(G868), .ZN(G284));
  OAI21_X1  g214(.A(new_n612), .B1(new_n638), .B2(G868), .ZN(G321));
  NAND2_X1  g215(.A1(G286), .A2(G868), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT82), .ZN(new_n642));
  INV_X1    g217(.A(G299), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(G868), .ZN(G297));
  OAI21_X1  g219(.A(new_n642), .B1(new_n643), .B2(G868), .ZN(G280));
  INV_X1    g220(.A(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n638), .B1(new_n646), .B2(G860), .ZN(G148));
  INV_X1    g222(.A(G868), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n551), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n627), .A2(new_n637), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n650), .A2(G559), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n649), .B1(new_n651), .B2(new_n648), .ZN(G323));
  XNOR2_X1  g227(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g228(.A1(new_n476), .A2(G135), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n462), .A2(G111), .ZN(new_n655));
  OAI21_X1  g230(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n656));
  INV_X1    g231(.A(G123), .ZN(new_n657));
  OAI221_X1 g232(.A(new_n654), .B1(new_n655), .B2(new_n656), .C1(new_n657), .C2(new_n482), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT83), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT12), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT13), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n664), .ZN(G156));
  XNOR2_X1  g240(.A(KEYINPUT15), .B(G2435), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2438), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2427), .B(G2430), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT14), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n667), .B2(new_n668), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1341), .B(G1348), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2451), .B(G2454), .Z(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2443), .B(G2446), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(G14), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n678), .ZN(G401));
  XOR2_X1   g257(.A(G2084), .B(G2090), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT86), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n686), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(KEYINPUT17), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G2072), .B(G2078), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n692), .B(new_n693), .C1(new_n691), .C2(new_n687), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n692), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g270(.A(G2096), .B(G2100), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G227));
  XOR2_X1   g272(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n698));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1956), .B(G2474), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1961), .B(G1966), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT20), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n701), .A2(new_n702), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n703), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n705), .B(new_n707), .C1(new_n700), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(G1991), .B(G1996), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1981), .B(G1986), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(G229));
  INV_X1    g292(.A(KEYINPUT94), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n719));
  NAND2_X1  g294(.A1(G288), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n594), .A2(KEYINPUT92), .A3(new_n595), .A4(new_n596), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G23), .B(new_n722), .S(G16), .Z(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT33), .B(G1976), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G6), .B(G305), .S(G16), .Z(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT32), .B(G1981), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G22), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G166), .B2(new_n732), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1971), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n728), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n726), .B1(new_n724), .B2(new_n727), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n718), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n738), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n740), .A2(new_n728), .A3(KEYINPUT94), .A4(new_n736), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n739), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT89), .B(G29), .Z(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(G25), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n476), .A2(G131), .ZN(new_n748));
  OR2_X1    g323(.A1(G95), .A2(G2105), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n749), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n750));
  INV_X1    g325(.A(G119), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n750), .C1(new_n751), .C2(new_n482), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n747), .B1(new_n753), .B2(new_n746), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT90), .Z(new_n755));
  XOR2_X1   g330(.A(KEYINPUT35), .B(G1991), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G24), .B(G290), .S(G16), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1986), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n744), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n743), .B1(new_n739), .B2(new_n741), .ZN(new_n762));
  OAI21_X1  g337(.A(KEYINPUT36), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n739), .A2(new_n741), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(new_n742), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT36), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n765), .A2(new_n766), .A3(new_n744), .A4(new_n760), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n746), .A2(G35), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n746), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT29), .B(G2090), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT31), .B(G11), .Z(new_n773));
  INV_X1    g348(.A(G29), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G28), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(KEYINPUT100), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n776), .A2(KEYINPUT100), .B1(new_n775), .B2(G28), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n658), .B2(new_n745), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n771), .A2(new_n772), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G1966), .ZN(new_n782));
  NOR2_X1   g357(.A1(G168), .A2(new_n732), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n732), .B2(G21), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n781), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n774), .A2(G33), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT25), .Z(new_n788));
  INV_X1    g363(.A(G139), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n498), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(new_n462), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT98), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n786), .B1(new_n797), .B2(new_n774), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G2072), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n732), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n732), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(G1961), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n785), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n483), .A2(G129), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n476), .A2(G141), .ZN(new_n806));
  NAND3_X1  g381(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT26), .Z(new_n808));
  NAND4_X1  g383(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G32), .B(new_n809), .S(G29), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT99), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT27), .B(G1996), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G2072), .B2(new_n798), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT24), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G34), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(G34), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n745), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n480), .B2(new_n774), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G2084), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n746), .A2(G27), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G164), .B2(new_n746), .ZN(new_n822));
  INV_X1    g397(.A(G2078), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n782), .B2(new_n784), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n811), .A2(new_n812), .B1(G1961), .B2(new_n801), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n803), .A2(new_n814), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(G299), .A2(G16), .ZN(new_n830));
  INV_X1    g405(.A(G1956), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n732), .A2(G20), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT101), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT23), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n831), .B1(new_n830), .B2(new_n834), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n829), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n732), .A2(G4), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n650), .B2(G16), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT95), .B(G1348), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n732), .A2(G19), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n552), .B2(new_n732), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(G1341), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n476), .A2(G140), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n462), .A2(G116), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n848));
  INV_X1    g423(.A(G128), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n846), .B1(new_n847), .B2(new_n848), .C1(new_n849), .C2(new_n482), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G29), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n745), .A2(G26), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT28), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(G2067), .Z(new_n855));
  NAND4_X1  g430(.A1(new_n841), .A2(new_n842), .A3(new_n845), .A4(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n837), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT102), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n837), .A2(new_n859), .A3(new_n862), .A4(new_n858), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n763), .A2(new_n767), .B1(new_n861), .B2(new_n863), .ZN(G311));
  NAND2_X1  g439(.A1(new_n763), .A2(new_n767), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n863), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(G150));
  NAND2_X1  g442(.A1(new_n638), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT38), .ZN(new_n869));
  INV_X1    g444(.A(G67), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n514), .B2(new_n515), .ZN(new_n871));
  AND2_X1   g446(.A1(G80), .A2(G543), .ZN(new_n872));
  OAI21_X1  g447(.A(G651), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(KEYINPUT103), .B(G55), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n531), .A2(G543), .A3(new_n532), .A4(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n531), .A2(G93), .A3(new_n532), .A4(new_n516), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n551), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n551), .A2(new_n877), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n869), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n883));
  AOI21_X1  g458(.A(G860), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n883), .B2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n877), .A2(G860), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT37), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(G145));
  XNOR2_X1  g463(.A(new_n850), .B(KEYINPUT105), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n796), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n796), .A2(new_n889), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n752), .B(KEYINPUT106), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n662), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n502), .A2(KEYINPUT104), .A3(new_n503), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT104), .B1(new_n502), .B2(new_n503), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n495), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n809), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n476), .A2(G142), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n462), .A2(G118), .ZN(new_n904));
  OAI21_X1  g479(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n905));
  INV_X1    g480(.A(G130), .ZN(new_n906));
  OAI221_X1 g481(.A(new_n903), .B1(new_n904), .B2(new_n905), .C1(new_n906), .C2(new_n482), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n902), .B(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n898), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n896), .A2(new_n908), .A3(new_n897), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n490), .B(new_n658), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n480), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  INV_X1    g491(.A(new_n914), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n910), .A2(new_n917), .A3(new_n911), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n916), .A4(new_n918), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n921), .A2(KEYINPUT40), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT40), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(G395));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  OR2_X1    g502(.A1(G303), .A2(G305), .ZN(new_n928));
  NAND2_X1  g503(.A1(G303), .A2(G305), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(KEYINPUT110), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n931));
  AND2_X1   g506(.A1(G303), .A2(G305), .ZN(new_n932));
  NOR2_X1   g507(.A1(G303), .A2(G305), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  XNOR2_X1  g511(.A(G290), .B(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n720), .A3(new_n721), .ZN(new_n938));
  XNOR2_X1  g513(.A(G290), .B(KEYINPUT109), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n722), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n935), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n932), .A2(new_n933), .A3(new_n931), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n940), .A2(new_n938), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n927), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT111), .B1(new_n941), .B2(new_n943), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(new_n926), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n940), .A2(new_n938), .A3(new_n942), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n940), .A2(new_n938), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n947), .B(new_n948), .C1(new_n949), .C2(new_n935), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT42), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n944), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n952), .A2(KEYINPUT113), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n651), .A2(new_n881), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n880), .B1(new_n650), .B2(G559), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n626), .B1(new_n585), .B2(new_n586), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n562), .A2(new_n566), .A3(KEYINPUT76), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n584), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT78), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n573), .A2(KEYINPUT78), .A3(new_n584), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n635), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n954), .A2(new_n955), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n954), .A2(new_n955), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT41), .B1(new_n956), .B2(new_n963), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n956), .A2(new_n963), .A3(KEYINPUT41), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n965), .A2(new_n966), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n952), .A2(KEYINPUT113), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n953), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n953), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g551(.A(G868), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n877), .A2(new_n648), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(G295));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n978), .ZN(G331));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT114), .B(KEYINPUT44), .Z(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n945), .A2(new_n950), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n985));
  NAND2_X1  g560(.A1(G286), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n530), .A2(new_n533), .A3(new_n534), .A4(KEYINPUT115), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n986), .B(new_n987), .C1(new_n878), .C2(new_n879), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n987), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n551), .A2(new_n877), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n551), .A2(new_n877), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n988), .A2(new_n992), .A3(G171), .ZN(new_n993));
  AOI21_X1  g568(.A(G171), .B1(new_n988), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n964), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT41), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n585), .A2(new_n626), .A3(new_n586), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n635), .B1(new_n961), .B2(new_n962), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n956), .A2(new_n963), .A3(KEYINPUT41), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n995), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n996), .B1(new_n1002), .B2(KEYINPUT116), .ZN(new_n1003));
  INV_X1    g578(.A(new_n994), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n988), .A2(new_n992), .A3(G171), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT116), .B(new_n1006), .C1(new_n970), .C2(new_n969), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n984), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n964), .A2(new_n1005), .A3(new_n1004), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n984), .ZN(new_n1012));
  AOI21_X1  g587(.A(G37), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1009), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n984), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1006), .B1(new_n970), .B2(new_n969), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1017), .A2(new_n945), .A3(new_n950), .A4(new_n996), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n916), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n983), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1014), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1016), .A2(new_n1018), .A3(new_n1014), .A4(new_n916), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT44), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n981), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1010), .B1(new_n1017), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1012), .B1(new_n1028), .B2(new_n1007), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1018), .A2(new_n916), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1029), .A2(new_n1030), .A3(KEYINPUT43), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1014), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n982), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT43), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(KEYINPUT44), .A3(new_n1023), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(KEYINPUT117), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1026), .A2(new_n1036), .ZN(G397));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n1038));
  INV_X1    g613(.A(new_n495), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n502), .A2(new_n503), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT104), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n502), .A2(KEYINPUT104), .A3(new_n503), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1039), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1038), .B1(new_n1044), .B2(G1384), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n472), .A2(G40), .A3(new_n479), .ZN(new_n1046));
  OR3_X1    g621(.A1(new_n1045), .A2(KEYINPUT118), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT118), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n850), .B(G2067), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT120), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1053), .A3(new_n1050), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n809), .B(G1996), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n753), .A2(new_n756), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1057), .A2(new_n1058), .B1(G2067), .B2(new_n850), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1049), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT46), .ZN(new_n1062));
  OR3_X1    g637(.A1(new_n1061), .A2(new_n1062), .A3(G1996), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1049), .B1(new_n809), .B2(new_n1050), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1061), .B2(G1996), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT47), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1057), .ZN(new_n1068));
  XOR2_X1   g643(.A(new_n752), .B(new_n756), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n1049), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G290), .A2(G1986), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1049), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1072), .B(KEYINPUT48), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1060), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G8), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1044), .A2(G1384), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1046), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(G305), .B(G1981), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT122), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1080), .A2(KEYINPUT122), .A3(new_n1081), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1079), .B(new_n1082), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1976), .ZN(new_n1086));
  INV_X1    g661(.A(G288), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(G1981), .B2(G305), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1079), .B(KEYINPUT123), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n720), .A2(G1976), .A3(new_n721), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1079), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT52), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n1086), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1094), .B(KEYINPUT121), .Z(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n1079), .A3(new_n1091), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1093), .A2(new_n1085), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1038), .A2(G1384), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n901), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1384), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n504), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1046), .B1(new_n1101), .B2(new_n1038), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1971), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT50), .B1(new_n901), .B2(new_n1100), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT50), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1101), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1078), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1105), .B1(new_n1109), .B2(G2090), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G303), .A2(G8), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT55), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(G8), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1089), .A2(new_n1090), .B1(new_n1097), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1107), .B1(new_n901), .B2(new_n1100), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1078), .B1(new_n1101), .B2(KEYINPUT50), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(G2090), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1104), .B2(new_n1103), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1112), .B1(new_n1120), .B2(new_n1076), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT45), .B1(new_n901), .B2(new_n1100), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n504), .A2(new_n1098), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1078), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n782), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1046), .A2(G2084), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1076), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1128), .A2(G168), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1097), .A2(new_n1121), .A3(new_n1114), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(KEYINPUT63), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1093), .A2(new_n1096), .A3(new_n1085), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1113), .B1(new_n1110), .B2(G8), .ZN(new_n1135));
  NOR4_X1   g710(.A1(new_n1133), .A2(new_n1115), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1116), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1125), .A2(new_n1127), .A3(G168), .ZN(new_n1138));
  OAI21_X1  g713(.A(G8), .B1(KEYINPUT126), .B2(KEYINPUT51), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT51), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1138), .B(new_n1140), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1128), .A2(G286), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT62), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1099), .A2(new_n1102), .A3(new_n823), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(G2078), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1045), .A2(new_n1078), .A3(new_n1153), .A4(new_n1123), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1107), .B1(new_n1044), .B2(G1384), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1108), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1046), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1152), .B(new_n1154), .C1(new_n1157), .C2(G1961), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1158), .A2(new_n1159), .A3(G171), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1158), .B2(G171), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1141), .A2(new_n1144), .B1(G286), .B2(new_n1128), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n1146), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1149), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1158), .A2(G171), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT54), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1045), .A2(new_n1099), .A3(new_n1078), .A4(new_n1153), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1152), .B(new_n1169), .C1(new_n1157), .C2(G1961), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1170), .B2(G171), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1163), .A2(new_n1146), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1170), .A2(G171), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1160), .A2(new_n1161), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n1174), .B2(KEYINPUT54), .ZN(new_n1175));
  INV_X1    g750(.A(new_n840), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1157), .A2(new_n1176), .B1(new_n1177), .B2(G2067), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n831), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1179));
  INV_X1    g754(.A(new_n584), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT57), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(new_n562), .B2(new_n566), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1183), .B1(new_n959), .B2(KEYINPUT57), .ZN(new_n1184));
  XNOR2_X1  g759(.A(KEYINPUT56), .B(G2072), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1099), .A2(new_n1102), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1179), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1178), .A2(new_n635), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1184), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1177), .A2(G2067), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1193), .B1(new_n840), .B2(new_n1109), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT60), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1195), .B1(new_n635), .B2(KEYINPUT125), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n626), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1194), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  OAI211_X1 g774(.A(new_n1197), .B(new_n626), .C1(new_n1178), .C2(new_n1195), .ZN(new_n1200));
  OAI211_X1 g775(.A(new_n1199), .B(new_n1200), .C1(KEYINPUT60), .C2(new_n1194), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1187), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1184), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1203));
  OAI21_X1  g778(.A(KEYINPUT61), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1191), .A2(new_n1205), .A3(new_n1187), .ZN(new_n1206));
  XOR2_X1   g781(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n1207));
  INV_X1    g782(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1103), .A2(G1996), .ZN(new_n1209));
  XNOR2_X1  g784(.A(KEYINPUT58), .B(G1341), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1210), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n552), .B(new_n1208), .C1(new_n1209), .C2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n552), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n1207), .ZN(new_n1214));
  AOI22_X1  g789(.A1(new_n1204), .A2(new_n1206), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1192), .B1(new_n1201), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1166), .B1(new_n1175), .B2(new_n1216), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1097), .A2(new_n1121), .A3(new_n1114), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1137), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  AND2_X1   g794(.A1(G290), .A2(G1986), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1049), .B1(new_n1220), .B2(new_n1071), .ZN(new_n1221));
  XOR2_X1   g796(.A(new_n1221), .B(KEYINPUT119), .Z(new_n1222));
  NAND3_X1  g797(.A1(new_n1222), .A2(new_n1070), .A3(new_n1068), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1075), .B1(new_n1219), .B2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g799(.A1(new_n921), .A2(new_n922), .ZN(new_n1226));
  INV_X1    g800(.A(G319), .ZN(new_n1227));
  NOR2_X1   g801(.A1(G227), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g802(.A(new_n1228), .B1(new_n715), .B2(new_n716), .ZN(new_n1229));
  NOR2_X1   g803(.A1(G401), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g804(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1231));
  NAND3_X1  g805(.A1(new_n1226), .A2(new_n1230), .A3(new_n1231), .ZN(G225));
  INV_X1    g806(.A(G225), .ZN(G308));
endmodule


