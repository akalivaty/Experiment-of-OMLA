

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U549 ( .A1(n804), .A2(n803), .ZN(n817) );
  NOR2_X1 U550 ( .A1(G1384), .A2(G164), .ZN(n773) );
  INV_X1 U551 ( .A(KEYINPUT26), .ZN(n690) );
  INV_X1 U552 ( .A(KEYINPUT29), .ZN(n710) );
  NAND2_X1 U553 ( .A1(n773), .A2(n681), .ZN(n728) );
  XNOR2_X1 U554 ( .A(KEYINPUT12), .B(KEYINPUT68), .ZN(n569) );
  XNOR2_X1 U555 ( .A(n570), .B(n569), .ZN(n572) );
  NOR2_X2 U556 ( .A1(G2104), .A2(n516), .ZN(n844) );
  NOR2_X1 U557 ( .A1(G651), .A2(n646), .ZN(n640) );
  NOR2_X1 U558 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U559 ( .A1(n579), .A2(n578), .ZN(n965) );
  XNOR2_X1 U560 ( .A(n522), .B(KEYINPUT82), .ZN(G164) );
  AND2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n843) );
  NAND2_X1 U562 ( .A1(G114), .A2(n843), .ZN(n515) );
  INV_X1 U563 ( .A(G2105), .ZN(n516) );
  NAND2_X1 U564 ( .A1(G126), .A2(n844), .ZN(n514) );
  AND2_X1 U565 ( .A1(n515), .A2(n514), .ZN(n518) );
  AND2_X1 U566 ( .A1(n516), .A2(G2104), .ZN(n847) );
  NAND2_X1 U567 ( .A1(G102), .A2(n847), .ZN(n517) );
  AND2_X1 U568 ( .A1(n518), .A2(n517), .ZN(n521) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n519), .Z(n848) );
  NAND2_X1 U571 ( .A1(n848), .A2(G138), .ZN(n520) );
  AND2_X1 U572 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n523) );
  XOR2_X2 U574 ( .A(KEYINPUT65), .B(n523), .Z(n631) );
  NAND2_X1 U575 ( .A1(G85), .A2(n631), .ZN(n525) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n646) );
  INV_X1 U577 ( .A(G651), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n646), .A2(n526), .ZN(n634) );
  NAND2_X1 U579 ( .A1(G72), .A2(n634), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U581 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n527), .Z(n645) );
  NAND2_X1 U583 ( .A1(G60), .A2(n645), .ZN(n529) );
  NAND2_X1 U584 ( .A1(G47), .A2(n640), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n530) );
  OR2_X1 U586 ( .A1(n531), .A2(n530), .ZN(G290) );
  XOR2_X1 U587 ( .A(G2446), .B(G2451), .Z(n533) );
  XNOR2_X1 U588 ( .A(G2454), .B(KEYINPUT97), .ZN(n532) );
  XNOR2_X1 U589 ( .A(n533), .B(n532), .ZN(n540) );
  XOR2_X1 U590 ( .A(G2438), .B(G2430), .Z(n535) );
  XNOR2_X1 U591 ( .A(G2435), .B(G2443), .ZN(n534) );
  XNOR2_X1 U592 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U593 ( .A(n536), .B(G2427), .Z(n538) );
  XNOR2_X1 U594 ( .A(G1341), .B(G1348), .ZN(n537) );
  XNOR2_X1 U595 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U596 ( .A(n540), .B(n539), .ZN(n541) );
  AND2_X1 U597 ( .A1(n541), .A2(G14), .ZN(G401) );
  XNOR2_X1 U598 ( .A(KEYINPUT9), .B(KEYINPUT67), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G90), .A2(n631), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G77), .A2(n634), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n545), .B(n544), .ZN(n550) );
  NAND2_X1 U603 ( .A1(n645), .A2(G64), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n546), .B(KEYINPUT66), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G52), .A2(n640), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n550), .A2(n549), .ZN(G171) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  NAND2_X1 U612 ( .A1(G65), .A2(n645), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G53), .A2(n640), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G91), .A2(n631), .ZN(n554) );
  NAND2_X1 U616 ( .A1(G78), .A2(n634), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n705) );
  INV_X1 U619 ( .A(n705), .ZN(G299) );
  NAND2_X1 U620 ( .A1(n631), .A2(G89), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G76), .A2(n634), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(KEYINPUT5), .ZN(n565) );
  NAND2_X1 U625 ( .A1(G63), .A2(n645), .ZN(n562) );
  NAND2_X1 U626 ( .A1(G51), .A2(n640), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n566), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n820) );
  NAND2_X1 U635 ( .A1(n820), .A2(G567), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  XNOR2_X1 U637 ( .A(KEYINPUT13), .B(KEYINPUT69), .ZN(n574) );
  NAND2_X1 U638 ( .A1(G81), .A2(n631), .ZN(n570) );
  NAND2_X1 U639 ( .A1(G68), .A2(n634), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n645), .A2(G56), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(n575), .Z(n576) );
  NAND2_X1 U644 ( .A1(n640), .A2(G43), .ZN(n578) );
  INV_X1 U645 ( .A(G860), .ZN(n616) );
  OR2_X1 U646 ( .A1(n965), .A2(n616), .ZN(G153) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  INV_X1 U648 ( .A(G868), .ZN(n594) );
  NOR2_X1 U649 ( .A1(G301), .A2(n594), .ZN(n593) );
  INV_X1 U650 ( .A(KEYINPUT15), .ZN(n590) );
  NAND2_X1 U651 ( .A1(G79), .A2(n634), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G54), .A2(n640), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n631), .A2(G92), .ZN(n582) );
  XNOR2_X1 U655 ( .A(n582), .B(KEYINPUT70), .ZN(n584) );
  NAND2_X1 U656 ( .A1(G66), .A2(n645), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n586) );
  INV_X1 U658 ( .A(KEYINPUT71), .ZN(n585) );
  XNOR2_X1 U659 ( .A(n586), .B(n585), .ZN(n587) );
  NOR2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U661 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U662 ( .A(KEYINPUT72), .B(n591), .ZN(n959) );
  INV_X1 U663 ( .A(n959), .ZN(n871) );
  NOR2_X1 U664 ( .A1(n871), .A2(G868), .ZN(n592) );
  NOR2_X1 U665 ( .A1(n593), .A2(n592), .ZN(G284) );
  NOR2_X1 U666 ( .A1(G286), .A2(n594), .ZN(n596) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U669 ( .A1(G559), .A2(n616), .ZN(n597) );
  XOR2_X1 U670 ( .A(KEYINPUT73), .B(n597), .Z(n598) );
  NAND2_X1 U671 ( .A1(n959), .A2(n598), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n965), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n959), .A2(G868), .ZN(n600) );
  NOR2_X1 U675 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U677 ( .A(KEYINPUT74), .B(n603), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G111), .A2(n843), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT76), .ZN(n608) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n606) );
  NAND2_X1 U681 ( .A1(G123), .A2(n844), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n606), .B(n605), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U684 ( .A1(G99), .A2(n847), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G135), .A2(n848), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n908) );
  XNOR2_X1 U688 ( .A(n908), .B(G2096), .ZN(n614) );
  INV_X1 U689 ( .A(G2100), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U691 ( .A1(n959), .A2(G559), .ZN(n615) );
  XOR2_X1 U692 ( .A(n965), .B(n615), .Z(n654) );
  NAND2_X1 U693 ( .A1(n616), .A2(n654), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G67), .A2(n645), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G55), .A2(n640), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G93), .A2(n631), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G80), .A2(n634), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n656) );
  XOR2_X1 U701 ( .A(n623), .B(n656), .Z(G145) );
  NAND2_X1 U702 ( .A1(G88), .A2(n631), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G75), .A2(n634), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G62), .A2(n645), .ZN(n627) );
  NAND2_X1 U706 ( .A1(G50), .A2(n640), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U709 ( .A(KEYINPUT78), .B(n630), .Z(G303) );
  NAND2_X1 U710 ( .A1(G86), .A2(n631), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G61), .A2(n645), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n634), .A2(G73), .ZN(n635) );
  XOR2_X1 U714 ( .A(KEYINPUT2), .B(n635), .Z(n636) );
  NOR2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(G48), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(G305) );
  NAND2_X1 U718 ( .A1(G49), .A2(n640), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U721 ( .A(KEYINPUT77), .B(n643), .Z(n644) );
  NOR2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n646), .A2(G87), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(G288) );
  XNOR2_X1 U725 ( .A(n705), .B(n656), .ZN(n651) );
  XNOR2_X1 U726 ( .A(G303), .B(G305), .ZN(n649) );
  XNOR2_X1 U727 ( .A(n649), .B(G288), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U729 ( .A(KEYINPUT19), .B(n652), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(G290), .ZN(n869) );
  XNOR2_X1 U731 ( .A(n869), .B(n654), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n655), .A2(G868), .ZN(n658) );
  OR2_X1 U733 ( .A1(G868), .A2(n656), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(G295) );
  XOR2_X1 U735 ( .A(KEYINPUT79), .B(KEYINPUT21), .Z(n662) );
  NAND2_X1 U736 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U738 ( .A1(n660), .A2(G2090), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U740 ( .A1(G2072), .A2(n663), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U742 ( .A1(G120), .A2(G69), .ZN(n664) );
  NOR2_X1 U743 ( .A1(G237), .A2(n664), .ZN(n665) );
  XOR2_X1 U744 ( .A(KEYINPUT81), .B(n665), .Z(n666) );
  NAND2_X1 U745 ( .A1(G108), .A2(n666), .ZN(n824) );
  NAND2_X1 U746 ( .A1(n824), .A2(G567), .ZN(n672) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U749 ( .A1(G218), .A2(n668), .ZN(n669) );
  XNOR2_X1 U750 ( .A(KEYINPUT80), .B(n669), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n670), .A2(G96), .ZN(n825) );
  NAND2_X1 U752 ( .A1(n825), .A2(G2106), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n875) );
  NAND2_X1 U754 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U755 ( .A1(n875), .A2(n673), .ZN(n823) );
  NAND2_X1 U756 ( .A1(n823), .A2(G36), .ZN(G176) );
  NAND2_X1 U757 ( .A1(n843), .A2(G113), .ZN(n676) );
  NAND2_X1 U758 ( .A1(G101), .A2(n847), .ZN(n674) );
  XOR2_X1 U759 ( .A(KEYINPUT23), .B(n674), .Z(n675) );
  NAND2_X1 U760 ( .A1(n676), .A2(n675), .ZN(n680) );
  NAND2_X1 U761 ( .A1(G125), .A2(n844), .ZN(n678) );
  NAND2_X1 U762 ( .A1(G137), .A2(n848), .ZN(n677) );
  NAND2_X1 U763 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U764 ( .A1(n680), .A2(n679), .ZN(G160) );
  INV_X1 U765 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U766 ( .A(KEYINPUT96), .B(KEYINPUT40), .ZN(n819) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n772) );
  INV_X1 U768 ( .A(n772), .ZN(n681) );
  INV_X1 U769 ( .A(n728), .ZN(n712) );
  NAND2_X1 U770 ( .A1(n712), .A2(G2072), .ZN(n683) );
  INV_X1 U771 ( .A(KEYINPUT27), .ZN(n682) );
  XNOR2_X1 U772 ( .A(n683), .B(n682), .ZN(n685) );
  NAND2_X1 U773 ( .A1(G1956), .A2(n728), .ZN(n684) );
  NAND2_X1 U774 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U775 ( .A(KEYINPUT90), .B(n686), .Z(n704) );
  NOR2_X1 U776 ( .A1(n705), .A2(n704), .ZN(n688) );
  XNOR2_X1 U777 ( .A(KEYINPUT28), .B(KEYINPUT91), .ZN(n687) );
  XNOR2_X1 U778 ( .A(n688), .B(n687), .ZN(n709) );
  NAND2_X1 U779 ( .A1(n728), .A2(G1341), .ZN(n693) );
  INV_X1 U780 ( .A(G1996), .ZN(n933) );
  NOR2_X1 U781 ( .A1(n772), .A2(n933), .ZN(n689) );
  AND2_X1 U782 ( .A1(n773), .A2(n689), .ZN(n691) );
  XNOR2_X1 U783 ( .A(n691), .B(n690), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U785 ( .A1(n694), .A2(n965), .ZN(n695) );
  XOR2_X1 U786 ( .A(n695), .B(KEYINPUT64), .Z(n700) );
  OR2_X1 U787 ( .A1(n700), .A2(n871), .ZN(n699) );
  NOR2_X1 U788 ( .A1(n712), .A2(G1348), .ZN(n697) );
  NOR2_X1 U789 ( .A1(G2067), .A2(n728), .ZN(n696) );
  NOR2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n871), .A2(n700), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U794 ( .A(n703), .B(KEYINPUT92), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U797 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U798 ( .A(n711), .B(n710), .ZN(n717) );
  OR2_X1 U799 ( .A1(n712), .A2(G1961), .ZN(n714) );
  XNOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .ZN(n936) );
  NAND2_X1 U801 ( .A1(n712), .A2(n936), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n721) );
  AND2_X1 U803 ( .A1(n721), .A2(G171), .ZN(n715) );
  XNOR2_X1 U804 ( .A(n715), .B(KEYINPUT89), .ZN(n716) );
  NAND2_X1 U805 ( .A1(n717), .A2(n716), .ZN(n726) );
  NAND2_X1 U806 ( .A1(G8), .A2(n728), .ZN(n767) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n767), .ZN(n741) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n728), .ZN(n738) );
  NOR2_X1 U809 ( .A1(n741), .A2(n738), .ZN(n718) );
  NAND2_X1 U810 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U811 ( .A(KEYINPUT30), .B(n719), .ZN(n720) );
  NOR2_X1 U812 ( .A1(G168), .A2(n720), .ZN(n723) );
  NOR2_X1 U813 ( .A1(G171), .A2(n721), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U815 ( .A(KEYINPUT31), .B(n724), .Z(n725) );
  NAND2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n742) );
  AND2_X1 U817 ( .A1(G286), .A2(G8), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n742), .A2(n727), .ZN(n736) );
  INV_X1 U819 ( .A(G8), .ZN(n734) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n728), .ZN(n729) );
  XNOR2_X1 U821 ( .A(KEYINPUT93), .B(n729), .ZN(n732) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n767), .ZN(n730) );
  NOR2_X1 U823 ( .A1(G166), .A2(n730), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n733) );
  OR2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  AND2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U827 ( .A(n737), .B(KEYINPUT32), .ZN(n745) );
  NAND2_X1 U828 ( .A1(G8), .A2(n738), .ZN(n739) );
  XOR2_X1 U829 ( .A(KEYINPUT88), .B(n739), .Z(n740) );
  NOR2_X1 U830 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n761) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n977) );
  NOR2_X1 U834 ( .A1(G303), .A2(G1971), .ZN(n746) );
  NOR2_X1 U835 ( .A1(n977), .A2(n746), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n761), .A2(n747), .ZN(n748) );
  XNOR2_X1 U837 ( .A(n748), .B(KEYINPUT94), .ZN(n751) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n978) );
  INV_X1 U839 ( .A(n978), .ZN(n749) );
  NOR2_X1 U840 ( .A1(n767), .A2(n749), .ZN(n750) );
  NAND2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n753) );
  INV_X1 U842 ( .A(KEYINPUT33), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n758) );
  NAND2_X1 U844 ( .A1(n977), .A2(KEYINPUT33), .ZN(n754) );
  NOR2_X1 U845 ( .A1(n754), .A2(n767), .ZN(n756) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n961) );
  INV_X1 U847 ( .A(n961), .ZN(n755) );
  NOR2_X1 U848 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n771) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U851 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n767), .A2(n762), .ZN(n763) );
  XNOR2_X1 U854 ( .A(n763), .B(KEYINPUT95), .ZN(n769) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XNOR2_X1 U856 ( .A(n764), .B(KEYINPUT24), .ZN(n765) );
  XNOR2_X1 U857 ( .A(n765), .B(KEYINPUT87), .ZN(n766) );
  NOR2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n785) );
  NOR2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n814) );
  XNOR2_X1 U862 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NAND2_X1 U863 ( .A1(n848), .A2(G140), .ZN(n774) );
  XOR2_X1 U864 ( .A(KEYINPUT83), .B(n774), .Z(n776) );
  NAND2_X1 U865 ( .A1(n847), .A2(G104), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n778) );
  XNOR2_X1 U867 ( .A(KEYINPUT34), .B(KEYINPUT84), .ZN(n777) );
  XNOR2_X1 U868 ( .A(n778), .B(n777), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G116), .A2(n843), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G128), .A2(n844), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U872 ( .A(KEYINPUT35), .B(n781), .Z(n782) );
  NOR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U874 ( .A(KEYINPUT36), .B(n784), .ZN(n866) );
  NOR2_X1 U875 ( .A1(n812), .A2(n866), .ZN(n913) );
  NAND2_X1 U876 ( .A1(n814), .A2(n913), .ZN(n810) );
  NAND2_X1 U877 ( .A1(n785), .A2(n810), .ZN(n804) );
  XNOR2_X1 U878 ( .A(G1986), .B(G290), .ZN(n973) );
  AND2_X1 U879 ( .A1(n973), .A2(n814), .ZN(n802) );
  NAND2_X1 U880 ( .A1(G95), .A2(n847), .ZN(n787) );
  NAND2_X1 U881 ( .A1(G131), .A2(n848), .ZN(n786) );
  NAND2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U883 ( .A1(G107), .A2(n843), .ZN(n789) );
  NAND2_X1 U884 ( .A1(G119), .A2(n844), .ZN(n788) );
  NAND2_X1 U885 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n855) );
  XNOR2_X1 U887 ( .A(KEYINPUT85), .B(G1991), .ZN(n942) );
  NOR2_X1 U888 ( .A1(n855), .A2(n942), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G117), .A2(n843), .ZN(n793) );
  NAND2_X1 U890 ( .A1(G129), .A2(n844), .ZN(n792) );
  NAND2_X1 U891 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n847), .A2(G105), .ZN(n794) );
  XOR2_X1 U893 ( .A(KEYINPUT38), .B(n794), .Z(n795) );
  NOR2_X1 U894 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U895 ( .A1(n848), .A2(G141), .ZN(n797) );
  NAND2_X1 U896 ( .A1(n798), .A2(n797), .ZN(n858) );
  AND2_X1 U897 ( .A1(G1996), .A2(n858), .ZN(n799) );
  NOR2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n910) );
  XOR2_X1 U899 ( .A(n814), .B(KEYINPUT86), .Z(n801) );
  NOR2_X1 U900 ( .A1(n910), .A2(n801), .ZN(n807) );
  OR2_X1 U901 ( .A1(n802), .A2(n807), .ZN(n803) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n858), .ZN(n921) );
  AND2_X1 U903 ( .A1(n942), .A2(n855), .ZN(n909) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U905 ( .A1(n909), .A2(n805), .ZN(n806) );
  NOR2_X1 U906 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U907 ( .A1(n921), .A2(n808), .ZN(n809) );
  XNOR2_X1 U908 ( .A(KEYINPUT39), .B(n809), .ZN(n811) );
  NAND2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n812), .A2(n866), .ZN(n917) );
  NAND2_X1 U911 ( .A1(n813), .A2(n917), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U914 ( .A(n819), .B(n818), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n820), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U917 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(G188) );
  XOR2_X1 U920 ( .A(G120), .B(KEYINPUT98), .Z(G236) );
  XNOR2_X1 U921 ( .A(G96), .B(KEYINPUT99), .ZN(G221) );
  XOR2_X1 U922 ( .A(G69), .B(KEYINPUT100), .Z(G235) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  NOR2_X1 U925 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  NAND2_X1 U927 ( .A1(G124), .A2(n844), .ZN(n826) );
  XNOR2_X1 U928 ( .A(n826), .B(KEYINPUT44), .ZN(n828) );
  NAND2_X1 U929 ( .A1(n843), .A2(G112), .ZN(n827) );
  NAND2_X1 U930 ( .A1(n828), .A2(n827), .ZN(n832) );
  NAND2_X1 U931 ( .A1(G100), .A2(n847), .ZN(n830) );
  NAND2_X1 U932 ( .A1(G136), .A2(n848), .ZN(n829) );
  NAND2_X1 U933 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U934 ( .A1(n832), .A2(n831), .ZN(G162) );
  NAND2_X1 U935 ( .A1(G139), .A2(n848), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n847), .A2(G103), .ZN(n833) );
  XNOR2_X1 U937 ( .A(KEYINPUT105), .B(n833), .ZN(n839) );
  NAND2_X1 U938 ( .A1(G115), .A2(n843), .ZN(n835) );
  NAND2_X1 U939 ( .A1(G127), .A2(n844), .ZN(n834) );
  NAND2_X1 U940 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U941 ( .A(KEYINPUT47), .B(n836), .Z(n837) );
  XNOR2_X1 U942 ( .A(KEYINPUT106), .B(n837), .ZN(n838) );
  NOR2_X1 U943 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U944 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n842), .B(KEYINPUT107), .ZN(n903) );
  NAND2_X1 U946 ( .A1(G118), .A2(n843), .ZN(n846) );
  NAND2_X1 U947 ( .A1(G130), .A2(n844), .ZN(n845) );
  NAND2_X1 U948 ( .A1(n846), .A2(n845), .ZN(n853) );
  NAND2_X1 U949 ( .A1(G106), .A2(n847), .ZN(n850) );
  NAND2_X1 U950 ( .A1(G142), .A2(n848), .ZN(n849) );
  NAND2_X1 U951 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(KEYINPUT45), .B(n851), .Z(n852) );
  NOR2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n903), .B(n854), .ZN(n865) );
  XOR2_X1 U955 ( .A(KEYINPUT104), .B(KEYINPUT46), .Z(n857) );
  XNOR2_X1 U956 ( .A(n855), .B(KEYINPUT48), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n862) );
  XOR2_X1 U958 ( .A(n908), .B(G162), .Z(n860) );
  XOR2_X1 U959 ( .A(G160), .B(n858), .Z(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(n862), .B(n861), .Z(n863) );
  XNOR2_X1 U962 ( .A(G164), .B(n863), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n867) );
  XOR2_X1 U964 ( .A(n867), .B(n866), .Z(n868) );
  NOR2_X1 U965 ( .A1(G37), .A2(n868), .ZN(G395) );
  XNOR2_X1 U966 ( .A(G171), .B(n965), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n870), .B(n869), .ZN(n873) );
  XOR2_X1 U968 ( .A(G286), .B(n871), .Z(n872) );
  XNOR2_X1 U969 ( .A(n873), .B(n872), .ZN(n874) );
  NOR2_X1 U970 ( .A1(G37), .A2(n874), .ZN(G397) );
  INV_X1 U971 ( .A(n875), .ZN(G319) );
  XOR2_X1 U972 ( .A(KEYINPUT42), .B(G2090), .Z(n877) );
  XNOR2_X1 U973 ( .A(G2072), .B(G2078), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(n878), .B(G2100), .Z(n880) );
  XNOR2_X1 U976 ( .A(G2067), .B(G2084), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n884) );
  XOR2_X1 U978 ( .A(G2096), .B(KEYINPUT43), .Z(n882) );
  XNOR2_X1 U979 ( .A(KEYINPUT101), .B(G2678), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U981 ( .A(n884), .B(n883), .Z(G227) );
  XOR2_X1 U982 ( .A(KEYINPUT41), .B(G1961), .Z(n886) );
  XNOR2_X1 U983 ( .A(G1981), .B(G1966), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U985 ( .A(n887), .B(KEYINPUT102), .Z(n889) );
  XNOR2_X1 U986 ( .A(G1996), .B(G1991), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n893) );
  XOR2_X1 U988 ( .A(G1971), .B(G1956), .Z(n891) );
  XNOR2_X1 U989 ( .A(G1986), .B(G1976), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U991 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U992 ( .A(KEYINPUT103), .B(G2474), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(G229) );
  NOR2_X1 U994 ( .A1(G395), .A2(G397), .ZN(n896) );
  XOR2_X1 U995 ( .A(KEYINPUT109), .B(n896), .Z(n902) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n897) );
  XOR2_X1 U997 ( .A(KEYINPUT49), .B(n897), .Z(n898) );
  NAND2_X1 U998 ( .A1(G319), .A2(n898), .ZN(n899) );
  NOR2_X1 U999 ( .A1(G401), .A2(n899), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(KEYINPUT108), .B(n900), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1003 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(G2072), .B(n903), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(G164), .B(G2078), .ZN(n904) );
  NAND2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n928) );
  NOR2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(G160), .B(G2084), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1013 ( .A(KEYINPUT110), .B(n916), .Z(n918) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n925) );
  XOR2_X1 U1015 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n923) );
  XNOR2_X1 U1016 ( .A(G2090), .B(G162), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(KEYINPUT111), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1019 ( .A(n923), .B(n922), .Z(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(n926), .B(KEYINPUT113), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1023 ( .A(KEYINPUT52), .B(n929), .Z(n930) );
  NOR2_X1 U1024 ( .A1(KEYINPUT55), .A2(n930), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(KEYINPUT115), .B(n931), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n932), .A2(G29), .ZN(n1017) );
  XOR2_X1 U1027 ( .A(G2067), .B(G26), .Z(n935) );
  XNOR2_X1 U1028 ( .A(n933), .B(G32), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n940) );
  XOR2_X1 U1030 ( .A(G2072), .B(G33), .Z(n938) );
  XNOR2_X1 U1031 ( .A(n936), .B(G27), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT118), .B(n941), .ZN(n947) );
  XNOR2_X1 U1035 ( .A(KEYINPUT116), .B(G25), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(n943), .B(n942), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(G28), .A2(n944), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT117), .B(n945), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(n948), .B(KEYINPUT53), .ZN(n951) );
  XOR2_X1 U1041 ( .A(G2084), .B(G34), .Z(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(n949), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(G35), .B(G2090), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(KEYINPUT55), .B(n954), .ZN(n956) );
  INV_X1 U1047 ( .A(G29), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1049 ( .A1(n957), .A2(G11), .ZN(n1015) );
  INV_X1 U1050 ( .A(G16), .ZN(n1011) );
  XNOR2_X1 U1051 ( .A(KEYINPUT56), .B(KEYINPUT119), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(n1011), .B(n958), .ZN(n986) );
  XNOR2_X1 U1053 ( .A(G1348), .B(n959), .ZN(n984) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n960), .B(KEYINPUT120), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n963), .B(KEYINPUT57), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(G171), .B(G1961), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT121), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1341), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n982) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G303), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(n970), .B(KEYINPUT123), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(G1956), .B(KEYINPUT122), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(n971), .B(G299), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(KEYINPUT124), .B(n980), .ZN(n981) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n1013) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(G1961), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(n987), .B(G5), .ZN(n1006) );
  XOR2_X1 U1077 ( .A(G1348), .B(KEYINPUT59), .Z(n988) );
  XNOR2_X1 U1078 ( .A(G4), .B(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G20), .B(G1956), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(G1981), .B(G6), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(KEYINPUT60), .ZN(n1004) );
  XNOR2_X1 U1086 ( .A(G1976), .B(G23), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1089 ( .A(KEYINPUT126), .B(n998), .Z(n1000) );
  XNOR2_X1 U1090 ( .A(G1986), .B(G24), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT127), .B(n1001), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT58), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G21), .B(G1966), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT61), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1018), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

