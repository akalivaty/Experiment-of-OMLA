//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(G137), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT69), .Z(G160));
  AND2_X1   g050(.A1(new_n462), .A2(KEYINPUT70), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(KEYINPUT70), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n468), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n480), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n468), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT72), .A4(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n462), .A2(G126), .A3(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n462), .B2(new_n499), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n496), .B(new_n497), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(G126), .A2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n502), .ZN(new_n510));
  INV_X1    g085(.A(new_n501), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n499), .B1(new_n502), .B2(new_n501), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT4), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n514), .B2(new_n503), .ZN(new_n515));
  AOI21_X1  g090(.A(KEYINPUT73), .B1(new_n515), .B2(new_n496), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n508), .A2(new_n516), .ZN(G164));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g096(.A(KEYINPUT5), .B(G543), .Z(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(G88), .B1(new_n528), .B2(G50), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n521), .A2(new_n529), .ZN(G166));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n523), .A2(new_n524), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n518), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT74), .B(G89), .Z(new_n535));
  OAI22_X1  g110(.A1(new_n531), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n536), .A2(new_n540), .ZN(G168));
  AOI22_X1  g116(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n520), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n526), .A2(G90), .B1(new_n528), .B2(G52), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT75), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n550), .A2(new_n533), .B1(new_n534), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n520), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n528), .A2(G53), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n522), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(new_n526), .B2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  XNOR2_X1  g144(.A(G166), .B(KEYINPUT76), .ZN(G303));
  NAND2_X1  g145(.A1(new_n526), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n528), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(new_n526), .A2(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n528), .A2(G48), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(new_n520), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(G305));
  INV_X1    g155(.A(G47), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n581), .A2(new_n533), .B1(new_n534), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n520), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n534), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n590), .A2(new_n591), .B1(G54), .B2(new_n528), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n520), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n594), .B2(new_n593), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(G868), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g174(.A(new_n598), .B1(G171), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n562), .A2(new_n566), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(new_n597), .ZN(new_n605));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(KEYINPUT78), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(KEYINPUT78), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n610), .B(new_n611), .C1(G868), .C2(new_n555), .ZN(G323));
  XNOR2_X1  g187(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n613));
  XNOR2_X1  g188(.A(G323), .B(new_n613), .ZN(G282));
  NAND2_X1  g189(.A1(new_n479), .A2(G135), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT80), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n482), .A2(G123), .ZN(new_n617));
  NOR3_X1   g192(.A1(new_n468), .A2(KEYINPUT81), .A3(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n468), .B2(G111), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(G2104), .A3(new_n620), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n621), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n462), .A2(new_n471), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(G156));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n633), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT83), .B(G2100), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n646), .A2(new_n647), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n652), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n664), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n666), .B(new_n668), .C1(new_n661), .C2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G229));
  NOR2_X1   g251(.A1(G29), .A2(G35), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G162), .B2(G29), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT29), .Z(new_n679));
  INV_X1    g254(.A(G2090), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT98), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT23), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n602), .B2(new_n684), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(G1956), .ZN(new_n688));
  NOR2_X1   g263(.A1(G16), .A2(G19), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n555), .B2(G16), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(G1341), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(G1956), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT31), .B(G11), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT30), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n695), .A2(G28), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n695), .B2(G28), .ZN(new_n698));
  OAI221_X1 g273(.A(new_n694), .B1(new_n696), .B2(new_n698), .C1(new_n622), .C2(new_n697), .ZN(new_n699));
  INV_X1    g274(.A(G2084), .ZN(new_n700));
  INV_X1    g275(.A(G34), .ZN(new_n701));
  AOI21_X1  g276(.A(G29), .B1(new_n701), .B2(KEYINPUT24), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(KEYINPUT24), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G160), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n697), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n693), .B(new_n699), .C1(new_n700), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n697), .A2(G32), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n479), .A2(G141), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n482), .A2(G129), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT26), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n712), .A2(new_n713), .B1(G105), .B2(new_n471), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n708), .A2(new_n709), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n707), .B1(new_n716), .B2(new_n697), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT27), .B(G1996), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT94), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n717), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(G164), .A2(G29), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G27), .B2(G29), .ZN(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n706), .A2(new_n720), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n684), .A2(G4), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n605), .B2(new_n684), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1348), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n697), .A2(G26), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n479), .A2(G140), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n482), .A2(G128), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n468), .A2(G116), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n730), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2067), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n723), .B2(new_n722), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n725), .A2(new_n728), .A3(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n679), .A2(new_n680), .ZN(new_n740));
  NAND2_X1  g315(.A1(G168), .A2(G16), .ZN(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(KEYINPUT95), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(KEYINPUT95), .B2(new_n741), .ZN(new_n744));
  INV_X1    g319(.A(G1966), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT25), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n479), .B2(G139), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n462), .A2(G127), .ZN(new_n750));
  INV_X1    g325(.A(G115), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n470), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n468), .B1(new_n752), .B2(KEYINPUT92), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT92), .B2(new_n752), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  MUX2_X1   g330(.A(G33), .B(new_n755), .S(G29), .Z(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G2072), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(G2072), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n746), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G5), .A2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT96), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G171), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT97), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G1961), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n705), .A2(new_n700), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT93), .Z(new_n767));
  AOI211_X1 g342(.A(new_n765), .B(new_n767), .C1(G1961), .C2(new_n763), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n683), .A2(new_n739), .A3(new_n740), .A4(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n697), .A2(G25), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n771));
  INV_X1    g346(.A(G119), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n481), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n771), .B1(new_n481), .B2(new_n772), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(new_n468), .B2(G107), .ZN(new_n777));
  OR3_X1    g352(.A1(KEYINPUT86), .A2(G95), .A3(G2105), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT86), .B1(G95), .B2(G2105), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n479), .B2(G131), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n770), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT35), .B(G1991), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n784), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n697), .B1(new_n776), .B2(new_n781), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n770), .ZN(new_n788));
  OR3_X1    g363(.A1(new_n583), .A2(KEYINPUT87), .A3(new_n585), .ZN(new_n789));
  OAI21_X1  g364(.A(KEYINPUT87), .B1(new_n583), .B2(new_n585), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n684), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G24), .ZN(new_n792));
  OAI21_X1  g367(.A(G1986), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n791), .A2(G1986), .A3(new_n792), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n785), .B(new_n788), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G6), .A2(G16), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n575), .A2(new_n576), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n578), .A2(new_n520), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n797), .B1(new_n800), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT32), .B(G1981), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n684), .A2(G23), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G288), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n801), .A2(new_n802), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n803), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n684), .A2(G22), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G166), .B2(new_n684), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1971), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n810), .A2(new_n813), .A3(KEYINPUT34), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT88), .B1(new_n796), .B2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n795), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n816), .A2(new_n793), .B1(new_n783), .B2(new_n784), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT88), .ZN(new_n818));
  INV_X1    g393(.A(G1971), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n812), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n802), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n801), .B(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n807), .A2(new_n809), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT34), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n820), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n817), .A2(new_n818), .A3(new_n825), .A4(new_n788), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT34), .B1(new_n810), .B2(new_n813), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT90), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n829), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n828), .B1(new_n832), .B2(KEYINPUT89), .ZN(new_n833));
  INV_X1    g408(.A(new_n829), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n815), .B2(new_n826), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT89), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n831), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT36), .B1(new_n835), .B2(new_n836), .ZN(new_n839));
  AOI211_X1 g414(.A(KEYINPUT89), .B(new_n834), .C1(new_n815), .C2(new_n826), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n839), .A2(KEYINPUT90), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT91), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT90), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n835), .B2(new_n828), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n839), .B2(new_n840), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n832), .A2(KEYINPUT89), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n846), .A2(new_n843), .A3(KEYINPUT36), .A4(new_n837), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT91), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n769), .B1(new_n842), .B2(new_n849), .ZN(G311));
  AND4_X1   g425(.A1(new_n740), .A2(new_n683), .A3(new_n739), .A4(new_n768), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n848), .B1(new_n845), .B2(new_n847), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(G150));
  NAND2_X1  g429(.A1(new_n605), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  INV_X1    g431(.A(G55), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n857), .A2(new_n533), .B1(new_n534), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n520), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n555), .A2(new_n862), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n554), .A2(new_n552), .B1(new_n859), .B2(new_n861), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n856), .B(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n868), .A2(new_n869), .A3(G860), .ZN(new_n870));
  INV_X1    g445(.A(new_n862), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G860), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT99), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  OR2_X1    g449(.A1(new_n870), .A2(new_n874), .ZN(G145));
  OR2_X1    g450(.A1(G162), .A2(new_n622), .ZN(new_n876));
  NAND2_X1  g451(.A1(G162), .A2(new_n622), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT100), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n880), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n704), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(G160), .A3(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n735), .A2(new_n506), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n735), .A2(new_n506), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n886), .A2(new_n715), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n715), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n888), .A2(new_n889), .A3(new_n755), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n755), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n782), .B(new_n626), .ZN(new_n893));
  OR2_X1    g468(.A1(G106), .A2(G2105), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n894), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n895));
  INV_X1    g470(.A(G130), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n481), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(G142), .B2(new_n479), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n893), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n892), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  INV_X1    g477(.A(new_n899), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n903), .A2(new_n890), .A3(new_n891), .A4(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n892), .B1(KEYINPUT101), .B2(new_n899), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n883), .A2(new_n905), .A3(new_n884), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n901), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g484(.A(G305), .B(new_n586), .ZN(new_n910));
  XNOR2_X1  g485(.A(G166), .B(G288), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(KEYINPUT104), .B2(KEYINPUT42), .ZN(new_n913));
  NAND2_X1  g488(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT105), .Z(new_n915));
  XOR2_X1   g490(.A(new_n913), .B(new_n915), .Z(new_n916));
  XNOR2_X1  g491(.A(new_n865), .B(KEYINPUT102), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n608), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n605), .A2(new_n602), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND2_X1  g495(.A1(G299), .A2(new_n597), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT103), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n921), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT103), .B1(new_n925), .B2(KEYINPUT41), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n918), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n925), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n918), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n916), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G868), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(G868), .B2(new_n862), .ZN(G295));
  OAI21_X1  g508(.A(new_n932), .B1(G868), .B2(new_n862), .ZN(G331));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n547), .B2(new_n548), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n937), .A2(new_n865), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n547), .A2(new_n936), .A3(new_n548), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(G286), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n865), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n938), .B2(new_n942), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n944), .A2(new_n945), .B1(new_n923), .B2(new_n922), .ZN(new_n946));
  INV_X1    g521(.A(new_n942), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n937), .A2(new_n865), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n940), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(new_n943), .A3(new_n929), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n912), .ZN(new_n952));
  AOI21_X1  g527(.A(G37), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n924), .A2(new_n927), .B1(new_n949), .B2(new_n943), .ZN(new_n955));
  INV_X1    g530(.A(new_n950), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n954), .B1(new_n957), .B2(new_n912), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n925), .A2(KEYINPUT41), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n919), .A2(new_n921), .A3(new_n920), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n962), .A2(new_n926), .B1(new_n944), .B2(new_n945), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(new_n912), .A3(new_n950), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(KEYINPUT108), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n953), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n957), .A2(new_n954), .A3(new_n912), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n964), .A2(KEYINPUT108), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT107), .B1(new_n955), .B2(new_n956), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n963), .A2(new_n973), .A3(new_n950), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n974), .A3(new_n952), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n970), .A2(new_n971), .A3(new_n902), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n935), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n970), .A2(new_n902), .A3(new_n975), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT43), .B1(new_n968), .B2(new_n969), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n978), .A2(KEYINPUT43), .B1(new_n953), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n935), .B2(new_n980), .ZN(G397));
  XNOR2_X1  g556(.A(KEYINPUT109), .B(G1384), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n515), .B2(new_n496), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n467), .A2(new_n473), .A3(G40), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n983), .A2(new_n984), .A3(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT110), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n988), .A2(new_n716), .ZN(new_n989));
  INV_X1    g564(.A(new_n985), .ZN(new_n990));
  INV_X1    g565(.A(G2067), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n735), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n715), .A2(G1996), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n782), .B(new_n784), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1986), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n586), .B(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n985), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n508), .B2(new_n516), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n468), .B1(new_n463), .B2(new_n465), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n469), .A2(new_n472), .ZN(new_n1006));
  INV_X1    g581(.A(G40), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n983), .A2(new_n1009), .A3(KEYINPUT45), .ZN(new_n1010));
  INV_X1    g585(.A(new_n982), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT111), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT56), .B(G2072), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1004), .A2(new_n1008), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1956), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n506), .A2(new_n507), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n515), .A2(KEYINPUT73), .A3(new_n496), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT50), .B(G1384), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n515), .B2(new_n496), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1008), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1017), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1016), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n1026));
  XNOR2_X1  g601(.A(G299), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n984), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n1022), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT118), .ZN(new_n1033));
  INV_X1    g608(.A(G1348), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1030), .B(new_n1035), .C1(new_n1031), .C2(new_n1022), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n506), .A2(new_n1001), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(new_n984), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n991), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT119), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n1043), .A3(new_n1040), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1016), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n605), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1029), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT61), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1016), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1027), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT122), .B(new_n1049), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1029), .A2(KEYINPUT61), .A3(new_n1046), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1029), .A2(KEYINPUT123), .A3(new_n1046), .A4(KEYINPUT61), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1039), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1008), .B1(new_n1031), .B2(KEYINPUT45), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1009), .B1(new_n983), .B2(KEYINPUT45), .ZN(new_n1067));
  AND4_X1   g642(.A1(new_n1009), .A2(new_n506), .A3(KEYINPUT45), .A4(new_n1011), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1070), .B2(new_n986), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n555), .A2(KEYINPUT120), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT121), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1004), .A2(new_n986), .A3(new_n1008), .A4(new_n1014), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1064), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1072), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1074), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1077), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1081));
  AOI211_X1 g656(.A(KEYINPUT121), .B(new_n1072), .C1(new_n1075), .C2(new_n1064), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT59), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1056), .A2(new_n1061), .A3(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1037), .A2(new_n1043), .A3(new_n1040), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1043), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1087));
  OR3_X1    g662(.A1(new_n1086), .A2(new_n1087), .A3(KEYINPUT60), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n597), .B1(new_n1045), .B2(KEYINPUT60), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT60), .B(new_n597), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1048), .B1(new_n1085), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1961), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1033), .A2(new_n1094), .A3(new_n1036), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1004), .A2(KEYINPUT112), .A3(new_n1008), .A4(new_n1014), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n723), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1096), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n473), .B(KEYINPUT124), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(G2078), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(G40), .A3(new_n467), .A4(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n983), .A2(KEYINPUT45), .ZN(new_n1107));
  OR3_X1    g682(.A1(new_n1069), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1103), .A2(KEYINPUT125), .A3(G301), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1008), .B1(new_n1021), .B2(KEYINPUT45), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(KEYINPUT45), .B2(new_n1031), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1105), .ZN(new_n1113));
  AOI21_X1  g688(.A(G2078), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1095), .B(new_n1113), .C1(new_n1114), .C2(KEYINPUT53), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G171), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1095), .B(new_n1108), .C1(new_n1114), .C2(KEYINPUT53), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n1119), .B2(G171), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1109), .B(new_n1110), .C1(new_n1117), .C2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1110), .B1(new_n1119), .B2(G171), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(G171), .B2(new_n1115), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1030), .B(new_n700), .C1(new_n1031), .C2(new_n1022), .ZN(new_n1124));
  OAI211_X1 g699(.A(G168), .B(new_n1124), .C1(new_n1112), .C2(G1966), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G8), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1003), .B(G1384), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n745), .B1(new_n1127), .B2(new_n1111), .ZN(new_n1128));
  AOI21_X1  g703(.A(G168), .B1(new_n1128), .B2(new_n1124), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT51), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1125), .A2(new_n1131), .A3(G8), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1098), .A2(new_n819), .A3(new_n1099), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1032), .A2(G2090), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(G303), .A2(G8), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT55), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1139), .A3(G8), .ZN(new_n1140));
  INV_X1    g715(.A(G1981), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n579), .A2(new_n1141), .A3(new_n575), .A4(new_n576), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT113), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n577), .A2(KEYINPUT113), .A3(new_n1141), .A4(new_n579), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1144), .A2(new_n1145), .B1(G1981), .B2(G305), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT49), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(G8), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1039), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n1146), .B2(KEYINPUT49), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(G1976), .ZN(new_n1153));
  OR2_X1    g728(.A1(G288), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT52), .B1(G288), .B2(new_n1153), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1150), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT52), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1152), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1140), .A2(new_n1160), .ZN(new_n1161));
  OR3_X1    g736(.A1(new_n1020), .A2(G2090), .A3(new_n1023), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1134), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT117), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT117), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1134), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1164), .A2(G8), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1139), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1161), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1121), .A2(new_n1123), .A3(new_n1133), .A4(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1093), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT114), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1158), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n1157), .B2(new_n1155), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1175), .B(KEYINPUT114), .C1(new_n1148), .C2(new_n1151), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1149), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n1178), .A3(new_n1139), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1150), .B(KEYINPUT115), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1152), .A2(G1976), .A3(G288), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT116), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1180), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1130), .A2(new_n1186), .A3(new_n1132), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1186), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1187), .A2(new_n1188), .A3(new_n1116), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1185), .B1(new_n1189), .B2(new_n1169), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1149), .B(G286), .C1(new_n1128), .C2(new_n1124), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n1169), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1191), .A2(KEYINPUT63), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1177), .A2(new_n1140), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1178), .A2(new_n1139), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1190), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1000), .B1(new_n1171), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT46), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n988), .B(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n992), .A2(new_n716), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n985), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT47), .ZN(new_n1204));
  NOR4_X1   g779(.A1(new_n989), .A2(new_n994), .A3(new_n786), .A4(new_n782), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n735), .A2(G2067), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n985), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n985), .A2(new_n998), .A3(new_n586), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT48), .Z(new_n1209));
  OR2_X1    g784(.A1(new_n997), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1204), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1211), .B(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1198), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g789(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n908), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1217), .A2(new_n980), .ZN(G308));
  OR2_X1    g792(.A1(new_n1217), .A2(new_n980), .ZN(G225));
endmodule


