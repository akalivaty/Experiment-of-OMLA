//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n601, new_n603, new_n604, new_n605,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1119, new_n1120;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g039(.A(G2105), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n461), .A2(G137), .ZN(new_n467));
  AND2_X1   g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  MUX2_X1   g051(.A(G100), .B(G112), .S(G2105), .Z(new_n477));
  AOI22_X1  g052(.A1(new_n476), .A2(G124), .B1(G2104), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n466), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n466), .C1(new_n472), .C2(new_n473), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n461), .A2(new_n487), .A3(G138), .A4(new_n466), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  INV_X1    g066(.A(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n466), .A2(G102), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2105), .ZN(new_n494));
  AOI211_X1 g069(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G102), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT69), .B1(new_n497), .B2(G2104), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n490), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n484), .B1(new_n489), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n474), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(new_n491), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n497), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n486), .A2(new_n488), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(KEYINPUT70), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n512), .B1(new_n511), .B2(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g093(.A(KEYINPUT5), .B(G543), .Z(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(G88), .B1(new_n525), .B2(G50), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n518), .A2(new_n526), .ZN(G166));
  XNOR2_X1  g102(.A(new_n525), .B(KEYINPUT73), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(new_n522), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT74), .B(G89), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(new_n533), .B1(G63), .B2(G651), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n531), .B1(new_n534), .B2(new_n519), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n529), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AND2_X1   g112(.A1(new_n528), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n523), .A2(G90), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n538), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n519), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G651), .B1(new_n523), .B2(G81), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n525), .B(KEYINPUT73), .Z(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  XOR2_X1   g130(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n556));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT76), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n519), .B2(new_n562), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(KEYINPUT77), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(KEYINPUT77), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(G651), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n525), .A2(G53), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT9), .Z(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n523), .A2(G91), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(G299));
  INV_X1    g146(.A(G166), .ZN(G303));
  NAND2_X1  g147(.A1(new_n523), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n525), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n525), .A2(G48), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  INV_X1    g154(.A(new_n523), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n578), .B1(new_n579), .B2(new_n540), .C1(new_n580), .C2(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n523), .A2(G85), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  XOR2_X1   g159(.A(KEYINPUT78), .B(G47), .Z(new_n585));
  OAI221_X1 g160(.A(new_n583), .B1(new_n540), .B2(new_n584), .C1(new_n549), .C2(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n590));
  OR3_X1    g165(.A1(new_n580), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n580), .B2(new_n589), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n540), .C2(new_n593), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n528), .A2(G54), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n588), .B1(new_n587), .B2(new_n596), .ZN(G284));
  AOI21_X1  g172(.A(new_n588), .B1(new_n587), .B2(new_n596), .ZN(G321));
  MUX2_X1   g173(.A(G286), .B(G299), .S(new_n587), .Z(G297));
  MUX2_X1   g174(.A(G286), .B(G299), .S(new_n587), .Z(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n596), .B1(new_n601), .B2(G860), .ZN(G148));
  NOR2_X1   g177(.A1(new_n551), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(new_n596), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G559), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n603), .B1(new_n605), .B2(G868), .ZN(G323));
  XOR2_X1   g181(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n607));
  XNOR2_X1  g182(.A(G323), .B(new_n607), .ZN(G282));
  NAND2_X1  g183(.A1(new_n480), .A2(G135), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n476), .A2(G123), .ZN(new_n610));
  MUX2_X1   g185(.A(G99), .B(G111), .S(G2105), .Z(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G2104), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G2096), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n613), .A2(G2096), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT12), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n619), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n616), .A2(new_n617), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2438), .Z(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2430), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(KEYINPUT14), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT82), .ZN(new_n629));
  INV_X1    g204(.A(new_n625), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n626), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2443), .B(G2446), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  OAI21_X1  g212(.A(G14), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n636), .B2(new_n637), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  INV_X1    g221(.A(new_n642), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n643), .B1(new_n649), .B2(new_n640), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n641), .B2(new_n648), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n641), .A2(new_n644), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n647), .B1(new_n652), .B2(KEYINPUT17), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n646), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(new_n615), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT84), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n659), .A2(new_n660), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n658), .A2(new_n661), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n658), .B2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1981), .B(G1986), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1991), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT85), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NOR2_X1   g254(.A1(G171), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G5), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(G1961), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(G1961), .ZN(new_n684));
  NOR2_X1   g259(.A1(G168), .A2(new_n679), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n679), .B2(G21), .ZN(new_n686));
  INV_X1    g261(.A(G1966), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n683), .A2(new_n684), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(G4), .A2(G16), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT90), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n604), .B2(new_n679), .ZN(new_n693));
  INV_X1    g268(.A(G1348), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G19), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n552), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G1341), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n614), .A2(G29), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT31), .B(G11), .Z(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT30), .B(G28), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(KEYINPUT24), .A2(G34), .ZN(new_n704));
  NOR2_X1   g279(.A1(KEYINPUT24), .A2(G34), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n470), .B2(new_n701), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2084), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n698), .A2(new_n699), .A3(new_n703), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n701), .A2(G26), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G104), .B(G116), .S(G2105), .Z(new_n713));
  AOI22_X1  g288(.A1(new_n476), .A2(G128), .B1(G2104), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G140), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n479), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n712), .B1(new_n716), .B2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G2067), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OR4_X1    g294(.A1(new_n690), .A2(new_n695), .A3(new_n709), .A4(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G29), .A2(G32), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n480), .A2(G141), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n476), .A2(G129), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n722), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT95), .Z(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n679), .A2(G20), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT23), .Z(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G299), .B2(G16), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1956), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n734), .A2(new_n735), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G29), .A2(G35), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G162), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT29), .ZN(new_n743));
  INV_X1    g318(.A(G2090), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n746));
  NAND3_X1  g321(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  INV_X1    g324(.A(G139), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n748), .B1(new_n466), .B2(new_n749), .C1(new_n479), .C2(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G33), .B(new_n751), .S(G29), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT93), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2072), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n701), .A2(G27), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G164), .B2(new_n701), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n745), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n720), .A2(new_n740), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G6), .A2(G16), .ZN(new_n761));
  INV_X1    g336(.A(G305), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G16), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT32), .B(G1981), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n679), .A2(G22), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(KEYINPUT89), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(KEYINPUT89), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(G166), .C2(new_n679), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(G1971), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(G1971), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n679), .A2(G23), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n576), .B2(new_n679), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT33), .B(G1976), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n765), .A2(new_n770), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(KEYINPUT34), .ZN(new_n777));
  NOR2_X1   g352(.A1(G25), .A2(G29), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n466), .A2(G95), .ZN(new_n779));
  NAND2_X1  g354(.A1(G107), .A2(G2105), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n492), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n480), .B2(G131), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n476), .A2(KEYINPUT87), .A3(G119), .ZN(new_n783));
  AOI21_X1  g358(.A(KEYINPUT87), .B1(new_n476), .B2(G119), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n778), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT35), .B(G1991), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT88), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n787), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n776), .A2(KEYINPUT34), .ZN(new_n791));
  MUX2_X1   g366(.A(G24), .B(G290), .S(G16), .Z(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1986), .Z(new_n793));
  NAND4_X1  g368(.A1(new_n777), .A2(new_n790), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT36), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n760), .A2(new_n795), .ZN(G150));
  INV_X1    g371(.A(G150), .ZN(G311));
  AOI22_X1  g372(.A1(new_n528), .A2(G55), .B1(G93), .B2(new_n523), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n540), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT96), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G860), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT37), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n551), .B(KEYINPUT97), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(new_n802), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT38), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n604), .A2(new_n601), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT39), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n811), .A2(KEYINPUT98), .ZN(new_n812));
  AOI21_X1  g387(.A(G860), .B1(new_n810), .B2(KEYINPUT39), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n811), .B2(KEYINPUT98), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n804), .B1(new_n812), .B2(new_n814), .ZN(G145));
  NAND2_X1  g390(.A1(new_n506), .A2(new_n507), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n716), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n729), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(KEYINPUT99), .B2(new_n751), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n785), .B(new_n621), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT101), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT101), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n822), .B(new_n823), .C1(G118), .C2(new_n466), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n476), .A2(G130), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n480), .A2(new_n826), .A3(G142), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n480), .B2(G142), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n824), .B(new_n825), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n820), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n819), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n751), .A2(KEYINPUT99), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n833), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n482), .B(G160), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n614), .ZN(new_n837));
  OR3_X1    g412(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G37), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n837), .B1(new_n834), .B2(new_n835), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g417(.A1(new_n802), .A2(G868), .ZN(new_n843));
  XNOR2_X1  g418(.A(G299), .B(new_n596), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT41), .Z(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n806), .B(new_n605), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n844), .B2(new_n847), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT42), .ZN(new_n850));
  XNOR2_X1  g425(.A(G290), .B(G288), .ZN(new_n851));
  XNOR2_X1  g426(.A(G166), .B(G305), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT102), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n850), .B(new_n854), .Z(new_n855));
  AOI21_X1  g430(.A(new_n843), .B1(new_n855), .B2(G868), .ZN(G295));
  AOI21_X1  g431(.A(new_n843), .B1(new_n855), .B2(G868), .ZN(G331));
  XOR2_X1   g432(.A(G286), .B(G301), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n806), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n844), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(KEYINPUT103), .ZN(new_n862));
  INV_X1    g437(.A(new_n853), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n845), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(KEYINPUT103), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n862), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n866), .A2(new_n839), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n853), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(KEYINPUT43), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n866), .A2(new_n839), .ZN(new_n873));
  INV_X1    g448(.A(new_n861), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n874), .A2(new_n875), .B1(new_n845), .B2(new_n859), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n861), .A2(KEYINPUT104), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n863), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n870), .A2(new_n871), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n870), .A2(KEYINPUT105), .A3(new_n879), .A4(new_n871), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n867), .A2(new_n872), .A3(new_n869), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT43), .B1(new_n873), .B2(new_n878), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(KEYINPUT44), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(G397));
  AOI21_X1  g462(.A(G1384), .B1(new_n506), .B2(new_n507), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n465), .A2(new_n469), .A3(G40), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT45), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n786), .A2(new_n789), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n716), .B(new_n718), .ZN(new_n892));
  INV_X1    g467(.A(G1996), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n729), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n786), .A2(new_n789), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n891), .A2(new_n892), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G290), .B(G1986), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n890), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n888), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(new_n889), .ZN(new_n900));
  INV_X1    g475(.A(G8), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT109), .Z(new_n903));
  INV_X1    g478(.A(KEYINPUT49), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n579), .A2(new_n540), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n906));
  OAI21_X1  g481(.A(G1981), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n762), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(G305), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n904), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n762), .A2(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(G305), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT49), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n902), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G1976), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n915), .A2(new_n916), .A3(new_n576), .ZN(new_n917));
  NOR2_X1   g492(.A1(G305), .A2(G1981), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n903), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(G166), .A2(new_n901), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT50), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n889), .B1(new_n888), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  AOI21_X1  g500(.A(G1384), .B1(new_n500), .B2(new_n508), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n922), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n489), .A2(new_n499), .A3(new_n484), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT70), .B1(new_n506), .B2(new_n507), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(KEYINPUT106), .A3(KEYINPUT50), .ZN(new_n932));
  AOI211_X1 g507(.A(G2090), .B(new_n924), .C1(new_n927), .C2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n889), .B1(new_n888), .B2(KEYINPUT45), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n926), .B2(KEYINPUT45), .ZN(new_n935));
  INV_X1    g510(.A(G1971), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(G8), .B(new_n921), .C1(new_n933), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n576), .A2(G1976), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT52), .B1(G288), .B2(new_n916), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n902), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n940), .B(G8), .C1(new_n899), .C2(new_n889), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n943), .A2(KEYINPUT107), .A3(KEYINPUT52), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT107), .B1(new_n943), .B2(KEYINPUT52), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n915), .B(new_n942), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n919), .B1(new_n939), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G2084), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT106), .B1(new_n931), .B2(KEYINPUT50), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n926), .A2(new_n925), .A3(new_n922), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n948), .B(new_n923), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n926), .A2(KEYINPUT45), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n889), .B1(new_n899), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n687), .ZN(new_n956));
  AOI211_X1 g531(.A(new_n901), .B(G286), .C1(new_n951), .C2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n921), .ZN(new_n958));
  INV_X1    g533(.A(new_n889), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT50), .B1(new_n509), .B2(new_n928), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n899), .A2(new_n922), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n744), .B(new_n959), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n962), .A2(new_n937), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n958), .B1(new_n963), .B2(new_n901), .ZN(new_n964));
  INV_X1    g539(.A(new_n946), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n957), .A2(new_n964), .A3(new_n939), .A4(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n744), .B(new_n923), .C1(new_n949), .C2(new_n950), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n901), .B1(new_n970), .B2(new_n937), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n946), .B1(new_n971), .B2(new_n921), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(KEYINPUT110), .A3(new_n964), .A4(new_n957), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT63), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n968), .A2(new_n969), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n971), .A2(new_n921), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n976), .A2(new_n972), .A3(KEYINPUT63), .A4(new_n957), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n968), .A2(new_n974), .A3(new_n973), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT111), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n947), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n982));
  NOR2_X1   g557(.A1(G299), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n566), .A2(new_n570), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n566), .A2(KEYINPUT113), .A3(new_n570), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n568), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT112), .B(KEYINPUT57), .Z(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(KEYINPUT114), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  INV_X1    g567(.A(new_n990), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n983), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n935), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT56), .B(G2072), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n960), .A2(new_n961), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n889), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1001), .B2(G1956), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n1002), .A2(KEYINPUT117), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(KEYINPUT117), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n996), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n923), .B1(new_n949), .B2(new_n950), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT115), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n924), .B1(new_n927), .B2(new_n932), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n694), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n1012));
  INV_X1    g587(.A(new_n900), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(G2067), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1012), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1002), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n604), .B1(new_n996), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1005), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1025));
  AOI211_X1 g600(.A(KEYINPUT115), .B(new_n924), .C1(new_n927), .C2(new_n932), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1025), .A2(new_n1026), .A3(G1348), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT116), .B1(new_n1027), .B2(new_n1014), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n604), .B1(new_n1030), .B2(KEYINPUT60), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1023), .B(new_n596), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1024), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT61), .B1(new_n995), .B2(new_n1002), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1005), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT118), .B(KEYINPUT61), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n996), .A2(new_n1019), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n995), .A2(new_n1002), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT58), .B(G1341), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n935), .A2(G1996), .B1(new_n900), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n552), .ZN(new_n1042));
  XOR2_X1   g617(.A(new_n1042), .B(KEYINPUT59), .Z(new_n1043));
  NOR3_X1   g618(.A1(new_n1035), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1022), .B1(new_n1033), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT121), .B(G1961), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1007), .A2(new_n1010), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n935), .B2(G2078), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT53), .B1(new_n1051), .B2(G2078), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1051), .B2(G2078), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n954), .B(new_n1053), .C1(new_n953), .C2(new_n899), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1048), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1046), .B1(new_n1056), .B2(G171), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n952), .A2(KEYINPUT53), .A3(new_n757), .A4(new_n954), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1050), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1048), .A2(G301), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1057), .A2(KEYINPUT123), .A3(new_n1060), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n901), .B1(new_n951), .B2(new_n956), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G286), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G286), .A2(G8), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(KEYINPUT119), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT51), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1066), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1067), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n972), .A2(new_n964), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1056), .A2(G171), .ZN(new_n1079));
  AOI21_X1  g654(.A(G301), .B1(new_n1048), .B2(new_n1059), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1046), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1065), .A2(new_n1077), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT124), .B(new_n981), .C1(new_n1045), .C2(new_n1082), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1077), .A2(KEYINPUT62), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1077), .A2(KEYINPUT62), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1078), .A3(new_n1080), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT60), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n596), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1089), .A2(new_n1090), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1035), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1021), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1081), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT124), .B1(new_n1098), .B2(new_n981), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n898), .B1(new_n1087), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(G290), .A2(G1986), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n890), .ZN(new_n1102));
  XOR2_X1   g677(.A(new_n1102), .B(KEYINPUT48), .Z(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(new_n896), .B2(new_n890), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n892), .A2(new_n730), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n890), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT126), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n890), .B(new_n893), .C1(KEYINPUT125), .C2(KEYINPUT46), .ZN(new_n1108));
  NAND2_X1  g683(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n892), .A2(new_n894), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1114), .A2(new_n895), .B1(G2067), .B2(new_n716), .ZN(new_n1115));
  AOI211_X1 g690(.A(new_n1104), .B(new_n1113), .C1(new_n890), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1100), .A2(new_n1116), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g692(.A1(new_n870), .A2(new_n879), .ZN(new_n1119));
  NOR4_X1   g693(.A1(G229), .A2(G401), .A3(new_n459), .A4(G227), .ZN(new_n1120));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n841), .A3(new_n1120), .ZN(G225));
  INV_X1    g695(.A(G225), .ZN(G308));
endmodule


