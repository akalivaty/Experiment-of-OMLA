//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n440, new_n441, new_n443, new_n444, new_n445,
    new_n453, new_n457, new_n458, new_n459, new_n460, new_n461, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n565, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n439));
  OR2_X1    g014(.A1(new_n439), .A2(G69), .ZN(new_n440));
  NAND2_X1  g015(.A1(new_n439), .A2(G69), .ZN(new_n441));
  NAND2_X1  g016(.A1(new_n440), .A2(new_n441), .ZN(G235));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n443));
  OR2_X1    g018(.A1(new_n443), .A2(G120), .ZN(new_n444));
  NAND2_X1  g019(.A1(new_n443), .A2(G120), .ZN(new_n445));
  NAND2_X1  g020(.A1(new_n444), .A2(new_n445), .ZN(G236));
  INV_X1    g021(.A(G57), .ZN(G237));
  INV_X1    g022(.A(G108), .ZN(G238));
  NAND4_X1  g023(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g024(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g025(.A(G452), .Z(G391));
  AND2_X1   g026(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g027(.A1(G7), .A2(G661), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g029(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g030(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g031(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT2), .Z(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR4_X1   g034(.A1(G235), .A2(G236), .A3(G237), .A4(G238), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(G325));
  INV_X1    g037(.A(G325), .ZN(G261));
  NAND2_X1  g038(.A1(new_n459), .A2(G2106), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G567), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT66), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(G101), .A2(new_n470), .B1(new_n476), .B2(G137), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n478), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(new_n475), .A2(new_n468), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n476), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n475), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(new_n468), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n472), .A2(new_n474), .A3(G126), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n472), .A2(new_n474), .A3(G138), .A4(new_n468), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT67), .B(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n495), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT68), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n495), .A2(new_n499), .A3(new_n505), .A4(new_n502), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT69), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n508), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n511), .A2(new_n517), .B1(new_n522), .B2(G88), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n518), .A2(new_n520), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n523), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n518), .A2(new_n520), .ZN(new_n531));
  INV_X1    g106(.A(G63), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n515), .A2(G51), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT70), .B(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n524), .A2(new_n508), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n534), .A2(new_n537), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  INV_X1    g117(.A(G77), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n531), .A2(new_n542), .B1(new_n543), .B2(new_n512), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT71), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n546));
  OAI221_X1 g121(.A(new_n546), .B1(new_n543), .B2(new_n512), .C1(new_n531), .C2(new_n542), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(G651), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n521), .A2(new_n549), .B1(new_n509), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  AOI22_X1  g129(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n526), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n524), .A2(G81), .A3(new_n508), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n515), .A2(G43), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n557), .A2(KEYINPUT72), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT72), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G188));
  NAND3_X1  g144(.A1(new_n515), .A2(KEYINPUT73), .A3(G53), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n515), .A2(KEYINPUT73), .A3(KEYINPUT9), .A4(G53), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n531), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n524), .A2(G91), .A3(new_n508), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n522), .A2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n515), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT74), .B1(new_n521), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n524), .A2(new_n589), .A3(G86), .A4(new_n508), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n531), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(G48), .B2(new_n515), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(G305));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n521), .A2(new_n597), .B1(new_n509), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n524), .A2(G60), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n526), .B1(new_n601), .B2(new_n602), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT75), .B1(new_n607), .B2(new_n599), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G171), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT77), .B(KEYINPUT78), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(KEYINPUT10), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n522), .A2(G92), .A3(new_n614), .A4(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n617), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n615), .A2(new_n616), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI22_X1  g196(.A1(new_n619), .A2(new_n620), .B1(new_n521), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(G79), .A2(G543), .ZN(new_n623));
  INV_X1    g198(.A(G66), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n531), .B2(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n625), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n618), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n612), .B1(G868), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT76), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(KEYINPUT76), .B2(new_n611), .ZN(G284));
  OAI21_X1  g205(.A(new_n629), .B1(KEYINPUT76), .B2(new_n611), .ZN(G321));
  NAND2_X1  g206(.A1(G286), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n581), .B2(G868), .ZN(G297));
  OAI21_X1  g208(.A(new_n632), .B1(new_n581), .B2(G868), .ZN(G280));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n627), .B1(new_n635), .B2(G860), .ZN(G148));
  NAND2_X1  g211(.A1(new_n627), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g215(.A(new_n475), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n470), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT79), .B(G2100), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n484), .A2(G123), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n476), .A2(G135), .ZN(new_n648));
  OR2_X1    g223(.A1(G99), .A2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n649), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT80), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XOR2_X1   g231(.A(G2443), .B(G2446), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1341), .B(G1348), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT15), .B(G2435), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT14), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n660), .B(new_n665), .Z(new_n666));
  INV_X1    g241(.A(G14), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n677), .A2(KEYINPUT82), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n670), .A2(new_n671), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(KEYINPUT82), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n679), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n673), .B(KEYINPUT17), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n683), .A3(new_n672), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n676), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n690), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  AOI22_X1  g271(.A1(new_n694), .A2(KEYINPUT20), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n698), .A2(new_n690), .A3(new_n693), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n697), .B(new_n699), .C1(KEYINPUT20), .C2(new_n694), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1986), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1981), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1991), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n702), .B(new_n705), .ZN(G229));
  MUX2_X1   g281(.A(G35), .B(new_n489), .S(G29), .Z(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT29), .Z(new_n708));
  INV_X1    g283(.A(G2090), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G4), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n627), .B2(new_n710), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n708), .A2(new_n709), .B1(G1348), .B2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(KEYINPUT24), .A2(G34), .ZN(new_n714));
  NOR2_X1   g289(.A1(KEYINPUT24), .A2(G34), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n714), .A2(new_n715), .A3(G29), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n482), .B2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT92), .Z(new_n718));
  OAI221_X1 g293(.A(new_n713), .B1(G2084), .B2(new_n718), .C1(new_n709), .C2(new_n708), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n712), .A2(G1348), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT28), .ZN(new_n721));
  INV_X1    g296(.A(G26), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n484), .A2(G128), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n476), .A2(G140), .ZN(new_n726));
  OR2_X1    g301(.A1(G104), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n724), .B1(new_n729), .B2(G29), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n723), .B1(new_n730), .B2(new_n721), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G2067), .ZN(new_n732));
  OAI21_X1  g307(.A(KEYINPUT96), .B1(G5), .B2(G16), .ZN(new_n733));
  OR3_X1    g308(.A1(KEYINPUT96), .A2(G5), .A3(G16), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n733), .B(new_n734), .C1(G301), .C2(new_n710), .ZN(new_n735));
  INV_X1    g310(.A(G1961), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n731), .A2(G2067), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n732), .A2(new_n737), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n719), .A2(new_n720), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n651), .ZN(new_n742));
  INV_X1    g317(.A(G28), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n743), .B2(KEYINPUT30), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n742), .A2(G29), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G21), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G168), .B2(G16), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n484), .A2(G129), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT93), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  AOI22_X1  g327(.A1(G105), .A2(new_n470), .B1(new_n476), .B2(G141), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G29), .B2(G32), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n746), .B1(G1966), .B2(new_n748), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n710), .A2(G20), .ZN(new_n759));
  OAI211_X1 g334(.A(KEYINPUT23), .B(new_n759), .C1(new_n581), .C2(new_n710), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(KEYINPUT23), .B2(new_n759), .ZN(new_n761));
  INV_X1    g336(.A(G1956), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT31), .B(G11), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n748), .A2(G1966), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT95), .Z(new_n766));
  NOR4_X1   g341(.A1(new_n758), .A2(new_n763), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G27), .A2(G29), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G164), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT97), .B(G2078), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n741), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n476), .A2(G139), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT25), .Z(new_n775));
  AOI22_X1  g350(.A1(new_n641), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n775), .C1(new_n776), .C2(new_n468), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT90), .ZN(new_n778));
  MUX2_X1   g353(.A(G33), .B(new_n778), .S(G29), .Z(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT91), .B(G2072), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n756), .A2(new_n757), .B1(new_n718), .B2(G2084), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n772), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n710), .A2(G19), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n563), .B2(new_n710), .ZN(new_n787));
  MUX2_X1   g362(.A(new_n786), .B(new_n787), .S(KEYINPUT89), .Z(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1341), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n710), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n710), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT87), .B(G1971), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(G288), .A2(KEYINPUT85), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT85), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n583), .A2(new_n795), .A3(new_n584), .A4(new_n585), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G16), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n710), .A2(G23), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT33), .B(G1976), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT86), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n710), .A2(G6), .ZN(new_n804));
  INV_X1    g379(.A(G305), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n710), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n802), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n798), .A2(new_n809), .A3(new_n799), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n793), .A2(new_n803), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT88), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT88), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n814), .A3(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G25), .A2(G29), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n484), .A2(G119), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n476), .A2(G131), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n817), .B1(new_n823), .B2(G29), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT83), .Z(new_n825));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G1991), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n798), .A2(new_n809), .A3(new_n799), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n809), .B1(new_n798), .B2(new_n799), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT34), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n830), .A2(new_n831), .A3(new_n808), .A4(new_n793), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n710), .A2(G24), .ZN(new_n833));
  INV_X1    g408(.A(G290), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n710), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT84), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(KEYINPUT84), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G1986), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(G1986), .A3(new_n837), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n832), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n816), .A2(new_n827), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT36), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n832), .A2(new_n840), .A3(new_n841), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n813), .B2(new_n815), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n845), .B1(new_n847), .B2(new_n827), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n785), .B(new_n789), .C1(new_n844), .C2(new_n848), .ZN(G150));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n850));
  NAND2_X1  g425(.A1(G150), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n843), .B(KEYINPUT36), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n852), .A2(KEYINPUT98), .A3(new_n789), .A4(new_n785), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(G311));
  NAND2_X1  g429(.A1(new_n515), .A2(G55), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT100), .B(G93), .Z(new_n856));
  NAND3_X1  g431(.A1(new_n524), .A2(new_n856), .A3(new_n508), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n857), .C1(new_n858), .C2(new_n526), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  INV_X1    g436(.A(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n562), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n859), .B(new_n556), .C1(new_n560), .C2(new_n561), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n618), .A2(new_n622), .A3(new_n626), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n635), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT39), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n867), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n861), .B1(new_n871), .B2(G860), .ZN(G145));
  XNOR2_X1  g447(.A(new_n643), .B(new_n489), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n742), .B(new_n482), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n873), .B(new_n874), .Z(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n777), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n503), .B(new_n729), .Z(new_n879));
  NAND3_X1  g454(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n503), .B(new_n729), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n754), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n778), .B(new_n878), .C1(new_n881), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n777), .A2(KEYINPUT101), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n754), .A2(new_n882), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n822), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n822), .B1(new_n884), .B2(new_n888), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n484), .A2(G130), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n892), .A2(KEYINPUT102), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(KEYINPUT102), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n893), .A2(new_n894), .B1(G142), .B2(new_n476), .ZN(new_n895));
  OR2_X1    g470(.A1(G106), .A2(G2105), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n896), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n890), .A2(new_n891), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n884), .A2(new_n888), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n823), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n898), .B1(new_n902), .B2(new_n889), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n876), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G37), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n899), .B1(new_n890), .B2(new_n891), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n898), .A3(new_n889), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n875), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n904), .A2(KEYINPUT103), .A3(new_n905), .A4(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT40), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(G395));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n862), .A2(G868), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT104), .B1(new_n574), .B2(new_n580), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n522), .A2(G91), .B1(new_n577), .B2(G651), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n572), .A4(new_n573), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n924), .A3(new_n868), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n627), .A2(new_n581), .A3(new_n923), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT41), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n925), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n865), .B(new_n637), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n925), .A2(new_n926), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(new_n935), .B2(new_n933), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT42), .ZN(new_n937));
  NAND2_X1  g512(.A1(G290), .A2(G303), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n794), .A2(new_n796), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n606), .A2(new_n527), .A3(new_n608), .A4(new_n523), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n938), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(G305), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n938), .A2(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n797), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n805), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n937), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n950));
  INV_X1    g525(.A(new_n948), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n918), .B(new_n920), .C1(new_n954), .C2(new_n610), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n610), .B1(new_n949), .B2(new_n953), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT105), .B1(new_n956), .B2(new_n919), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(G295));
  OAI21_X1  g533(.A(new_n920), .B1(new_n954), .B2(new_n610), .ZN(G331));
  INV_X1    g534(.A(new_n864), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n557), .A2(new_n558), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT72), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n559), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n859), .B1(new_n964), .B2(new_n556), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n548), .A2(G286), .A3(new_n552), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(G286), .B1(new_n548), .B2(new_n552), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n960), .A2(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(G301), .A2(G168), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n863), .A2(new_n864), .A3(new_n970), .A4(new_n966), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n935), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n935), .A2(new_n969), .A3(new_n974), .A4(new_n971), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n865), .B(KEYINPUT106), .C1(new_n968), .C2(new_n967), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n969), .A2(new_n978), .A3(new_n971), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n931), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n948), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT108), .B1(new_n981), .B2(G37), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n979), .A2(new_n977), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n984), .A2(new_n931), .B1(new_n973), .B2(new_n975), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n983), .B(new_n905), .C1(new_n985), .C2(new_n948), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n948), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n982), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n984), .A2(new_n927), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n932), .A2(new_n991), .B1(new_n969), .B2(new_n971), .ZN(new_n993));
  OAI221_X1 g568(.A(new_n951), .B1(new_n991), .B2(new_n928), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(new_n905), .A3(new_n987), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n990), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT44), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n988), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT109), .B1(new_n988), .B2(KEYINPUT43), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n1001), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g577(.A(KEYINPUT126), .B(KEYINPUT46), .Z(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n503), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n477), .A2(G40), .A3(new_n481), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1005), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1003), .B1(new_n1008), .B2(G1996), .ZN(new_n1009));
  INV_X1    g584(.A(G2067), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n729), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1007), .B1(new_n1012), .B2(new_n880), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT126), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1007), .B(new_n1014), .C1(new_n1015), .C2(KEYINPUT46), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1009), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT47), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n880), .B(new_n1014), .ZN(new_n1019));
  AND4_X1   g594(.A1(new_n826), .A2(new_n1019), .A3(new_n823), .A4(new_n1011), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n729), .A2(G2067), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1007), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1011), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n822), .B(new_n826), .Z(new_n1025));
  OAI21_X1  g600(.A(new_n1007), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1007), .A2(new_n839), .A3(new_n834), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1028));
  XNOR2_X1  g603(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1023), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n591), .A2(new_n1031), .A3(new_n595), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n595), .B1(new_n587), .B2(new_n521), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G1981), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1032), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n503), .A2(new_n1004), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(new_n1006), .ZN(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1032), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1032), .B1(new_n1045), .B2(G288), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1041), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G303), .A2(G8), .ZN(new_n1048));
  NAND2_X1  g623(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n504), .A2(new_n1004), .A3(new_n506), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1006), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT112), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1971), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1053), .A2(KEYINPUT50), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1006), .B1(new_n1005), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G2090), .ZN(new_n1066));
  OAI211_X1 g641(.A(G8), .B(new_n1052), .C1(new_n1061), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1006), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1005), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G8), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1044), .B1(new_n794), .B2(new_n796), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT52), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n939), .A2(G1976), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT114), .B(G1976), .Z(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1041), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1043), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1047), .B1(new_n1067), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1072), .A2(new_n1043), .A3(new_n1076), .A4(KEYINPUT116), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1971), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1055), .A2(new_n1059), .A3(new_n1056), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1059), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(KEYINPUT115), .B(new_n1068), .C1(new_n1005), .C2(new_n1063), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n504), .A2(new_n1063), .A3(new_n1004), .A4(new_n506), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1063), .B1(new_n503), .B2(new_n1004), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1006), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1088), .A3(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1092), .A2(G2090), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1040), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1067), .B(new_n1082), .C1(new_n1052), .C2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G2078), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1058), .A2(new_n1096), .A3(new_n1060), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1065), .A2(new_n736), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1006), .B1(new_n1038), .B2(new_n1054), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n1004), .A4(new_n506), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1101), .A2(new_n1102), .A3(KEYINPUT53), .A4(new_n1096), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1099), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G171), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1095), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1107));
  INV_X1    g682(.A(G1966), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G2084), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1062), .A2(new_n1064), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1111), .A3(G168), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT51), .ZN(new_n1114));
  AOI21_X1  g689(.A(G168), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n1116));
  OAI211_X1 g691(.A(G8), .B(new_n1112), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1114), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1078), .B1(new_n1106), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1112), .A2(G8), .A3(G168), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1123), .B1(new_n1095), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(G8), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1052), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1077), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1128), .A2(KEYINPUT63), .A3(new_n1129), .A4(new_n1067), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1122), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  INV_X1    g708(.A(G1348), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1065), .A2(new_n1134), .B1(new_n1010), .B2(new_n1039), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1133), .B1(new_n1135), .B2(new_n868), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1135), .A2(new_n868), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT121), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1092), .A2(new_n762), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1092), .A2(KEYINPUT117), .A3(new_n762), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1057), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(G2072), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1141), .A2(new_n1142), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n574), .B(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n922), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1149), .A2(KEYINPUT119), .A3(new_n1150), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1153), .B(new_n1154), .C1(new_n1150), .C2(G299), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1136), .B(new_n1138), .C1(new_n1146), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1146), .A2(new_n1155), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT61), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1162));
  XNOR2_X1  g737(.A(G301), .B(KEYINPUT54), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1096), .A2(KEYINPUT125), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT53), .B1(new_n1165), .B2(G2078), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1164), .B(new_n1166), .C1(new_n1005), .C2(KEYINPUT45), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1167), .B2(new_n1101), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1099), .A2(new_n1100), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1163), .B2(new_n1104), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1155), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1174), .A2(new_n1175), .B1(KEYINPUT121), .B2(new_n1137), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1176), .A2(KEYINPUT61), .A3(new_n1157), .A4(new_n1136), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1095), .ZN(new_n1178));
  AND4_X1   g753(.A1(new_n1161), .A2(new_n1171), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(KEYINPUT58), .B(G1341), .Z(new_n1180));
  AND2_X1   g755(.A1(new_n1069), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1143), .A2(KEYINPUT122), .A3(new_n1014), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(new_n1057), .B2(G1996), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1181), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g762(.A(KEYINPUT123), .B(new_n1181), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n563), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1135), .A2(KEYINPUT60), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(new_n627), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1193), .B1(KEYINPUT60), .B2(new_n1135), .ZN(new_n1194));
  OAI211_X1 g769(.A(KEYINPUT59), .B(new_n563), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1191), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1158), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1132), .B1(new_n1179), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1007), .A2(G1986), .A3(G290), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1027), .A2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT111), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1026), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1030), .B1(new_n1198), .B2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g778(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n1205));
  INV_X1    g779(.A(KEYINPUT109), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OR2_X1    g781(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1208));
  NAND3_X1  g782(.A1(new_n988), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n1209));
  NAND3_X1  g783(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g784(.A(new_n687), .B1(new_n666), .B2(new_n667), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1211), .B1(new_n911), .B2(new_n912), .ZN(new_n1212));
  NOR2_X1   g786(.A1(G229), .A2(new_n466), .ZN(new_n1213));
  AND3_X1   g787(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(G308));
  NAND3_X1  g788(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(G225));
endmodule


