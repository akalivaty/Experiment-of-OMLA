//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  XOR2_X1   g000(.A(KEYINPUT21), .B(G898), .Z(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT90), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  OAI211_X1 g004(.A(G902), .B(G953), .C1(new_n189), .C2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT89), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G952), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n189), .B2(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(G214), .B1(G237), .B2(G902), .ZN(new_n198));
  XOR2_X1   g012(.A(new_n198), .B(KEYINPUT81), .Z(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(G210), .B1(G237), .B2(G902), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT78), .A3(G104), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n203), .A2(KEYINPUT78), .A3(KEYINPUT3), .A4(G104), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n203), .A2(G104), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT4), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G101), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT2), .B(G113), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT67), .A2(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT67), .A2(G119), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(G116), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G119), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n215), .B(new_n218), .C1(G116), .C2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT67), .A2(G119), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT67), .A2(G119), .ZN(new_n222));
  INV_X1    g036(.A(G116), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n219), .A2(G116), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n214), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n213), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n209), .A2(G101), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n208), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT4), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n208), .B2(new_n210), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n229), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n211), .A2(G101), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n212), .B1(new_n208), .B2(new_n230), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(KEYINPUT79), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n228), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n218), .B(KEYINPUT5), .C1(G116), .C2(new_n219), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT5), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n224), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(G113), .A3(new_n242), .ZN(new_n243));
  XOR2_X1   g057(.A(G104), .B(G107), .Z(new_n244));
  AOI22_X1  g058(.A1(new_n208), .A2(new_n230), .B1(G101), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n220), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G110), .B(G122), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n239), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n248), .B(KEYINPUT8), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n245), .B1(new_n243), .B2(new_n220), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT65), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n257), .A3(G143), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n258), .A2(new_n259), .A3(G128), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n254), .A2(G143), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n255), .A2(new_n257), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(new_n260), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n262), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G125), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(G143), .B1(new_n255), .B2(new_n257), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n266), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n258), .A2(new_n261), .A3(new_n272), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(G125), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n194), .A2(G224), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT7), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n271), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n253), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n250), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n280), .B1(new_n271), .B2(new_n278), .ZN(new_n286));
  OAI22_X1  g100(.A1(new_n286), .A2(KEYINPUT83), .B1(new_n281), .B2(new_n282), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n286), .A2(KEYINPUT83), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n232), .A2(new_n229), .A3(new_n234), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT79), .B1(new_n236), .B2(new_n237), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n246), .B(new_n248), .C1(new_n293), .C2(new_n228), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n249), .B1(new_n239), .B2(new_n247), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT6), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT6), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n249), .C1(new_n239), .C2(new_n247), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n271), .A2(new_n278), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(new_n279), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n202), .B1(new_n290), .B2(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n290), .A2(new_n301), .A3(new_n202), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT84), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n290), .A2(new_n301), .A3(new_n202), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT84), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n201), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G113), .B(G122), .ZN(new_n309));
  INV_X1    g123(.A(G104), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n190), .A2(KEYINPUT68), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G237), .ZN(new_n314));
  AOI21_X1  g128(.A(G953), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G214), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n260), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(G143), .A3(G214), .ZN(new_n318));
  INV_X1    g132(.A(G131), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT18), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n270), .A2(G140), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT65), .B(G146), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n254), .B2(new_n326), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n315), .A2(G143), .A3(G214), .ZN(new_n330));
  AOI21_X1  g144(.A(G143), .B1(new_n315), .B2(G214), .ZN(new_n331));
  OAI21_X1  g145(.A(G131), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n322), .B(new_n329), .C1(new_n321), .C2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n317), .A2(new_n319), .A3(new_n318), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(KEYINPUT17), .B(G131), .C1(new_n330), .C2(new_n331), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT73), .A4(KEYINPUT16), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT16), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT73), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n324), .B2(KEYINPUT16), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n339), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n338), .B1(new_n343), .B2(G146), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(G146), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT16), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n346), .B(new_n341), .C1(KEYINPUT16), .C2(new_n324), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(KEYINPUT74), .A3(new_n254), .A4(new_n339), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n337), .A2(new_n344), .A3(new_n345), .A4(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n311), .B(new_n333), .C1(new_n336), .C2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT86), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n344), .A2(new_n345), .A3(new_n348), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n337), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n355), .A2(KEYINPUT86), .A3(new_n311), .A4(new_n333), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n332), .A2(new_n334), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n326), .B(KEYINPUT19), .Z(new_n359));
  OAI21_X1  g173(.A(new_n345), .B1(new_n359), .B2(new_n267), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n333), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n311), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n365));
  NOR2_X1   g179(.A1(G475), .A2(G902), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n352), .A2(new_n356), .B1(new_n361), .B2(new_n362), .ZN(new_n368));
  INV_X1    g182(.A(new_n366), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT20), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT70), .B(G217), .Z(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT9), .B(G234), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n372), .A2(G953), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n223), .A2(G122), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT14), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT88), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n375), .A2(KEYINPUT14), .ZN(new_n379));
  OR3_X1    g193(.A1(new_n223), .A2(KEYINPUT87), .A3(G122), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT87), .B1(new_n223), .B2(G122), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n203), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n381), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n203), .A3(new_n375), .ZN(new_n385));
  XNOR2_X1  g199(.A(G128), .B(G143), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n386), .A2(G134), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(G134), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n375), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G107), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n391), .A2(new_n385), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT13), .B1(new_n263), .B2(G143), .ZN(new_n393));
  INV_X1    g207(.A(G134), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n395), .A2(new_n386), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n386), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI221_X1 g212(.A(new_n374), .B1(new_n383), .B2(new_n389), .C1(new_n392), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n374), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n383), .A2(new_n389), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n391), .A2(new_n385), .B1(new_n396), .B2(new_n397), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(G902), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G478), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(KEYINPUT15), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n404), .A2(new_n407), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n355), .A2(new_n333), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n352), .A2(new_n356), .B1(new_n362), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G475), .B1(new_n412), .B2(G902), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n371), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G221), .B1(new_n373), .B2(G902), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n276), .A2(new_n277), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n212), .B2(new_n234), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n291), .B2(new_n292), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n269), .A2(new_n245), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT10), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT10), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT80), .B1(new_n266), .B2(new_n259), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n259), .B1(G143), .B2(new_n254), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT80), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n263), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n422), .A2(new_n425), .B1(new_n258), .B2(new_n261), .ZN(new_n426));
  INV_X1    g240(.A(new_n262), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n421), .B(new_n245), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n420), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT11), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n394), .B2(G137), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n394), .A2(G137), .ZN(new_n432));
  INV_X1    g246(.A(G137), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT11), .A3(G134), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G131), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n431), .A2(new_n434), .A3(new_n319), .A4(new_n432), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n418), .A2(new_n429), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n245), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n265), .B1(new_n327), .B2(G143), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n259), .B1(new_n327), .B2(G143), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(new_n263), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n443), .A3(new_n262), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n245), .B1(new_n426), .B2(new_n427), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n436), .A2(new_n437), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT12), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT12), .ZN(new_n449));
  AOI211_X1 g263(.A(new_n449), .B(new_n438), .C1(new_n444), .C2(new_n445), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n439), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G140), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n194), .A2(G227), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n235), .A2(new_n238), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n456), .A2(new_n417), .B1(new_n420), .B2(new_n428), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n457), .B2(new_n438), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n418), .A2(new_n429), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n447), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(G469), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(G469), .A2(G902), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n418), .A2(new_n429), .A3(new_n438), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n438), .B1(new_n418), .B2(new_n429), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n454), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n454), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n439), .B(new_n468), .C1(new_n448), .C2(new_n450), .ZN(new_n469));
  AOI211_X1 g283(.A(G469), .B(G902), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n415), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n414), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT32), .ZN(new_n473));
  INV_X1    g287(.A(new_n432), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n394), .A2(G137), .ZN(new_n475));
  OAI21_X1  g289(.A(G131), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n437), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n269), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n447), .A2(new_n276), .A3(new_n277), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n477), .B1(new_n443), .B2(new_n262), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n416), .A2(KEYINPUT66), .B1(new_n437), .B2(new_n436), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n276), .A2(new_n484), .A3(new_n277), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n227), .B(new_n481), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n227), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n479), .A2(new_n490), .A3(new_n480), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n315), .A2(G210), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT27), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT27), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n315), .A2(new_n494), .A3(G210), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT26), .B(G101), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n493), .B2(new_n495), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n491), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT31), .ZN(new_n501));
  INV_X1    g315(.A(new_n416), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n502), .A2(new_n447), .B1(new_n269), .B2(new_n478), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(new_n490), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n491), .A2(KEYINPUT28), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n276), .A2(new_n484), .A3(new_n277), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n484), .B1(new_n276), .B2(new_n277), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n508), .A2(new_n509), .A3(new_n438), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n227), .B1(new_n510), .B2(new_n482), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n499), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT31), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n489), .A2(new_n515), .A3(new_n491), .A4(new_n499), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n501), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(G472), .A2(G902), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n473), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n517), .A2(new_n473), .A3(new_n518), .ZN(new_n520));
  INV_X1    g334(.A(G472), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n499), .B1(new_n490), .B2(new_n503), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT29), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n489), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G902), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n504), .B1(new_n503), .B2(new_n490), .ZN(new_n527));
  AND4_X1   g341(.A1(new_n504), .A2(new_n479), .A3(new_n490), .A4(new_n480), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n511), .B(new_n523), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n503), .A2(new_n490), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(new_n506), .B2(new_n505), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n529), .B(new_n499), .C1(new_n531), .C2(new_n523), .ZN(new_n532));
  AOI211_X1 g346(.A(KEYINPUT69), .B(new_n521), .C1(new_n526), .C2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n529), .A2(new_n499), .ZN(new_n535));
  INV_X1    g349(.A(new_n530), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n523), .B1(new_n507), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n525), .B(new_n524), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n534), .B1(new_n538), .B2(G472), .ZN(new_n539));
  OAI22_X1  g353(.A1(new_n519), .A2(new_n520), .B1(new_n533), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n372), .B1(G234), .B2(new_n525), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n263), .B1(new_n221), .B2(new_n222), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT23), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(KEYINPUT23), .A2(G119), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT72), .B1(new_n546), .B2(G128), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT72), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n548), .A2(new_n263), .A3(KEYINPUT23), .A4(G119), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n216), .A2(G128), .A3(new_n217), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n545), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G110), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT71), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n216), .A2(new_n554), .A3(G128), .A4(new_n217), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n221), .A2(new_n222), .A3(new_n263), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT71), .B1(new_n219), .B2(G128), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT24), .B(G110), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G110), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n545), .A2(new_n550), .A3(new_n563), .A4(new_n551), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT75), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n559), .B(new_n555), .C1(new_n556), .C2(new_n557), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n345), .A3(new_n328), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n569));
  OAI22_X1  g383(.A1(new_n353), .A2(new_n562), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT76), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n344), .A2(new_n345), .A3(new_n348), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n553), .A3(new_n561), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT76), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n573), .B(new_n574), .C1(new_n569), .C2(new_n568), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT22), .B(G137), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT77), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n571), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n570), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n578), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n525), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n580), .A2(KEYINPUT25), .A3(new_n525), .A4(new_n582), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n542), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n580), .A2(new_n582), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n541), .A2(G902), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n308), .A2(new_n472), .A3(new_n540), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  NOR3_X1   g408(.A1(new_n471), .A2(new_n587), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n517), .A2(new_n525), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n517), .A2(new_n518), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT92), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n368), .A2(KEYINPUT20), .A3(new_n369), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n413), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n404), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(KEYINPUT91), .A3(new_n405), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT91), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n404), .B2(G478), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n399), .A2(new_n403), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT33), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n399), .A2(new_n612), .A3(new_n403), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n405), .A2(G902), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n607), .A2(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n605), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n197), .B(new_n200), .C1(new_n303), .C2(new_n302), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n602), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n616), .B1(new_n371), .B2(new_n413), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n290), .A2(new_n301), .ZN(new_n622));
  INV_X1    g436(.A(new_n202), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n199), .B1(new_n624), .B2(new_n306), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n621), .A2(new_n625), .A3(KEYINPUT92), .A4(new_n197), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n601), .B1(new_n620), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT34), .B(G104), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  INV_X1    g443(.A(new_n410), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n371), .A2(new_n630), .A3(new_n413), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n619), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n595), .A3(new_n600), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  OR2_X1    g449(.A1(new_n579), .A2(KEYINPUT36), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n636), .A2(KEYINPUT93), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(KEYINPUT93), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n571), .ZN(new_n640));
  INV_X1    g454(.A(new_n575), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n637), .A2(new_n571), .A3(new_n575), .A4(new_n638), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n642), .A2(new_n643), .A3(new_n589), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n587), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n308), .A2(new_n472), .A3(new_n600), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT94), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT37), .B(G110), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  INV_X1    g463(.A(new_n196), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n192), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n631), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n200), .B1(new_n303), .B2(new_n302), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n471), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n653), .A2(new_n655), .A3(new_n540), .A4(new_n645), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  INV_X1    g471(.A(new_n415), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n451), .A2(new_n454), .B1(new_n458), .B2(new_n460), .ZN(new_n659));
  OAI21_X1  g473(.A(G469), .B1(new_n659), .B2(G902), .ZN(new_n660));
  INV_X1    g474(.A(G469), .ZN(new_n661));
  INV_X1    g475(.A(new_n467), .ZN(new_n662));
  INV_X1    g476(.A(new_n469), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n661), .B(new_n525), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n658), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n652), .B(KEYINPUT39), .Z(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT40), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT96), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n290), .A2(new_n301), .A3(new_n304), .A4(new_n202), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n307), .A2(new_n671), .A3(new_n624), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n587), .A2(new_n644), .ZN(new_n675));
  AOI21_X1  g489(.A(G902), .B1(new_n536), .B2(new_n522), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n513), .B1(new_n489), .B2(new_n491), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n520), .B2(new_n519), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n674), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n670), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n411), .A2(new_n362), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n357), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n525), .ZN(new_n685));
  AOI22_X1  g499(.A1(new_n367), .A2(new_n370), .B1(new_n685), .B2(G475), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n410), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n200), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n668), .B2(new_n669), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT97), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT97), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n682), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n260), .ZN(G45));
  AOI211_X1 g509(.A(new_n616), .B(new_n652), .C1(new_n371), .C2(new_n413), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n655), .A2(new_n696), .A3(new_n540), .A4(new_n645), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT98), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n675), .A2(new_n654), .A3(new_n471), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(KEYINPUT98), .A3(new_n540), .A4(new_n696), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT99), .B(G146), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G48));
  NAND2_X1  g518(.A1(new_n620), .A2(new_n626), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n467), .A2(new_n469), .ZN(new_n706));
  OAI21_X1  g520(.A(G469), .B1(new_n706), .B2(G902), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n415), .A3(new_n664), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n540), .A2(new_n709), .A3(new_n592), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT100), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT100), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n705), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND4_X1  g531(.A1(new_n632), .A2(new_n540), .A3(new_n592), .A4(new_n709), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NOR2_X1   g533(.A1(new_n619), .A2(new_n708), .ZN(new_n720));
  INV_X1    g534(.A(new_n414), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n540), .A3(new_n721), .A4(new_n645), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  NAND2_X1  g537(.A1(new_n585), .A2(new_n586), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n541), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n590), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT101), .B1(new_n587), .B2(new_n591), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n501), .B(new_n516), .C1(new_n499), .C2(new_n531), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n518), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n597), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n720), .A2(new_n687), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n736), .B(G122), .Z(G24));
  NOR2_X1   g551(.A1(new_n708), .A2(new_n654), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n696), .A3(new_n733), .A4(new_n645), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  AND3_X1   g554(.A1(new_n307), .A2(new_n671), .A3(new_n624), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT102), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n200), .A4(new_n665), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n307), .A2(new_n624), .A3(new_n671), .A4(new_n200), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT102), .B1(new_n744), .B2(new_n471), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n726), .B1(new_n725), .B2(new_n590), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n587), .A2(new_n591), .A3(KEYINPUT101), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n540), .B(new_n696), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT42), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n696), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(KEYINPUT42), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n540), .A2(new_n592), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n745), .A4(new_n743), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  NAND4_X1  g570(.A1(new_n753), .A2(new_n743), .A3(new_n653), .A4(new_n745), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NAND2_X1  g572(.A1(new_n686), .A2(new_n617), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n686), .A2(new_n761), .A3(new_n617), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n760), .A2(new_n599), .A3(new_n645), .A4(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(KEYINPUT44), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n744), .B(KEYINPUT105), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n766), .A2(KEYINPUT106), .A3(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n659), .A2(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n659), .A2(KEYINPUT45), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(G469), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n463), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT104), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n463), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT103), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(new_n664), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT104), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n773), .A2(new_n780), .A3(new_n774), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n776), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n778), .B1(new_n777), .B2(new_n664), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n415), .B(new_n666), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n769), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT106), .B1(new_n766), .B2(new_n768), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  OAI21_X1  g602(.A(new_n415), .B1(new_n782), .B2(new_n783), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT47), .B(new_n415), .C1(new_n782), .C2(new_n783), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n751), .A2(new_n540), .A3(new_n592), .A4(new_n744), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT107), .B(G140), .Z(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G42));
  NAND2_X1  g611(.A1(new_n707), .A2(new_n664), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n199), .B(new_n658), .C1(new_n798), .C2(KEYINPUT49), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(KEYINPUT49), .B2(new_n798), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n680), .A3(new_n759), .ZN(new_n801));
  INV_X1    g615(.A(new_n674), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n729), .ZN(new_n803));
  INV_X1    g617(.A(new_n409), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n404), .A2(new_n407), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT108), .B1(new_n408), .B2(new_n409), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n371), .A2(new_n809), .A3(new_n413), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n618), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n595), .A3(new_n308), .A4(new_n600), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n593), .A3(new_n646), .A4(new_n722), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n718), .B1(new_n734), .B2(new_n735), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n605), .A2(new_n652), .A3(new_n809), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n744), .A2(new_n471), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n540), .A4(new_n645), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n675), .A2(new_n732), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n743), .A2(new_n820), .A3(new_n745), .A4(new_n696), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n757), .A2(new_n819), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n755), .A2(new_n715), .A3(new_n815), .A4(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n757), .A2(new_n819), .A3(new_n821), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT109), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n654), .A2(new_n686), .A3(new_n410), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n471), .A2(new_n652), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n675), .A3(new_n680), .A4(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n831), .A2(new_n656), .A3(new_n739), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n832), .A2(new_n702), .A3(KEYINPUT112), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT112), .B1(new_n832), .B2(new_n702), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT52), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n699), .A2(new_n701), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n831), .A2(new_n739), .A3(new_n656), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(new_n702), .A3(KEYINPUT112), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n828), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n824), .A2(new_n827), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT113), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n833), .A2(new_n834), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n836), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n840), .A2(new_n849), .A3(new_n836), .A4(new_n841), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n832), .A2(new_n702), .A3(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT111), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT111), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n832), .A2(new_n702), .A3(new_n855), .A4(KEYINPUT52), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n848), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n845), .A2(new_n846), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n707), .A2(new_n658), .A3(new_n664), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n791), .A2(new_n792), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n760), .A2(new_n650), .A3(new_n762), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n864), .A2(new_n733), .A3(new_n729), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n865), .A2(new_n767), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n744), .A2(new_n708), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n864), .A2(new_n820), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n680), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n870), .A2(new_n872), .A3(new_n592), .A4(new_n650), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n686), .A2(new_n616), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n708), .A2(new_n200), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n802), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n802), .A2(KEYINPUT117), .A3(new_n876), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n865), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT50), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n879), .A2(new_n865), .A3(KEYINPUT50), .A4(new_n880), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n875), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n869), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n867), .A2(new_n868), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n861), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n195), .B1(new_n873), .B2(new_n618), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n864), .A2(new_n540), .A3(new_n729), .A4(new_n870), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT48), .Z(new_n891));
  AOI211_X1 g705(.A(new_n889), .B(new_n891), .C1(new_n738), .C2(new_n865), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n861), .B(new_n875), .C1(new_n883), .C2(new_n884), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n863), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n791), .A2(KEYINPUT118), .A3(new_n792), .A4(new_n862), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n866), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n893), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n893), .B2(new_n897), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n888), .B(new_n892), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n851), .A2(new_n858), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n755), .A2(new_n715), .A3(new_n815), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT110), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n826), .A4(new_n823), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT110), .B1(new_n824), .B2(new_n827), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n847), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT114), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT114), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n910), .B(new_n847), .C1(new_n902), .C2(new_n907), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n843), .A2(new_n844), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n909), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n860), .B(new_n901), .C1(new_n914), .C2(KEYINPUT54), .ZN(new_n915));
  NOR2_X1   g729(.A1(G952), .A2(G953), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n803), .B1(new_n915), .B2(new_n916), .ZN(G75));
  NOR2_X1   g731(.A1(new_n194), .A2(G952), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT120), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n525), .B1(new_n845), .B2(new_n859), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(G210), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n296), .A2(new_n298), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n300), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT55), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n929), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n920), .B1(new_n930), .B2(new_n931), .ZN(G51));
  XOR2_X1   g746(.A(new_n463), .B(KEYINPUT57), .Z(new_n933));
  AOI21_X1  g747(.A(new_n846), .B1(new_n845), .B2(new_n859), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n860), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n706), .ZN(new_n938));
  OAI211_X1 g752(.A(KEYINPUT121), .B(new_n933), .C1(new_n860), .C2(new_n934), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n923), .A2(new_n772), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n918), .B1(new_n940), .B2(new_n941), .ZN(G54));
  NAND2_X1  g756(.A1(KEYINPUT58), .A2(G475), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT122), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n922), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n368), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n364), .B1(new_n922), .B2(new_n944), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n946), .A2(new_n918), .A3(new_n947), .ZN(G60));
  NAND2_X1  g762(.A1(G478), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT59), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n614), .B(new_n951), .C1(new_n860), .C2(new_n934), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n919), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n912), .B1(new_n908), .B2(KEYINPUT114), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n846), .B1(new_n954), .B2(new_n911), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n951), .B1(new_n955), .B2(new_n860), .ZN(new_n956));
  INV_X1    g770(.A(new_n614), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G63));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n845), .B2(new_n859), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n642), .A2(new_n643), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n920), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n959), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n962), .A2(new_n588), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n967), .B(new_n964), .C1(new_n965), .C2(new_n959), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G66));
  INV_X1    g785(.A(G224), .ZN(new_n972));
  OAI21_X1  g786(.A(G953), .B1(new_n188), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT125), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n715), .A2(new_n815), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n974), .B1(new_n979), .B2(G953), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n926), .B1(G898), .B2(new_n194), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G69));
  OAI21_X1  g796(.A(new_n481), .B1(new_n486), .B2(new_n488), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(new_n359), .ZN(new_n984));
  NAND2_X1  g798(.A1(G900), .A2(G953), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n729), .A2(new_n540), .A3(new_n829), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n784), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n702), .A2(new_n656), .A3(new_n739), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n987), .A2(new_n757), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n787), .A2(new_n755), .A3(new_n795), .A4(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n984), .B(new_n985), .C1(new_n990), .C2(G953), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n691), .A2(new_n992), .A3(new_n693), .A4(new_n988), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n753), .A2(new_n666), .A3(new_n818), .A4(new_n811), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n787), .A2(new_n795), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n691), .A2(new_n693), .A3(new_n988), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(KEYINPUT126), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n991), .B1(new_n1001), .B2(new_n984), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1003), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n991), .B(new_n1005), .C1(new_n1001), .C2(new_n984), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(new_n990), .B2(new_n978), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n489), .A2(new_n522), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n918), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1009), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n1000), .B2(new_n979), .ZN(new_n1014));
  INV_X1    g828(.A(new_n678), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1011), .A2(new_n678), .A3(new_n1013), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n914), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n914), .A2(KEYINPUT127), .A3(new_n1017), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1016), .B1(new_n1020), .B2(new_n1021), .ZN(G57));
endmodule


