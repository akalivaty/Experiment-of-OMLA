//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n189));
  INV_X1    g003(.A(G101), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n193), .A2(KEYINPUT3), .A3(G104), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT3), .B1(new_n193), .B2(G104), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n190), .B(new_n192), .C1(new_n194), .C2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT74), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n191), .B2(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n193), .A2(KEYINPUT3), .A3(G104), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n200), .A2(new_n201), .B1(new_n191), .B2(G107), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n198), .B1(new_n202), .B2(new_n190), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT75), .B1(new_n193), .B2(G104), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT75), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(new_n191), .A3(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n193), .A2(G104), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n208), .A2(KEYINPUT76), .A3(G101), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT76), .B1(new_n208), .B2(G101), .ZN(new_n210));
  OAI22_X1  g024(.A1(new_n197), .A2(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n212), .A2(G143), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n216), .A2(new_n217), .B1(KEYINPUT1), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT10), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT4), .B1(new_n202), .B2(new_n190), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n202), .A2(new_n198), .A3(new_n190), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n196), .A2(KEYINPUT74), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n230), .A2(new_n213), .A3(new_n215), .ZN(new_n231));
  OR2_X1    g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n216), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n231), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G101), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n216), .A2(KEYINPUT64), .A3(new_n229), .A4(new_n232), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OAI22_X1  g054(.A1(new_n211), .A2(new_n224), .B1(new_n228), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n208), .A2(G101), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT76), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n208), .A2(KEYINPUT76), .A3(G101), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n244), .A2(new_n245), .B1(new_n227), .B2(new_n226), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n222), .A2(KEYINPUT77), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT77), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n220), .A2(new_n248), .A3(new_n221), .A4(G128), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n219), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT10), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n189), .B1(new_n241), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT11), .B1(new_n253), .B2(G137), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n256), .B2(G134), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(KEYINPUT65), .A3(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G131), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n258), .A2(new_n264), .A3(new_n260), .A4(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT10), .ZN(new_n267));
  INV_X1    g081(.A(new_n250), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n211), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n246), .A2(KEYINPUT10), .A3(new_n223), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n227), .A2(new_n226), .ZN(new_n271));
  INV_X1    g085(.A(new_n225), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n232), .A2(new_n229), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n234), .B1(new_n274), .B2(new_n220), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n220), .A2(new_n230), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n239), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(new_n278), .A3(new_n238), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n269), .A2(new_n270), .A3(new_n279), .A4(KEYINPUT80), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n252), .A2(new_n266), .A3(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n241), .A2(new_n251), .A3(new_n266), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G110), .B(G140), .ZN(new_n285));
  INV_X1    g099(.A(G953), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n286), .A2(G227), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n285), .B(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(KEYINPUT81), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n282), .A2(new_n288), .ZN(new_n290));
  XOR2_X1   g104(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n291));
  NAND2_X1  g105(.A1(new_n244), .A2(new_n245), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n292), .A2(new_n271), .A3(new_n250), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n223), .B1(new_n292), .B2(new_n271), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n266), .B(new_n291), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n266), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n246), .A2(new_n250), .ZN(new_n297));
  INV_X1    g111(.A(new_n223), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n211), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n295), .B(KEYINPUT79), .C1(new_n300), .C2(KEYINPUT12), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n302), .A3(new_n291), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n290), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n289), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT81), .B1(new_n284), .B2(new_n288), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n187), .B(new_n188), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n301), .A2(new_n283), .A3(new_n303), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n308), .A2(new_n288), .B1(new_n281), .B2(new_n290), .ZN(new_n309));
  OAI21_X1  g123(.A(G469), .B1(new_n309), .B2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT99), .ZN(new_n312));
  XNOR2_X1  g126(.A(G113), .B(G122), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT90), .B(G104), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(G237), .A2(G953), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(G143), .A3(G214), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(G143), .B1(new_n316), .B2(G214), .ZN(new_n319));
  OAI211_X1 g133(.A(KEYINPUT18), .B(G131), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G146), .ZN(new_n326));
  XNOR2_X1  g140(.A(G125), .B(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n212), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n319), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT18), .A2(G131), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n317), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n320), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT88), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT88), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n320), .A2(new_n332), .A3(new_n329), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT16), .ZN(new_n338));
  OR3_X1    g152(.A1(new_n323), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n338), .A2(G146), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G131), .B1(new_n318), .B2(new_n319), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n330), .A2(new_n264), .A3(new_n317), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n327), .A2(KEYINPUT89), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT19), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n343), .B1(new_n345), .B2(G146), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n315), .B1(new_n337), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n264), .B1(new_n330), .B2(new_n317), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT92), .A3(KEYINPUT17), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT92), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT17), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n341), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n338), .A2(new_n339), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n212), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n338), .A2(new_n339), .A3(G146), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n349), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(G146), .B1(new_n338), .B2(new_n339), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT91), .B1(new_n340), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n341), .A2(new_n342), .A3(new_n351), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n359), .A2(new_n364), .B1(new_n336), .B2(new_n334), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n347), .B1(new_n365), .B2(new_n315), .ZN(new_n366));
  NOR2_X1   g180(.A1(G475), .A2(G902), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT93), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT20), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n347), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n337), .B(new_n315), .C1(new_n358), .C2(new_n363), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n373));
  INV_X1    g187(.A(new_n368), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n337), .B1(new_n358), .B2(new_n363), .ZN(new_n377));
  INV_X1    g191(.A(new_n315), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n379), .A2(KEYINPUT94), .A3(new_n371), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT94), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n381), .A3(new_n378), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n188), .ZN(new_n383));
  OAI21_X1  g197(.A(G475), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n376), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G478), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT15), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT9), .B(G234), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n388), .A2(new_n389), .A3(G953), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n214), .A2(G128), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n217), .A2(G143), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n253), .ZN(new_n394));
  XNOR2_X1  g208(.A(G116), .B(G122), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n395), .A2(new_n193), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n193), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n214), .A2(KEYINPUT13), .A3(G128), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(KEYINPUT96), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n214), .A2(G128), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n401), .B2(KEYINPUT96), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n217), .A2(G143), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n403), .A2(KEYINPUT95), .A3(KEYINPUT13), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT13), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n405), .B1(new_n392), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n400), .B(new_n402), .C1(new_n404), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n398), .B1(new_n408), .B2(G134), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n395), .A2(new_n193), .ZN(new_n410));
  INV_X1    g224(.A(new_n394), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n253), .B1(new_n392), .B2(new_n393), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G116), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT14), .A3(G122), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G107), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n417), .B2(new_n395), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n391), .B1(new_n409), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n419), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n408), .A2(G134), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n421), .B(new_n390), .C1(new_n422), .C2(new_n398), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT97), .B1(new_n424), .B2(new_n188), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT97), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n426), .B(G902), .C1(new_n420), .C2(new_n423), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n387), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n188), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n426), .ZN(new_n430));
  INV_X1    g244(.A(new_n387), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(G234), .A2(G237), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n433), .A2(G952), .A3(new_n286), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(G898), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(G902), .A3(G953), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n439), .B(KEYINPUT98), .Z(new_n440));
  NAND3_X1  g254(.A1(new_n428), .A2(new_n432), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n312), .B1(new_n385), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n428), .A2(new_n440), .A3(new_n432), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n443), .A2(KEYINPUT99), .A3(new_n384), .A4(new_n376), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G221), .B1(new_n388), .B2(G902), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n311), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n450));
  OR3_X1    g264(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(KEYINPUT2), .A2(G113), .ZN(new_n454));
  INV_X1    g268(.A(G119), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G116), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n414), .A2(G119), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n453), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT5), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT5), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n455), .A3(G116), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n462), .A2(KEYINPUT82), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(KEYINPUT82), .ZN(new_n464));
  OAI211_X1 g278(.A(G113), .B(new_n460), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n459), .B1(new_n465), .B2(KEYINPUT83), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n465), .A2(KEYINPUT83), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n211), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n453), .A2(new_n454), .A3(new_n458), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT82), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n462), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n460), .A2(G113), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT84), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n465), .A2(KEYINPUT84), .A3(new_n469), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n246), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G122), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(KEYINPUT8), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n468), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n277), .A2(G125), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n219), .A2(new_n323), .A3(new_n222), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n286), .A2(G224), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n483), .A2(KEYINPUT7), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n480), .A2(new_n487), .A3(KEYINPUT85), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n453), .A2(new_n454), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(new_n458), .Z(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n273), .A3(new_n238), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n246), .A2(new_n466), .A3(new_n467), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n478), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT85), .B1(new_n480), .B2(new_n487), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n450), .B(new_n188), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n492), .ZN(new_n497));
  INV_X1    g311(.A(new_n478), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n493), .A3(KEYINPUT6), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n481), .A2(new_n482), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n503), .B(new_n483), .Z(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n480), .A2(new_n487), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT85), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n493), .A3(new_n488), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n450), .B1(new_n510), .B2(new_n188), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n449), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n188), .B1(new_n494), .B2(new_n495), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT86), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n515), .A2(new_n448), .A3(new_n505), .A4(new_n496), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G214), .B1(G237), .B2(G902), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n506), .A2(new_n511), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(KEYINPUT87), .A3(new_n448), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT22), .B(G137), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n286), .A2(G221), .A3(G234), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n455), .B2(G128), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n455), .A2(G128), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT70), .B(G110), .Z(new_n532));
  XOR2_X1   g346(.A(KEYINPUT24), .B(G110), .Z(new_n533));
  XNOR2_X1  g347(.A(G119), .B(G128), .ZN(new_n534));
  OAI22_X1  g348(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n356), .A3(new_n328), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n534), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n340), .B2(new_n360), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(KEYINPUT69), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n528), .A2(new_n529), .A3(new_n540), .A4(new_n530), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n539), .A2(G110), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT71), .B(new_n536), .C1(new_n538), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n354), .A2(new_n356), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n539), .A2(G110), .A3(new_n541), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n537), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT71), .B1(new_n547), .B2(new_n536), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n526), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n536), .B1(new_n538), .B2(new_n542), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n525), .ZN(new_n551));
  AOI21_X1  g365(.A(G902), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n522), .B1(new_n552), .B2(KEYINPUT25), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT71), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n525), .B1(new_n555), .B2(new_n543), .ZN(new_n556));
  INV_X1    g370(.A(new_n551), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT25), .B(new_n188), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n188), .B1(new_n556), .B2(new_n557), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT25), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(KEYINPUT72), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n549), .A2(new_n551), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n564), .A2(KEYINPUT73), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n553), .A2(new_n560), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n389), .B1(G234), .B2(new_n188), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(G902), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G472), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n253), .A2(G137), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n256), .A2(G134), .ZN(new_n574));
  OAI21_X1  g388(.A(G131), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n265), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n266), .A2(new_n278), .B1(new_n576), .B2(new_n223), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n489), .B(new_n458), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT28), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n277), .B1(new_n265), .B2(new_n263), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n223), .A2(new_n265), .A3(new_n575), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n490), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n265), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n260), .A2(new_n261), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n264), .B1(new_n584), .B2(new_n258), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n235), .B(new_n239), .C1(new_n583), .C2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n223), .A2(new_n265), .A3(new_n575), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n578), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n579), .B1(new_n589), .B2(KEYINPUT28), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n316), .A2(G210), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT27), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT26), .B(G101), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT29), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT30), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n586), .A2(new_n597), .A3(new_n587), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n586), .B2(new_n587), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n490), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n588), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n596), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n595), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n578), .B1(new_n586), .B2(new_n587), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT28), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n579), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT29), .A4(new_n594), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT68), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n590), .A2(KEYINPUT68), .A3(KEYINPUT29), .A4(new_n594), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n572), .B1(new_n604), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n600), .A2(KEYINPUT31), .A3(new_n594), .A4(new_n588), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n614), .A2(new_n188), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT28), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n582), .B2(new_n588), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n596), .B1(new_n617), .B2(new_n579), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n600), .A2(new_n594), .A3(new_n588), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT31), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n615), .A2(new_n621), .A3(KEYINPUT32), .A4(new_n572), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n615), .A2(new_n572), .A3(new_n621), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT67), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT32), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n615), .A2(new_n621), .A3(KEYINPUT67), .A4(new_n572), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n571), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n447), .A2(new_n521), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  INV_X1    g447(.A(new_n446), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n307), .B2(new_n310), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n568), .A2(new_n570), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n614), .A2(new_n188), .ZN(new_n638));
  OAI21_X1  g452(.A(G472), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n627), .A2(new_n629), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n635), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n518), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n386), .A2(G902), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n424), .A2(KEYINPUT100), .A3(KEYINPUT33), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT33), .B1(new_n424), .B2(KEYINPUT100), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n429), .A2(new_n386), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT20), .B(new_n368), .C1(new_n370), .C2(new_n371), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(G475), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n382), .A2(new_n188), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n379), .A2(KEYINPUT94), .A3(new_n371), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n440), .B(new_n649), .C1(new_n652), .C2(new_n656), .ZN(new_n657));
  AOI211_X1 g471(.A(new_n643), .B(new_n657), .C1(new_n512), .C2(new_n516), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n642), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G104), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT101), .B(KEYINPUT34), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  NAND2_X1  g476(.A1(new_n428), .A2(new_n432), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n663), .A2(new_n376), .A3(new_n384), .A4(new_n440), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n643), .B(new_n664), .C1(new_n512), .C2(new_n516), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n642), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  INV_X1    g483(.A(new_n567), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n552), .A2(new_n522), .A3(KEYINPUT25), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT72), .B1(new_n561), .B2(new_n562), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n560), .A2(new_n565), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n544), .A2(new_n548), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n526), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n678), .A2(new_n569), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n669), .B1(new_n675), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n679), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n568), .A2(KEYINPUT102), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n640), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n447), .A2(new_n521), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  NAND2_X1  g500(.A1(new_n624), .A2(new_n630), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n643), .B1(new_n512), .B2(new_n516), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT102), .B1(new_n568), .B2(new_n681), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n669), .B(new_n679), .C1(new_n566), .C2(new_n567), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n687), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n635), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n652), .A2(new_n656), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT103), .B(G900), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n694), .A2(new_n438), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n435), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n693), .A2(new_n663), .A3(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n691), .A2(new_n692), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n217), .ZN(G30));
  NAND2_X1  g513(.A1(new_n517), .A2(new_n520), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT38), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n596), .B1(new_n600), .B2(new_n588), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n188), .B1(new_n589), .B2(new_n594), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT104), .Z(new_n705));
  NAND3_X1  g519(.A1(new_n630), .A2(new_n622), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n689), .A2(new_n690), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n518), .A3(new_n385), .A4(new_n663), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n701), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n696), .B(KEYINPUT39), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n635), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT40), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT106), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT40), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n713), .B(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n711), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  AOI22_X1  g535(.A1(new_n680), .A2(new_n682), .B1(new_n630), .B2(new_n624), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n385), .A2(new_n649), .A3(new_n696), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(new_n635), .A3(new_n688), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  INV_X1    g540(.A(new_n307), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT81), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n269), .A2(new_n270), .A3(new_n279), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n296), .B1(new_n729), .B2(new_n189), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n282), .B1(new_n730), .B2(new_n280), .ZN(new_n731));
  INV_X1    g545(.A(new_n288), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n304), .A3(new_n289), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n187), .B1(new_n734), .B2(new_n188), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n727), .A2(new_n735), .A3(new_n634), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n658), .A3(new_n631), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT41), .B(G113), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G15));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n631), .A3(new_n665), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  NAND4_X1  g555(.A1(new_n722), .A2(new_n445), .A3(new_n736), .A4(new_n688), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NAND3_X1  g557(.A1(new_n639), .A2(KEYINPUT107), .A3(new_n625), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(G472), .C1(new_n637), .C2(new_n638), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n747), .A2(new_n636), .A3(new_n440), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n385), .A2(new_n663), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n643), .B(new_n749), .C1(new_n516), .C2(new_n512), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n736), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  OAI21_X1  g566(.A(new_n747), .B1(new_n689), .B2(new_n690), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g569(.A(KEYINPUT108), .B(new_n747), .C1(new_n689), .C2(new_n690), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n734), .A2(new_n188), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(G469), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n688), .A2(new_n759), .A3(new_n446), .A4(new_n307), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(new_n724), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  AOI21_X1  g577(.A(new_n643), .B1(new_n517), .B2(new_n520), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n631), .A3(new_n635), .A4(new_n724), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n700), .A2(new_n518), .A3(new_n635), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n604), .A2(new_n612), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n622), .B1(new_n768), .B2(new_n572), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n625), .A2(new_n628), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n636), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n724), .A2(KEYINPUT42), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n264), .ZN(G33));
  INV_X1    g589(.A(new_n697), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n767), .A2(new_n631), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NAND2_X1  g592(.A1(new_n693), .A2(new_n649), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT43), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n780), .A2(new_n709), .A3(new_n641), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n764), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n309), .A2(KEYINPUT45), .ZN(new_n787));
  OAI21_X1  g601(.A(G469), .B1(new_n309), .B2(KEYINPUT45), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(G469), .A2(G902), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n727), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n790), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n634), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n712), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(KEYINPUT110), .A3(new_n712), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n786), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n795), .A2(new_n807), .A3(new_n803), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n795), .B2(new_n803), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n764), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n811), .A2(new_n687), .A3(new_n636), .A4(new_n723), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n806), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  NAND2_X1  g628(.A1(new_n764), .A2(new_n736), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n815), .A2(new_n435), .A3(new_n780), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n769), .A2(new_n770), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n636), .A3(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT48), .Z(new_n819));
  XNOR2_X1  g633(.A(new_n706), .B(KEYINPUT105), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n820), .A2(new_n815), .A3(new_n571), .A4(new_n435), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n385), .A3(new_n649), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n747), .A2(new_n636), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n780), .A2(new_n823), .A3(new_n435), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n761), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n822), .A2(G952), .A3(new_n286), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n385), .A2(new_n649), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n821), .A2(new_n827), .B1(new_n757), .B2(new_n816), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n701), .A2(new_n643), .A3(new_n736), .A4(new_n824), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT50), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT50), .B1(new_n829), .B2(new_n830), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n727), .A2(new_n735), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n806), .A2(new_n810), .B1(new_n634), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n824), .A2(new_n764), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT117), .Z(new_n838));
  OAI21_X1  g652(.A(new_n834), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n819), .B(new_n826), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n723), .B1(new_n755), .B2(new_n756), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n663), .B(new_n385), .C1(new_n435), .C2(new_n695), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n722), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n767), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n765), .A2(new_n766), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n767), .A2(new_n773), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n848), .A2(new_n851), .A3(new_n777), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n736), .B(new_n631), .C1(new_n658), .C2(new_n665), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n742), .A2(new_n853), .A3(new_n751), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT113), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n742), .A2(new_n853), .A3(new_n751), .A4(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n447), .B(new_n521), .C1(new_n683), .C2(new_n631), .ZN(new_n859));
  INV_X1    g673(.A(new_n664), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n642), .A2(new_n521), .A3(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n657), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n517), .A2(new_n520), .A3(new_n518), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n642), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n852), .A2(new_n858), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n698), .B1(new_n761), .B2(new_n844), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n696), .B(KEYINPUT115), .Z(new_n874));
  NOR3_X1   g688(.A1(new_n675), .A2(new_n679), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n750), .A2(new_n635), .A3(new_n706), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n680), .A2(new_n682), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n687), .A3(new_n635), .A4(new_n688), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n878), .B2(new_n723), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT52), .B1(new_n873), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n723), .B(new_n760), .C1(new_n755), .C2(new_n756), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n882), .A2(new_n879), .A3(new_n698), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n872), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n855), .A2(new_n869), .A3(new_n862), .A4(new_n857), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n848), .A2(new_n851), .A3(new_n777), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n878), .A2(new_n697), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n762), .A2(new_n891), .A3(new_n725), .A4(new_n876), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n883), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n873), .A2(KEYINPUT52), .A3(new_n880), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT54), .B1(new_n887), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n886), .B1(new_n872), .B2(new_n885), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n742), .A2(new_n853), .A3(new_n751), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT116), .B1(new_n900), .B2(new_n851), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n774), .A2(new_n854), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n777), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n870), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n895), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n898), .A2(new_n899), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n843), .A2(new_n909), .B1(G952), .B2(G953), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n835), .B(KEYINPUT49), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n571), .A2(new_n779), .A3(new_n643), .A4(new_n634), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n701), .A2(new_n911), .A3(new_n708), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n910), .A2(new_n913), .ZN(G75));
  AND3_X1   g728(.A1(new_n895), .A2(new_n904), .A3(new_n906), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n896), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n188), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(G210), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n500), .A2(new_n502), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n504), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n918), .B2(new_n919), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n286), .A2(G952), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G51));
  NOR3_X1   g740(.A1(new_n916), .A2(new_n188), .A3(new_n789), .ZN(new_n927));
  INV_X1    g741(.A(new_n734), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT54), .B1(new_n915), .B2(new_n896), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n908), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n790), .B(KEYINPUT57), .Z(new_n931));
  AOI21_X1  g745(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n931), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n929), .B2(new_n908), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT119), .B1(new_n936), .B2(new_n928), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n925), .B1(new_n934), .B2(new_n937), .ZN(G54));
  INV_X1    g752(.A(KEYINPUT120), .ZN(new_n939));
  AND2_X1   g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n917), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n941), .B2(new_n366), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n925), .B1(new_n941), .B2(new_n366), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n917), .A2(KEYINPUT120), .A3(new_n372), .A4(new_n940), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(G60));
  OR2_X1    g759(.A1(new_n645), .A2(new_n646), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT59), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n909), .B2(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n930), .A2(new_n946), .A3(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n925), .ZN(G63));
  INV_X1    g765(.A(new_n925), .ZN(new_n952));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n898), .B2(new_n907), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n564), .B(KEYINPUT122), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT121), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n958), .A3(new_n678), .ZN(new_n959));
  INV_X1    g773(.A(new_n954), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n678), .B(new_n960), .C1(new_n915), .C2(new_n896), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT121), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n957), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n955), .B2(new_n956), .ZN(new_n965));
  INV_X1    g779(.A(new_n956), .ZN(new_n966));
  OAI211_X1 g780(.A(KEYINPUT123), .B(new_n966), .C1(new_n916), .C2(new_n954), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n965), .A2(new_n967), .A3(KEYINPUT61), .A4(new_n952), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n959), .A2(new_n962), .ZN(new_n969));
  OAI22_X1  g783(.A1(new_n963), .A2(KEYINPUT61), .B1(new_n968), .B2(new_n969), .ZN(G66));
  AOI21_X1  g784(.A(new_n286), .B1(new_n437), .B2(G224), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT124), .ZN(new_n972));
  INV_X1    g786(.A(new_n888), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(G953), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n920), .B1(G898), .B2(new_n286), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G69));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n785), .B1(new_n798), .B2(new_n799), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n873), .A2(new_n725), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n979), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n801), .A2(KEYINPUT127), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n800), .A2(new_n636), .A3(new_n750), .A4(new_n817), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n851), .A2(new_n777), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n813), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n986), .A3(new_n286), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n598), .A2(new_n599), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(new_n345), .Z(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(G900), .B2(G953), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n989), .B(KEYINPUT125), .ZN(new_n992));
  INV_X1    g806(.A(new_n631), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n385), .A2(new_n649), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n693), .B2(new_n663), .ZN(new_n995));
  NOR4_X1   g809(.A1(new_n811), .A2(new_n993), .A3(new_n713), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n786), .B2(new_n800), .ZN(new_n997));
  INV_X1    g811(.A(new_n720), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT62), .B1(new_n998), .B2(new_n979), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n981), .A2(new_n720), .A3(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n813), .A2(new_n997), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n992), .B1(new_n1002), .B2(new_n286), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1003), .A2(KEYINPUT126), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1005));
  AOI211_X1 g819(.A(new_n1005), .B(new_n992), .C1(new_n1002), .C2(new_n286), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n991), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n286), .B1(G227), .B2(G900), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1008), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n1010), .B(new_n991), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(G72));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  OAI21_X1  g828(.A(new_n1014), .B1(new_n1002), .B2(new_n888), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n702), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n603), .A2(new_n619), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1014), .B(new_n1017), .C1(new_n887), .C2(new_n896), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1016), .A2(new_n952), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n983), .A2(new_n986), .A3(new_n973), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n1014), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n601), .A2(new_n594), .A3(new_n602), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(G57));
endmodule


