//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(G131), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT80), .A2(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT80), .A2(G143), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(G237), .A2(G953), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n194), .B(G214), .C1(KEYINPUT80), .C2(G143), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n187), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT17), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT83), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(KEYINPUT83), .A3(KEYINPUT17), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT16), .B1(new_n202), .B2(G125), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT70), .B1(KEYINPUT69), .B2(G125), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT70), .A2(G125), .ZN(new_n205));
  OAI21_X1  g019(.A(G140), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT69), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT70), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n202), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n203), .B1(new_n211), .B2(KEYINPUT16), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n211), .A2(KEYINPUT16), .ZN(new_n215));
  OAI21_X1  g029(.A(G146), .B1(new_n215), .B2(new_n203), .ZN(new_n216));
  INV_X1    g030(.A(new_n196), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n193), .A2(new_n187), .A3(new_n195), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n201), .A2(new_n214), .A3(new_n216), .A4(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G113), .B(G122), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n193), .A2(new_n195), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT18), .A2(G131), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n206), .A2(new_n228), .A3(new_n210), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n206), .B2(new_n210), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n213), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n202), .A2(G125), .ZN(new_n234));
  INV_X1    g048(.A(G125), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G140), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n236), .A3(new_n213), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n227), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n221), .A2(new_n224), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT19), .B1(new_n229), .B2(new_n231), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT19), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n234), .A2(new_n236), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n213), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT82), .A3(new_n216), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n217), .A2(new_n219), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT82), .B1(new_n244), .B2(new_n216), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n239), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n224), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n240), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G475), .A2(G902), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT20), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT20), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n244), .A2(new_n216), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n245), .A3(new_n246), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n224), .B1(new_n259), .B2(new_n239), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n255), .B(new_n252), .C1(new_n260), .C2(new_n240), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G475), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n224), .B1(new_n221), .B2(new_n239), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT84), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n221), .A2(new_n224), .A3(new_n239), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G902), .B1(new_n264), .B2(KEYINPUT84), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n263), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT9), .B(G234), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(G217), .A3(new_n189), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G116), .B(G122), .ZN(new_n276));
  INV_X1    g090(.A(G107), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT64), .B(G134), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G128), .ZN(new_n281));
  INV_X1    g095(.A(G128), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G143), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT13), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n283), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n281), .A2(new_n285), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT85), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n281), .A2(new_n289), .A3(new_n285), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G134), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n278), .B(new_n284), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G116), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT14), .A3(G122), .ZN(new_n295));
  INV_X1    g109(.A(new_n276), .ZN(new_n296));
  OAI211_X1 g110(.A(G107), .B(new_n295), .C1(new_n296), .C2(KEYINPUT14), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n276), .A2(new_n277), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n299));
  INV_X1    g113(.A(new_n284), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(new_n298), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n275), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n293), .A2(new_n301), .A3(new_n275), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G478), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(KEYINPUT15), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n304), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n302), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n307), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(G234), .A2(G237), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(G952), .A3(new_n189), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT21), .B(G898), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(G902), .A3(G953), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT86), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n262), .A2(new_n271), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT87), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n270), .B1(new_n254), .B2(new_n261), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT87), .A3(new_n324), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n194), .A2(G210), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT27), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G101), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT2), .B(G113), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G116), .B(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(G116), .B(G119), .Z(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n336), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT11), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n279), .B2(G137), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n292), .A2(G137), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n279), .B2(G137), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n187), .B(new_n345), .C1(new_n347), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n292), .A2(KEYINPUT64), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT64), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G134), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G137), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n292), .A2(G137), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G131), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n213), .A2(G143), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n280), .A2(G146), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n361), .A2(KEYINPUT1), .A3(new_n282), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT65), .ZN(new_n363));
  AOI21_X1  g177(.A(G128), .B1(new_n359), .B2(new_n360), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n365), .A2(new_n213), .A3(G143), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n363), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n213), .A2(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT1), .ZN(new_n369));
  XNOR2_X1  g183(.A(G143), .B(G146), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n369), .B(KEYINPUT65), .C1(new_n370), .C2(G128), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n362), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n358), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT0), .B(G128), .Z(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(new_n370), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT0), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(new_n282), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n361), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n349), .A2(new_n351), .A3(G137), .ZN(new_n380));
  INV_X1    g194(.A(new_n346), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n344), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT11), .B1(new_n352), .B2(new_n353), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n379), .B1(new_n384), .B2(new_n348), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT30), .B1(new_n373), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n348), .ZN(new_n387));
  INV_X1    g201(.A(new_n379), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n370), .A2(new_n365), .A3(G128), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n280), .A2(G146), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n282), .B1(new_n391), .B2(new_n368), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT65), .B1(new_n392), .B2(new_n369), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n364), .A2(new_n363), .A3(new_n366), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n348), .A3(new_n357), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n389), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n343), .B1(new_n386), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT66), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n342), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n389), .A2(new_n401), .A3(new_n396), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n335), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n389), .A2(new_n396), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n342), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT28), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n187), .B1(new_n354), .B2(new_n355), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n382), .A2(new_n383), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(new_n187), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n395), .A2(new_n411), .B1(new_n387), .B2(new_n388), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n412), .B2(new_n401), .ZN(new_n413));
  AND4_X1   g227(.A1(new_n408), .A2(new_n389), .A3(new_n401), .A4(new_n396), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n407), .B(new_n334), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n404), .A2(new_n405), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT67), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n404), .A2(KEYINPUT67), .A3(new_n415), .A4(new_n405), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n402), .A2(KEYINPUT28), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n412), .A2(new_n408), .A3(new_n401), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n401), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n406), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n335), .A2(new_n405), .ZN(new_n426));
  AOI21_X1  g240(.A(G902), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G472), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n334), .B1(new_n422), .B2(new_n407), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n373), .A2(KEYINPUT30), .A3(new_n385), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n397), .B1(new_n389), .B2(new_n396), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n342), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n402), .A3(new_n334), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT31), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n386), .A2(new_n398), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n403), .B1(new_n437), .B2(new_n342), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT31), .A3(new_n334), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n430), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G472), .A2(G902), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n440), .A2(KEYINPUT32), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT32), .ZN(new_n444));
  INV_X1    g258(.A(new_n430), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT31), .B1(new_n438), .B2(new_n334), .ZN(new_n446));
  NOR4_X1   g260(.A1(new_n399), .A2(new_n403), .A3(new_n435), .A4(new_n335), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n444), .B1(new_n448), .B2(new_n441), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n429), .B1(new_n443), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G234), .ZN(new_n451));
  OAI21_X1  g265(.A(G217), .B1(new_n451), .B2(G902), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n452), .B(KEYINPUT68), .Z(new_n453));
  NAND2_X1  g267(.A1(new_n216), .A2(new_n214), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT23), .ZN(new_n455));
  INV_X1    g269(.A(G119), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n456), .B2(G128), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n282), .A2(KEYINPUT23), .A3(G119), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n457), .B(new_n458), .C1(G119), .C2(new_n282), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G110), .ZN(new_n460));
  XOR2_X1   g274(.A(KEYINPUT24), .B(G110), .Z(new_n461));
  XNOR2_X1  g275(.A(G119), .B(G128), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n212), .A2(new_n213), .ZN(new_n467));
  OAI22_X1  g281(.A1(new_n459), .A2(G110), .B1(new_n462), .B2(new_n461), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n237), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT22), .B(G137), .ZN(new_n472));
  INV_X1    g286(.A(G221), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(new_n451), .A3(G953), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n472), .B(new_n474), .Z(new_n475));
  NAND3_X1  g289(.A1(new_n466), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n475), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n464), .B1(new_n216), .B2(new_n214), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(new_n470), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n310), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT25), .A4(new_n310), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n453), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n476), .A2(new_n479), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n452), .A2(new_n310), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  INV_X1    g303(.A(G101), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n491));
  AOI22_X1  g305(.A1(KEYINPUT73), .A2(new_n491), .B1(new_n223), .B2(G107), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n493));
  AND4_X1   g307(.A1(new_n493), .A2(new_n277), .A3(KEYINPUT3), .A4(G104), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n493), .A2(KEYINPUT3), .B1(new_n277), .B2(G104), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n490), .B(new_n492), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n223), .A2(G107), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n277), .A2(G104), .ZN(new_n498));
  OAI21_X1  g312(.A(G101), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n496), .A2(KEYINPUT10), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT74), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n395), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n496), .A2(KEYINPUT10), .A3(new_n499), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT74), .B1(new_n372), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n387), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G101), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(KEYINPUT4), .A3(new_n496), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n510), .A3(G101), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n388), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n390), .A2(new_n392), .A3(new_n369), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n499), .A3(new_n496), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT10), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n505), .A2(new_n506), .A3(new_n512), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n189), .A2(G227), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT71), .ZN(new_n519));
  XNOR2_X1  g333(.A(G110), .B(G140), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n496), .A2(new_n499), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n514), .B1(new_n395), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT12), .A3(new_n387), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT12), .B1(new_n525), .B2(new_n387), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT12), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n372), .A2(new_n523), .ZN(new_n531));
  AOI221_X4 g345(.A(new_n530), .B1(new_n348), .B2(new_n384), .C1(new_n531), .C2(new_n514), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n529), .B1(new_n532), .B2(KEYINPUT75), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n522), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n501), .B1(new_n395), .B2(new_n500), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n372), .A2(new_n503), .A3(KEYINPUT74), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n512), .A2(new_n516), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n387), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n521), .B1(new_n539), .B2(new_n517), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n489), .B(new_n310), .C1(new_n534), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(G469), .A2(G902), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n517), .A2(new_n521), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n539), .ZN(new_n544));
  INV_X1    g358(.A(new_n517), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n533), .B2(new_n528), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n521), .B(KEYINPUT72), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n544), .B(G469), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n541), .A2(new_n542), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n473), .B1(new_n273), .B2(new_n310), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G214), .B1(G237), .B2(G902), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G210), .B1(G237), .B2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n509), .A2(new_n342), .A3(new_n511), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n338), .A2(KEYINPUT5), .ZN(new_n558));
  OR3_X1    g372(.A1(new_n294), .A2(KEYINPUT5), .A3(G119), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(G113), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT76), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n560), .A2(new_n561), .B1(new_n338), .B2(new_n337), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n558), .A2(KEYINPUT76), .A3(G113), .A4(new_n559), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n524), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G122), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n557), .A2(new_n564), .A3(new_n566), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(KEYINPUT6), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n370), .B1(new_n376), .B2(new_n282), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n571), .B(G125), .C1(new_n370), .C2(new_n374), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT77), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n372), .A2(new_n235), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT77), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G224), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G953), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n580), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n574), .A2(new_n575), .A3(new_n582), .A4(new_n577), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT6), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n565), .A2(new_n585), .A3(new_n567), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n570), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n562), .A2(new_n523), .A3(new_n563), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n560), .A2(new_n339), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n524), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT78), .B(KEYINPUT8), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n566), .B(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n582), .A2(KEYINPUT7), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n574), .A2(new_n575), .A3(new_n577), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n569), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n573), .B1(new_n575), .B2(KEYINPUT79), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT79), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n372), .A2(new_n599), .A3(new_n235), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n595), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n310), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n556), .B1(new_n587), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n569), .A2(new_n596), .A3(new_n593), .ZN(new_n604));
  INV_X1    g418(.A(new_n601), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n570), .A2(new_n584), .A3(new_n586), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(new_n555), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n554), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n552), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n330), .A2(new_n450), .A3(new_n488), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  INV_X1    g427(.A(KEYINPUT88), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n603), .A2(new_n614), .A3(new_n608), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n555), .B1(new_n606), .B2(new_n607), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n554), .B1(new_n616), .B2(KEYINPUT88), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n617), .A3(new_n322), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n303), .A2(KEYINPUT90), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n303), .A2(KEYINPUT90), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(KEYINPUT33), .A3(new_n304), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n311), .B2(new_n302), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n306), .A2(G902), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n624), .A2(new_n625), .B1(new_n306), .B2(new_n312), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n618), .A2(new_n328), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G472), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n448), .B2(new_n310), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n440), .A2(new_n442), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n488), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n552), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n627), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND3_X1  g450(.A1(new_n254), .A2(new_n261), .A3(KEYINPUT91), .ZN(new_n637));
  INV_X1    g451(.A(new_n251), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT91), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n255), .A4(new_n252), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n270), .A2(new_n314), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n618), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n633), .A3(new_n631), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT92), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT35), .B(G107), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NAND2_X1  g461(.A1(new_n466), .A2(new_n471), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n477), .A2(KEYINPUT36), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n486), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n484), .A2(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n629), .A2(new_n630), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n330), .A2(new_n611), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT93), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT37), .B(G110), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  NAND4_X1  g473(.A1(new_n549), .A2(new_n551), .A3(new_n615), .A4(new_n617), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n320), .A2(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n317), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n642), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n654), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n450), .A2(new_n661), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  NAND2_X1  g482(.A1(new_n262), .A2(new_n271), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n315), .A3(new_n553), .A4(new_n654), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT94), .Z(new_n671));
  AND3_X1   g485(.A1(new_n606), .A2(new_n607), .A3(new_n555), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n616), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT38), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT32), .B1(new_n440), .B2(new_n442), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n448), .A2(new_n444), .A3(new_n441), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n402), .A2(new_n335), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(G902), .B1(new_n680), .B2(new_n424), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n438), .A2(new_n335), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n675), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n671), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n663), .B(KEYINPUT39), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n549), .A2(new_n551), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT40), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT95), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT96), .ZN(new_n692));
  OR3_X1    g506(.A1(new_n687), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n692), .B1(new_n687), .B2(new_n691), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n280), .ZN(G45));
  NOR3_X1   g510(.A1(new_n328), .A2(new_n626), .A3(new_n664), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n450), .A2(new_n661), .A3(new_n666), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NAND4_X1  g513(.A1(new_n525), .A2(KEYINPUT75), .A3(KEYINPUT12), .A4(new_n387), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n506), .B1(new_n514), .B2(new_n531), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n528), .B(new_n700), .C1(KEYINPUT12), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n539), .A2(new_n517), .ZN(new_n703));
  INV_X1    g517(.A(new_n521), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n702), .A2(new_n543), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(G469), .B1(new_n705), .B2(G902), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n551), .A3(new_n541), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n627), .A2(new_n450), .A3(new_n488), .A4(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT41), .B(G113), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT97), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n709), .B(new_n711), .ZN(G15));
  NAND4_X1  g526(.A1(new_n643), .A2(new_n450), .A3(new_n488), .A4(new_n708), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT98), .B(G116), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G18));
  NAND2_X1  g529(.A1(new_n615), .A2(new_n617), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n707), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n330), .A2(new_n450), .A3(new_n666), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  XOR2_X1   g533(.A(KEYINPUT100), .B(G472), .Z(new_n720));
  OAI21_X1  g534(.A(new_n720), .B1(new_n440), .B2(G902), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT99), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n334), .B1(new_n422), .B2(new_n424), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n436), .B2(new_n439), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n722), .B1(new_n724), .B2(new_n442), .ZN(new_n725));
  OAI22_X1  g539(.A1(new_n446), .A2(new_n447), .B1(new_n334), .B2(new_n425), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(KEYINPUT99), .A3(new_n441), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n721), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n716), .A2(new_n328), .A3(new_n314), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n707), .A2(new_n323), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n729), .A3(new_n488), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND4_X1  g546(.A1(new_n728), .A2(new_n666), .A3(new_n697), .A4(new_n717), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  XNOR2_X1  g548(.A(new_n542), .B(KEYINPUT101), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n541), .A2(new_n548), .A3(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n672), .A2(new_n616), .A3(new_n554), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n736), .A2(new_n737), .A3(new_n551), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n450), .A2(new_n488), .A3(new_n697), .A4(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n676), .A2(new_n677), .B1(new_n428), .B2(G472), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n632), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(KEYINPUT42), .A3(new_n697), .A4(new_n738), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  AND4_X1   g560(.A1(new_n450), .A2(new_n665), .A3(new_n488), .A4(new_n738), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n292), .ZN(G36));
  AND2_X1   g562(.A1(new_n688), .A2(new_n551), .ZN(new_n749));
  INV_X1    g563(.A(new_n735), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n547), .B1(new_n702), .B2(new_n517), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n539), .A2(new_n517), .A3(new_n521), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n544), .B(KEYINPUT45), .C1(new_n546), .C2(new_n547), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT102), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n489), .B1(new_n759), .B2(new_n751), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(KEYINPUT102), .A3(new_n755), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n750), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n541), .B1(new_n762), .B2(KEYINPUT46), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n764), .B(new_n750), .C1(new_n758), .C2(new_n761), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n749), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT103), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT103), .B(new_n749), .C1(new_n763), .C2(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n669), .A2(new_n626), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n631), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n666), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n771), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n772), .B(KEYINPUT43), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n775), .A4(new_n666), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n777), .A2(new_n779), .A3(new_n737), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n770), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  OAI21_X1  g596(.A(new_n551), .B1(new_n763), .B2(new_n765), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n785), .B(new_n551), .C1(new_n763), .C2(new_n765), .ZN(new_n786));
  INV_X1    g600(.A(new_n626), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n669), .A2(new_n787), .A3(new_n663), .ZN(new_n788));
  INV_X1    g602(.A(new_n737), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n450), .A2(new_n788), .A3(new_n488), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n784), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NOR4_X1   g606(.A1(new_n675), .A2(new_n632), .A3(new_n554), .A4(new_n550), .ZN(new_n793));
  INV_X1    g607(.A(new_n685), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n706), .A2(new_n541), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT49), .Z(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n772), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n728), .A2(new_n488), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n674), .A2(new_n554), .A3(new_n708), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT107), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n774), .B2(new_n317), .ZN(new_n801));
  INV_X1    g615(.A(new_n317), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n778), .A2(KEYINPUT107), .A3(new_n802), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n798), .B(new_n799), .C1(new_n801), .C2(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(KEYINPUT109), .A2(KEYINPUT50), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n807));
  OAI21_X1  g621(.A(new_n806), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n784), .A2(new_n786), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n795), .A2(new_n551), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n801), .A2(new_n803), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n488), .A3(new_n728), .A4(new_n737), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n808), .B(KEYINPUT51), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n789), .A2(new_n707), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n794), .A2(new_n488), .A3(new_n802), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n328), .A3(new_n626), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT112), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n812), .A2(KEYINPUT110), .A3(new_n815), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT110), .B1(new_n812), .B2(new_n815), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n666), .B(new_n728), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n814), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n818), .A2(new_n819), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n669), .A2(new_n787), .ZN(new_n828));
  OAI211_X1 g642(.A(G952), .B(new_n189), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n812), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n798), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(new_n831), .B2(new_n717), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT48), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n822), .A2(new_n823), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(new_n743), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n833), .B(new_n743), .C1(new_n822), .C2(new_n823), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n832), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n826), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT108), .B1(new_n811), .B2(new_n813), .ZN(new_n841));
  INV_X1    g655(.A(new_n813), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT108), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n842), .B(new_n843), .C1(new_n809), .C2(new_n810), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n821), .A2(new_n808), .A3(new_n824), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(KEYINPUT113), .B(new_n840), .C1(new_n845), .C2(new_n846), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n839), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n667), .A2(new_n733), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n742), .A2(new_n654), .A3(new_n660), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n484), .A2(new_n653), .A3(new_n664), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n736), .A2(new_n854), .A3(new_n551), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n678), .B2(new_n684), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n853), .A2(new_n697), .B1(new_n729), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n852), .A2(new_n857), .A3(KEYINPUT105), .ZN(new_n858));
  INV_X1    g672(.A(new_n855), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n685), .A2(new_n729), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n667), .A2(new_n698), .A3(new_n733), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT105), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT52), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n747), .B1(new_n741), .B2(new_n744), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n612), .A2(new_n709), .A3(new_n713), .A4(new_n656), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n309), .A2(KEYINPUT104), .A3(new_n313), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT104), .B1(new_n309), .B2(new_n313), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n328), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n828), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n610), .A2(new_n323), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n633), .A3(new_n631), .A4(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n718), .A2(new_n731), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n721), .A2(new_n725), .A3(new_n727), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n875), .A2(new_n788), .A3(new_n654), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n742), .A2(new_n654), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n869), .A2(new_n664), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n737), .A2(new_n878), .A3(new_n271), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n637), .A2(new_n640), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n552), .A3(new_n880), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n876), .A2(new_n738), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n865), .A2(new_n866), .A3(new_n874), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n864), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n858), .A2(new_n863), .A3(KEYINPUT52), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n861), .A2(KEYINPUT52), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n864), .A2(new_n883), .A3(new_n887), .A4(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n886), .A2(new_n890), .A3(KEYINPUT54), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT105), .B1(new_n852), .B2(new_n857), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n861), .A2(new_n862), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n866), .A2(new_n874), .ZN(new_n897));
  INV_X1    g711(.A(new_n747), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n736), .A2(new_n737), .A3(new_n551), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n742), .A2(new_n632), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT42), .B1(new_n900), .B2(new_n697), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n739), .A2(new_n740), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n898), .B(new_n882), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n896), .A2(new_n904), .A3(new_n888), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n887), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n896), .A2(new_n904), .A3(KEYINPUT53), .A4(new_n885), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n892), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT106), .B1(new_n891), .B2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n864), .A2(new_n883), .A3(new_n889), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n907), .B1(new_n910), .B2(KEYINPUT53), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n884), .A2(KEYINPUT53), .A3(new_n888), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n896), .A2(new_n904), .A3(new_n885), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n913), .B(new_n892), .C1(new_n914), .C2(KEYINPUT53), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT106), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n851), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(G952), .A2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n797), .B1(new_n918), .B2(new_n919), .ZN(G75));
  OAI21_X1  g734(.A(new_n913), .B1(new_n914), .B2(KEYINPUT53), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(G210), .A3(G902), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n570), .A2(new_n586), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n584), .ZN(new_n925));
  XNOR2_X1  g739(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n925), .B(new_n926), .Z(new_n927));
  AND3_X1   g741(.A1(new_n922), .A2(new_n923), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n922), .B2(new_n923), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n189), .A2(G952), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(G51));
  NAND4_X1  g745(.A1(new_n921), .A2(G902), .A3(new_n758), .A4(new_n761), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT117), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n705), .B(KEYINPUT115), .Z(new_n935));
  NAND2_X1  g749(.A1(new_n921), .A2(KEYINPUT54), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n915), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n735), .B(KEYINPUT57), .Z(new_n938));
  AOI21_X1  g752(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT116), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n930), .B1(new_n941), .B2(new_n942), .ZN(G54));
  AND4_X1   g757(.A1(KEYINPUT58), .A2(new_n921), .A3(G475), .A4(G902), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(new_n638), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n638), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(new_n930), .ZN(G60));
  XNOR2_X1  g761(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n306), .A2(new_n310), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n909), .A2(new_n917), .A3(new_n951), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n624), .B(KEYINPUT118), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n950), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n930), .B1(new_n937), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(KEYINPUT120), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT120), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n954), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(G63));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT121), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n921), .A2(new_n650), .A3(new_n652), .A4(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n921), .A2(new_n965), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n930), .B1(new_n971), .B2(new_n485), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n968), .B2(new_n969), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI221_X1 g789(.A(new_n972), .B1(new_n962), .B2(KEYINPUT61), .C1(new_n968), .C2(new_n969), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G66));
  OAI21_X1  g791(.A(G953), .B1(new_n318), .B2(new_n579), .ZN(new_n978));
  INV_X1    g792(.A(new_n897), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(G953), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n924), .B1(G898), .B2(new_n189), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G69));
  AOI21_X1  g796(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n743), .A2(new_n729), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n770), .A2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n667), .A2(new_n698), .A3(new_n733), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n865), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n781), .A2(new_n988), .A3(new_n791), .A4(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g808(.A1(new_n809), .A2(new_n790), .B1(new_n770), .B2(new_n987), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n990), .B1(new_n770), .B2(new_n780), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT124), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n189), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n189), .A2(G900), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n998), .A2(KEYINPUT125), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n992), .A2(new_n993), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n995), .A2(KEYINPUT124), .A3(new_n996), .ZN(new_n1004));
  AOI21_X1  g818(.A(G953), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1002), .B1(new_n1005), .B2(new_n999), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n241), .A2(new_n243), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n437), .B(new_n1007), .Z(new_n1008));
  NAND3_X1  g822(.A1(new_n1001), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n693), .A2(new_n694), .A3(new_n989), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  INV_X1    g825(.A(new_n743), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1012), .A2(new_n689), .A3(new_n789), .ZN(new_n1013));
  AOI22_X1  g827(.A1(new_n770), .A2(new_n780), .B1(new_n871), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n693), .A2(new_n694), .A3(new_n1015), .A4(new_n989), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1011), .A2(new_n791), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n189), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1008), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n984), .B(new_n985), .C1(new_n1009), .C2(new_n1020), .ZN(new_n1021));
  AND4_X1   g835(.A1(KEYINPUT126), .A2(new_n1009), .A3(new_n983), .A4(new_n1020), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1021), .A2(new_n1022), .ZN(G72));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  NAND2_X1  g839(.A1(new_n404), .A2(new_n434), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n911), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1027), .B1(G952), .B2(new_n189), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1003), .A2(new_n1004), .A3(new_n979), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1025), .B(KEYINPUT127), .Z(new_n1030));
  AOI211_X1 g844(.A(new_n399), .B(new_n679), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1030), .B1(new_n1017), .B2(new_n897), .ZN(new_n1032));
  AOI211_X1 g846(.A(new_n1028), .B(new_n1031), .C1(new_n683), .C2(new_n1032), .ZN(G57));
endmodule


