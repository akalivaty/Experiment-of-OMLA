//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0004(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G116), .ZN(new_n206));
  INV_X1    g0006(.A(G270), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n208), .B(new_n214), .C1(G97), .C2(G257), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G1), .B2(G20), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT1), .Z(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G1), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n222), .A2(new_n219), .A3(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NOR3_X1   g0025(.A1(new_n217), .A2(new_n221), .A3(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND3_X1  g0041(.A1(new_n222), .A2(G13), .A3(G20), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  AND2_X1   g0044(.A1(new_n244), .A2(new_n220), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n245), .B1(G1), .B2(new_n219), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(new_n210), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n219), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n248), .A2(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n255), .B1(new_n252), .B2(new_n250), .C1(new_n248), .C2(new_n249), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n254), .B(new_n256), .C1(new_n219), .C2(new_n201), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n244), .A2(new_n220), .ZN(new_n258));
  AOI211_X1 g0058(.A(new_n243), .B(new_n247), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G179), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT64), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT64), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G33), .A3(G41), .ZN(new_n264));
  INV_X1    g0064(.A(new_n220), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n222), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G226), .A3(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n222), .B(G274), .C1(G41), .C2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n270), .A2(KEYINPUT65), .ZN(new_n271));
  OR2_X1    g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT66), .B(G223), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n274), .B(new_n276), .C1(new_n277), .C2(new_n275), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n265), .A2(new_n261), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n278), .B(new_n280), .C1(G77), .C2(new_n274), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n270), .A2(KEYINPUT65), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n271), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n259), .B1(new_n260), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(G169), .B2(new_n284), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  OR3_X1    g0088(.A1(new_n259), .A2(new_n288), .A3(KEYINPUT9), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n288), .B1(new_n259), .B2(KEYINPUT9), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(G200), .ZN(new_n292));
  AOI22_X1  g0092(.A1(G190), .A2(new_n284), .B1(new_n259), .B2(KEYINPUT9), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT10), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n291), .A2(new_n296), .A3(new_n292), .A4(new_n293), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n287), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(G58), .A2(G68), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G58), .A2(G68), .ZN(new_n300));
  OAI21_X1  g0100(.A(G20), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT75), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n251), .A2(G159), .ZN(new_n304));
  OAI211_X1 g0104(.A(KEYINPUT75), .B(G20), .C1(new_n299), .C2(new_n300), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n219), .A4(new_n273), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT74), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(KEYINPUT3), .A2(G33), .ZN(new_n310));
  NOR2_X1   g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT7), .B1(new_n312), .B2(new_n219), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n272), .A2(new_n219), .A3(new_n273), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(KEYINPUT74), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G68), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n306), .B(KEYINPUT16), .C1(new_n314), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n310), .A2(new_n311), .A3(G20), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT76), .B1(new_n321), .B2(KEYINPUT7), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT76), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n315), .A2(new_n323), .A3(new_n316), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n307), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n320), .B1(new_n325), .B2(G68), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n258), .B(new_n319), .C1(new_n326), .C2(KEYINPUT16), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n266), .A2(G232), .A3(new_n267), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n269), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n211), .A2(G1698), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n331), .B1(G223), .B2(G1698), .C1(new_n310), .C2(new_n311), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G87), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n279), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n328), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(KEYINPUT77), .ZN(new_n336));
  INV_X1    g0136(.A(new_n334), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT77), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n329), .A2(new_n338), .A3(new_n269), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n335), .B1(new_n340), .B2(G190), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n248), .A2(new_n242), .ZN(new_n342));
  INV_X1    g0142(.A(new_n246), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(new_n248), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n327), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT17), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n327), .A2(new_n341), .A3(KEYINPUT17), .A4(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n336), .A2(new_n337), .A3(new_n260), .A4(new_n339), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n330), .B2(new_n334), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AOI211_X1 g0155(.A(new_n351), .B(new_n355), .C1(new_n344), .C2(new_n327), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n319), .A2(new_n258), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n344), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n355), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT18), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT15), .B(G87), .Z(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n249), .A2(new_n364), .B1(new_n248), .B2(new_n252), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n219), .A2(new_n202), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n258), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT68), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n343), .A2(G77), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n369), .C1(G77), .C2(new_n242), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n275), .A2(G232), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n274), .B(new_n371), .C1(new_n213), .C2(new_n275), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n280), .C1(G107), .C2(new_n274), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n266), .A2(G244), .A3(new_n267), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(new_n269), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n375), .A2(G200), .ZN(new_n378));
  OR3_X1    g0178(.A1(new_n370), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n298), .A2(new_n350), .A3(new_n362), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n211), .A2(new_n275), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n274), .B(new_n381), .C1(G232), .C2(new_n275), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n280), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n266), .A2(G238), .A3(new_n267), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n386), .A2(new_n387), .A3(new_n269), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n386), .B2(new_n269), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT13), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n385), .B(new_n392), .C1(new_n388), .C2(new_n389), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G190), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n391), .A2(KEYINPUT72), .A3(new_n393), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT72), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n390), .A2(new_n397), .A3(KEYINPUT13), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(G200), .A3(new_n398), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n252), .A2(new_n210), .B1(new_n249), .B2(new_n202), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n219), .A2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n258), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT11), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n402), .A2(new_n403), .B1(new_n212), .B2(new_n246), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n402), .A2(new_n403), .ZN(new_n405));
  INV_X1    g0205(.A(G13), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(G1), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n401), .ZN(new_n408));
  XOR2_X1   g0208(.A(new_n408), .B(KEYINPUT12), .Z(new_n409));
  NOR3_X1   g0209(.A1(new_n404), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n395), .A2(new_n399), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n396), .A2(G169), .A3(new_n398), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(KEYINPUT73), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n394), .A2(G179), .ZN(new_n416));
  INV_X1    g0216(.A(new_n414), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n396), .A2(G169), .A3(new_n398), .A4(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n410), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n411), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n375), .A2(G179), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT69), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n375), .A2(new_n353), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n370), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n380), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n219), .B(G87), .C1(new_n310), .C2(new_n311), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT22), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT84), .B(G116), .ZN(new_n431));
  INV_X1    g0231(.A(new_n249), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT23), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n219), .B2(G107), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(KEYINPUT23), .A3(G20), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n431), .A2(new_n432), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n274), .A2(KEYINPUT22), .A3(new_n219), .A4(G87), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n430), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT90), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT90), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n437), .A2(new_n430), .A3(new_n438), .A4(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(KEYINPUT24), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT24), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n439), .A2(KEYINPUT90), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n258), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G257), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G1698), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n448), .B1(G250), .B2(G1698), .C1(new_n310), .C2(new_n311), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G294), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n279), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G45), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G1), .ZN(new_n454));
  NAND2_X1  g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n266), .A2(new_n458), .A3(G264), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n222), .A2(G45), .ZN(new_n460));
  INV_X1    g0260(.A(new_n457), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(new_n455), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G274), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n452), .A2(new_n459), .A3(new_n376), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n459), .ZN(new_n465));
  INV_X1    g0265(.A(new_n463), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n465), .A2(new_n451), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n467), .B2(G200), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n407), .A2(G20), .A3(new_n435), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT25), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n222), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n245), .A2(new_n471), .A3(new_n242), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n245), .A2(KEYINPUT79), .A3(new_n471), .A4(new_n242), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n470), .B1(new_n477), .B2(G107), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n446), .A2(new_n468), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n452), .A2(new_n459), .A3(new_n260), .A4(new_n463), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n467), .B2(G169), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n446), .B2(new_n478), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT91), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n446), .A2(new_n478), .ZN(new_n484));
  INV_X1    g0284(.A(new_n481), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT91), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n446), .A2(new_n468), .A3(new_n478), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n325), .A2(G107), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n251), .A2(G77), .ZN(new_n492));
  OR2_X1    g0292(.A1(KEYINPUT6), .A2(G97), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT78), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(new_n493), .B2(new_n494), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n435), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n498), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(G107), .A3(new_n496), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n501), .A3(G20), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n491), .A2(new_n492), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n258), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n242), .A2(G97), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G97), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n476), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(G250), .B1(new_n310), .B2(new_n311), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT80), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n275), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(new_n275), .C1(new_n310), .C2(new_n311), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n512), .B1(new_n518), .B2(KEYINPUT80), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G244), .ZN(new_n521));
  OAI211_X1 g0321(.A(KEYINPUT80), .B(new_n512), .C1(new_n312), .C2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n517), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n280), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n266), .A2(new_n458), .A3(G257), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n463), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n353), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n519), .A2(new_n514), .A3(new_n516), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n279), .B1(new_n530), .B2(new_n522), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT81), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n525), .A2(new_n463), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n525), .B2(new_n463), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT83), .ZN(new_n536));
  NOR4_X1   g0336(.A1(new_n531), .A2(new_n535), .A3(new_n536), .A4(G179), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n526), .A2(KEYINPUT81), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n525), .A2(new_n463), .A3(new_n532), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n523), .A2(new_n280), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT83), .B1(new_n540), .B2(new_n260), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n510), .B(new_n529), .C1(new_n537), .C2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT82), .B1(new_n531), .B2(new_n535), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n538), .A2(new_n539), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n524), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n546), .A3(G200), .ZN(new_n547));
  AOI211_X1 g0347(.A(new_n505), .B(new_n508), .C1(new_n503), .C2(new_n258), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n524), .A2(G190), .A3(new_n527), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n542), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n272), .A2(new_n273), .B1(new_n213), .B2(new_n275), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n521), .A2(G1698), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n431), .A2(G33), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n279), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g0356(.A1(new_n460), .A2(G274), .ZN(new_n557));
  INV_X1    g0357(.A(G250), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n460), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n557), .A2(new_n266), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n260), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n274), .A2(new_n219), .A3(G68), .ZN(new_n563));
  INV_X1    g0363(.A(G87), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n507), .A3(new_n435), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n383), .A2(new_n219), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT19), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n249), .B2(new_n507), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n563), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n258), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n363), .A2(new_n242), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n476), .C2(new_n364), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n562), .B(new_n573), .C1(G169), .C2(new_n561), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n474), .A2(G87), .A3(new_n475), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n575), .A2(new_n571), .A3(new_n572), .ZN(new_n576));
  OAI21_X1  g0376(.A(G200), .B1(new_n556), .B2(new_n560), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n554), .A2(new_n555), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n280), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT85), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n557), .A2(new_n266), .A3(new_n559), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(G190), .A4(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n552), .A2(new_n553), .B1(G33), .B2(new_n431), .ZN(new_n583));
  OAI211_X1 g0383(.A(G190), .B(new_n581), .C1(new_n583), .C2(new_n279), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT85), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n576), .A2(new_n577), .A3(new_n582), .A4(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n574), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n447), .A2(new_n275), .ZN(new_n588));
  INV_X1    g0388(.A(G264), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G1698), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n590), .C1(new_n310), .C2(new_n311), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n272), .A2(G303), .A3(new_n273), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(KEYINPUT87), .A3(new_n592), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n280), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n266), .A2(new_n458), .A3(G270), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT86), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n266), .A2(new_n458), .A3(KEYINPUT86), .A4(G270), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n597), .A2(new_n602), .A3(new_n463), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(KEYINPUT21), .A3(G169), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n279), .B1(new_n593), .B2(new_n594), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n466), .B1(new_n605), .B2(new_n596), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(G179), .A3(new_n602), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT88), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n515), .B(new_n219), .C1(G33), .C2(new_n507), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n258), .B(new_n610), .C1(new_n431), .C2(new_n219), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT20), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n611), .A2(new_n612), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n611), .A2(new_n609), .A3(new_n612), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n431), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(G20), .A3(new_n407), .ZN(new_n619));
  INV_X1    g0419(.A(new_n472), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G116), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n608), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n353), .B1(new_n606), .B2(new_n602), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g0425(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n617), .A2(new_n621), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n603), .A2(G200), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n606), .A2(G190), .A3(new_n602), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n619), .A4(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n587), .A2(new_n623), .A3(new_n627), .A4(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n490), .A2(new_n551), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n427), .A2(new_n633), .ZN(G372));
  INV_X1    g0434(.A(KEYINPUT92), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n560), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n581), .A2(KEYINPUT92), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n556), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n579), .A2(new_n581), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n638), .A2(G169), .B1(new_n639), .B2(G179), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT93), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n562), .B(KEYINPUT93), .C1(G169), .C2(new_n638), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n573), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n524), .A2(new_n545), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n536), .B1(new_n646), .B2(G179), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n540), .A2(KEYINPUT83), .A3(new_n260), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n587), .A3(new_n529), .A4(new_n510), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n623), .A2(new_n486), .A3(new_n627), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n652), .A2(new_n488), .A3(new_n542), .A4(new_n550), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n638), .A2(new_n328), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(new_n576), .A3(new_n585), .A4(new_n582), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n645), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n645), .B(new_n651), .C1(new_n653), .C2(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n656), .A2(KEYINPUT26), .A3(new_n542), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n427), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT94), .Z(new_n660));
  INV_X1    g0460(.A(new_n411), .ZN(new_n661));
  INV_X1    g0461(.A(new_n425), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n419), .B2(new_n420), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n362), .B1(new_n663), .B2(new_n349), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n295), .A2(new_n297), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n287), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(G369));
  AND2_X1   g0467(.A1(new_n623), .A2(new_n627), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n406), .A2(G20), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n222), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n622), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n668), .A2(new_n631), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n668), .B2(new_n676), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT95), .ZN(new_n679));
  INV_X1    g0479(.A(G330), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n675), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n446), .B2(new_n478), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n490), .A2(new_n683), .B1(new_n486), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n483), .A2(new_n489), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n668), .A2(new_n675), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n482), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n223), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n565), .A2(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n218), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  INV_X1    g0500(.A(new_n607), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n465), .A2(new_n451), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n524), .A2(new_n561), .A3(new_n527), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n704), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n702), .A4(new_n701), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n638), .A2(G179), .ZN(new_n708));
  INV_X1    g0508(.A(new_n467), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n646), .A2(new_n708), .A3(new_n709), .A4(new_n603), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n705), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n711), .A2(new_n712), .A3(new_n675), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n711), .B2(new_n675), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n551), .A2(new_n632), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n686), .A3(new_n682), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT96), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT96), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n633), .A2(new_n719), .A3(new_n682), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n715), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n680), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n682), .B1(new_n657), .B2(new_n658), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n645), .A2(new_n655), .ZN(new_n726));
  INV_X1    g0526(.A(new_n542), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(KEYINPUT26), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT26), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n650), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT97), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT97), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n650), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n645), .B1(new_n653), .B2(new_n656), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n675), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n722), .B1(new_n725), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n699), .B1(new_n739), .B2(G1), .ZN(G364));
  NAND2_X1  g0540(.A1(new_n669), .A2(G45), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n695), .A2(G1), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n681), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n679), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(G330), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n219), .A2(new_n376), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n260), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G58), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n274), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n328), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G87), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n219), .A2(G190), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n752), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G107), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n260), .A2(new_n328), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n747), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n755), .B(new_n759), .C1(new_n210), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n756), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n751), .B(new_n762), .C1(G68), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n219), .B1(new_n766), .B2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G97), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n756), .A2(new_n766), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT32), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n771), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n756), .A2(new_n748), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n765), .B(new_n775), .C1(new_n202), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  INV_X1    g0580(.A(G329), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n757), .A2(new_n780), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n779), .B(new_n782), .C1(G303), .C2(new_n754), .ZN(new_n783));
  INV_X1    g0583(.A(new_n761), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G326), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n768), .A2(G294), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n312), .B1(new_n749), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT33), .B(G317), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(new_n764), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n783), .A2(new_n785), .A3(new_n786), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n777), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n220), .B1(G20), .B2(new_n353), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n793), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n693), .A2(new_n274), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n218), .A2(G45), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(new_n237), .C2(new_n453), .ZN(new_n800));
  INV_X1    g0600(.A(G355), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n274), .A2(new_n223), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n800), .B1(G116), .B2(new_n223), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n792), .A2(new_n793), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n796), .B(KEYINPUT98), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n745), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n746), .B1(new_n742), .B2(new_n806), .ZN(G396));
  NAND2_X1  g0607(.A1(new_n370), .A2(new_n675), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n370), .A2(new_n377), .A3(new_n378), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n425), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n425), .A2(new_n675), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n723), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n379), .A2(new_n808), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n812), .B1(new_n816), .B2(new_n425), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n817), .B(new_n682), .C1(new_n657), .C2(new_n658), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n722), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n742), .ZN(new_n821));
  INV_X1    g0621(.A(new_n749), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G143), .A2(new_n822), .B1(new_n764), .B2(G150), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n824), .B2(new_n761), .C1(new_n771), .C2(new_n776), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n758), .A2(G68), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n825), .A2(new_n826), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n274), .B1(new_n770), .B2(new_n830), .C1(new_n210), .C2(new_n753), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G58), .B2(new_n768), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n753), .A2(new_n435), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n757), .A2(new_n564), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n763), .A2(new_n780), .B1(new_n770), .B2(new_n778), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(G303), .C2(new_n784), .ZN(new_n837));
  INV_X1    g0637(.A(G294), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n312), .B1(new_n749), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n776), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n431), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n837), .A2(new_n769), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n833), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT100), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n742), .B1(new_n844), .B2(new_n793), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n793), .A2(new_n794), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT99), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n202), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n845), .B(new_n848), .C1(new_n795), .C2(new_n817), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n821), .A2(new_n849), .ZN(G384));
  INV_X1    g0650(.A(new_n715), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n719), .B1(new_n633), .B2(new_n682), .ZN(new_n852));
  AND4_X1   g0652(.A1(new_n719), .A2(new_n716), .A3(new_n686), .A4(new_n682), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n306), .B1(new_n314), .B2(new_n318), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT101), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(KEYINPUT16), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n857), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n306), .B(new_n859), .C1(new_n314), .C2(new_n318), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n858), .A2(new_n258), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n673), .B1(new_n861), .B2(new_n344), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n356), .A2(new_n361), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(new_n349), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n359), .A2(new_n360), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n673), .B(KEYINPUT102), .Z(new_n866));
  NAND2_X1  g0666(.A1(new_n359), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n865), .A2(new_n867), .A3(new_n868), .A4(new_n345), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n327), .A2(new_n341), .A3(new_n344), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n355), .B1(new_n861), .B2(new_n344), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n870), .A2(new_n862), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n869), .B1(new_n872), .B2(new_n868), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n864), .A2(new_n873), .A3(KEYINPUT38), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n864), .B2(new_n873), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n410), .A2(new_n682), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n421), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n420), .B(new_n675), .C1(new_n419), .C2(new_n411), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n814), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n854), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n865), .A2(new_n867), .A3(new_n345), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(new_n868), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n867), .B1(new_n362), .B2(new_n350), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n864), .A2(new_n873), .A3(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n854), .A2(new_n891), .A3(new_n881), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n721), .A2(new_n426), .A3(new_n380), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n680), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT39), .B1(new_n889), .B2(new_n890), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n874), .A2(new_n875), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(KEYINPUT39), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n419), .A2(new_n420), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n675), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n877), .B(new_n411), .C1(new_n420), .C2(new_n419), .ZN(new_n903));
  INV_X1    g0703(.A(new_n880), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n818), .B2(new_n813), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n876), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n362), .A2(new_n866), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n738), .A2(new_n427), .A3(new_n725), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n666), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n896), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n222), .B2(new_n669), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n499), .A2(new_n501), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT35), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n219), .B(new_n220), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n917), .B(G116), .C1(new_n916), .C2(new_n915), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT36), .ZN(new_n919));
  OAI21_X1  g0719(.A(G77), .B1(new_n750), .B2(new_n212), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n920), .A2(new_n218), .B1(G50), .B2(new_n212), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(G1), .A3(new_n406), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n914), .A2(new_n919), .A3(new_n922), .ZN(G367));
  NOR2_X1   g0723(.A1(new_n548), .A2(new_n682), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n551), .A2(new_n924), .B1(new_n542), .B2(new_n682), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT103), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n688), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT42), .ZN(new_n931));
  INV_X1    g0731(.A(new_n929), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n727), .B1(new_n932), .B2(new_n482), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n675), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n685), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n932), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n576), .A2(new_n682), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n645), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n726), .B2(new_n937), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n936), .B1(new_n934), .B2(new_n941), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n945), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n694), .B(new_n949), .Z(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n932), .A2(new_n691), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n929), .A2(new_n690), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT44), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n953), .A2(new_n935), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n935), .B1(new_n953), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n688), .B1(new_n684), .B2(new_n687), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n681), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n739), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n956), .A2(new_n957), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n951), .B1(new_n962), .B2(new_n739), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n741), .A2(G1), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n947), .B(new_n948), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n798), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n797), .B1(new_n223), .B2(new_n364), .C1(new_n233), .C2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(G303), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n749), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n312), .B1(new_n776), .B2(new_n780), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(G107), .C2(new_n768), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n784), .A2(G311), .ZN(new_n972));
  INV_X1    g0772(.A(G317), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n763), .A2(new_n838), .B1(new_n770), .B2(new_n973), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n618), .A2(new_n753), .A3(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT46), .B1(new_n753), .B2(new_n206), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n757), .A2(new_n507), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n971), .A2(new_n972), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n758), .A2(G77), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n274), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT106), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n749), .A2(new_n250), .B1(new_n767), .B2(new_n212), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT105), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n753), .A2(new_n750), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n776), .A2(new_n210), .B1(new_n770), .B2(new_n824), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(G143), .C2(new_n784), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n763), .A2(new_n771), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n980), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT47), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n742), .B1(new_n992), .B2(new_n793), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n967), .B(new_n993), .C1(new_n940), .C2(new_n805), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n965), .A2(new_n994), .ZN(G387));
  NAND2_X1  g0795(.A1(new_n959), .A2(new_n964), .ZN(new_n996));
  INV_X1    g0796(.A(new_n770), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n997), .A2(G326), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G311), .A2(new_n764), .B1(new_n822), .B2(G317), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n968), .B2(new_n776), .C1(new_n787), .C2(new_n761), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT48), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n780), .B2(new_n767), .C1(new_n838), .C2(new_n753), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT49), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n274), .B(new_n998), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .C1(new_n618), .C2(new_n757), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n763), .A2(new_n248), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n754), .A2(G77), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n776), .B2(new_n212), .C1(new_n250), .C2(new_n770), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G159), .B2(new_n784), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n768), .A2(new_n363), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n312), .B(new_n978), .C1(G50), .C2(new_n822), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1005), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n798), .B1(new_n230), .B2(new_n453), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n696), .B2(new_n802), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n212), .A2(new_n202), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n248), .A2(G50), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G116), .B(new_n565), .C1(new_n1017), .C2(KEYINPUT50), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1018), .B(new_n453), .C1(KEYINPUT50), .C2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1015), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(G107), .B2(new_n223), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1013), .A2(new_n793), .B1(new_n797), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1022), .B(new_n743), .C1(new_n684), .C2(new_n805), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n694), .B1(new_n959), .B2(new_n739), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n996), .B(new_n1023), .C1(new_n961), .C2(new_n1024), .ZN(G393));
  NAND2_X1  g0825(.A1(new_n956), .A2(new_n957), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n695), .B1(new_n1026), .B2(new_n960), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1027), .A2(new_n962), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n929), .A2(new_n796), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n797), .B1(new_n507), .B2(new_n223), .C1(new_n240), .C2(new_n966), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n763), .A2(new_n210), .B1(new_n776), .B2(new_n248), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT107), .Z(new_n1032));
  OAI22_X1  g0832(.A1(new_n761), .A2(new_n250), .B1(new_n749), .B2(new_n771), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT51), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n274), .B1(new_n757), .B2(new_n564), .C1(new_n212), .C2(new_n753), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G77), .B2(new_n768), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n997), .A2(G143), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n763), .A2(new_n968), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n776), .A2(new_n838), .B1(new_n770), .B2(new_n787), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G283), .C2(new_n754), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n761), .A2(new_n973), .B1(new_n749), .B2(new_n778), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT52), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n274), .B1(new_n768), .B2(new_n431), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n1043), .A3(new_n759), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n742), .B1(new_n1046), .B2(new_n793), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1029), .A2(new_n1030), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n964), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(new_n1026), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1028), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(G390));
  NAND2_X1  g0852(.A1(new_n818), .A2(new_n813), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n905), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n901), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n728), .A2(new_n731), .A3(new_n733), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n682), .B(new_n811), .C1(new_n1056), .C2(new_n735), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n905), .B1(new_n1057), .B2(new_n813), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n901), .B1(new_n889), .B2(new_n890), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1055), .A2(new_n899), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n722), .A2(KEYINPUT108), .A3(new_n881), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n898), .A2(KEYINPUT39), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n901), .A2(new_n906), .B1(new_n1065), .B2(new_n897), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n812), .B1(new_n737), .B2(new_n811), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1059), .B1(new_n1067), .B2(new_n905), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1068), .A3(new_n1062), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1064), .A2(new_n964), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT110), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n894), .A2(G330), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n666), .A3(new_n910), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n854), .A2(G330), .A3(new_n881), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n721), .A2(new_n680), .A3(new_n814), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n1054), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n1053), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1074), .B(new_n1067), .C1(new_n1075), .C2(new_n1054), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1073), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT109), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1064), .B(new_n1069), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n854), .A2(G330), .A3(new_n817), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1083), .A2(new_n905), .B1(new_n722), .B2(new_n881), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1053), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1078), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1073), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1082), .A2(new_n1088), .A3(KEYINPUT109), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1081), .A2(new_n1089), .A3(new_n694), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n749), .A2(new_n830), .B1(new_n757), .B2(new_n210), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G137), .B2(new_n764), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n761), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n312), .B(new_n1094), .C1(G159), .C2(new_n768), .ZN(new_n1095));
  INV_X1    g0895(.A(G125), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(KEYINPUT54), .B(G143), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT111), .Z(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1095), .B1(new_n1096), .B2(new_n770), .C1(new_n776), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n754), .A2(G150), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n761), .A2(new_n780), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n749), .A2(new_n206), .B1(new_n770), .B2(new_n838), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(G97), .C2(new_n840), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n202), .B2(new_n767), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n764), .A2(G107), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n755), .A2(new_n1107), .A3(new_n828), .A4(new_n312), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1100), .A2(new_n1102), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1109), .A2(new_n793), .B1(new_n248), .B2(new_n847), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n743), .B(new_n1110), .C1(new_n899), .C2(new_n795), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1071), .A2(new_n1090), .A3(new_n1111), .ZN(G378));
  OAI21_X1  g0912(.A(new_n817), .B1(new_n903), .B2(new_n904), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n721), .A2(new_n1113), .A3(new_n898), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n892), .C1(new_n1114), .C2(KEYINPUT40), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT55), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n298), .A2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(KEYINPUT55), .B(new_n287), .C1(new_n295), .C2(new_n297), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n259), .A2(new_n673), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT56), .Z(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1121), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n298), .A2(new_n1116), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n1118), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1115), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1128), .A2(new_n884), .A3(G330), .A4(new_n892), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n909), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT116), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n909), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT116), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1127), .A2(new_n909), .A3(new_n1129), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT57), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1064), .A2(new_n1086), .A3(new_n1069), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n1087), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n694), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT117), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT114), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n909), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1132), .B2(KEYINPUT115), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1132), .A2(KEYINPUT115), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n909), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(KEYINPUT115), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1146), .B1(new_n1149), .B2(new_n1145), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1139), .A2(new_n1087), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1138), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT117), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1141), .A2(new_n1154), .A3(new_n694), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1143), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1150), .A2(new_n1049), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1128), .A2(new_n794), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n846), .A2(new_n210), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G128), .A2(new_n822), .B1(new_n764), .B2(G132), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1096), .B2(new_n761), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G150), .B2(new_n768), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n824), .B2(new_n776), .C1(new_n753), .C2(new_n1099), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT59), .Z(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n997), .B2(G124), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G33), .B1(new_n758), .B2(G159), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G58), .A2(new_n758), .B1(new_n997), .B2(G283), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n274), .A2(G41), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1007), .A3(new_n1169), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT112), .Z(new_n1171));
  AOI22_X1  g0971(.A1(G97), .A2(new_n764), .B1(new_n822), .B2(G107), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n206), .B2(new_n761), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G68), .B2(new_n768), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1171), .B(new_n1174), .C1(new_n364), .C2(new_n776), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT58), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n210), .B1(new_n310), .B2(G41), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1167), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT113), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n742), .B1(new_n1179), .B2(new_n793), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1158), .A2(new_n1159), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1157), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1156), .A2(new_n1183), .ZN(G375));
  NAND2_X1  g0984(.A1(new_n905), .A2(new_n794), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n981), .A2(new_n312), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT119), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n761), .A2(new_n838), .B1(new_n770), .B2(new_n968), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n618), .A2(new_n763), .B1(new_n753), .B2(new_n507), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1010), .B1(new_n780), .B2(new_n749), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT120), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n435), .C2(new_n776), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G137), .A2(new_n822), .B1(new_n754), .B2(G159), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n1093), .B2(new_n770), .C1(new_n250), .C2(new_n776), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G50), .B2(new_n768), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n312), .B1(new_n758), .B2(G58), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n763), .C2(new_n1099), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n784), .A2(G132), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT121), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1193), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1201), .A2(new_n793), .B1(new_n212), .B2(new_n847), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1185), .A2(new_n743), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1086), .B2(new_n964), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n950), .B(KEYINPUT118), .Z(new_n1205));
  NAND2_X1  g1005(.A1(new_n1088), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1204), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT122), .ZN(G381));
  NAND2_X1  g1009(.A1(G378), .A2(KEYINPUT123), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT123), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1071), .A2(new_n1090), .A3(new_n1211), .A4(new_n1111), .ZN(new_n1212));
  AOI21_X1  g1012(.A(G375), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1051), .A2(new_n994), .A3(new_n965), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n1213), .A2(new_n674), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(G407), .A2(G213), .A3(new_n1218), .ZN(G409));
  NAND2_X1  g1019(.A1(G390), .A2(G387), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1215), .ZN(new_n1221));
  XOR2_X1   g1021(.A(G393), .B(G396), .Z(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1222), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1220), .A2(new_n1215), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1156), .A2(G378), .A3(new_n1183), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1137), .A2(new_n964), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1181), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT124), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT115), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1134), .A2(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1232), .A2(new_n1147), .B1(new_n1144), .B2(new_n909), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1151), .B(new_n1205), .C1(new_n1233), .C2(new_n1146), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1228), .A2(new_n1235), .A3(new_n1181), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1230), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1227), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n674), .A2(G213), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1207), .A2(KEYINPUT60), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n694), .A3(new_n1088), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1207), .A2(KEYINPUT60), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1204), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G384), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT125), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n695), .B1(new_n1207), .B2(KEYINPUT60), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n1088), .C1(KEYINPUT60), .C2(new_n1207), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(G384), .A4(new_n1204), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1247), .A2(new_n1248), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1240), .A2(new_n1241), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT126), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT126), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1240), .A2(new_n1257), .A3(new_n1241), .A4(new_n1254), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT62), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n674), .A2(G213), .A3(G2897), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1253), .B(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1255), .A2(KEYINPUT62), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1226), .B1(new_n1259), .B2(new_n1265), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1240), .A2(new_n1241), .A3(new_n1254), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1226), .B1(new_n1267), .B2(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1263), .B(new_n1268), .C1(new_n1269), .C2(KEYINPUT63), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1266), .A2(new_n1270), .ZN(G405));
  NAND2_X1  g1071(.A1(G375), .A2(new_n1238), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1226), .A2(KEYINPUT127), .A3(new_n1227), .A4(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(KEYINPUT127), .A3(new_n1227), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT127), .B1(new_n1272), .B2(new_n1227), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(new_n1254), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1273), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(G402));
endmodule


