//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n211), .B1(new_n215), .B2(KEYINPUT0), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n216), .B1(KEYINPUT0), .B2(new_n215), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT64), .Z(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n218), .A2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(new_n208), .ZN(new_n251));
  INV_X1    g0051(.A(G223), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n252), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n261), .A2(G222), .A3(new_n258), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(new_n261), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n251), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(new_n250), .B2(new_n208), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n209), .A2(KEYINPUT68), .A3(new_n249), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n273), .A2(G226), .A3(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n271), .A2(new_n272), .A3(G274), .A4(new_n276), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G179), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT75), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT70), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(new_n208), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(new_n284), .B2(new_n208), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT72), .A2(G58), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n290), .A2(KEYINPUT8), .ZN(new_n291));
  AND3_X1   g0091(.A1(KEYINPUT71), .A2(KEYINPUT72), .A3(G58), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT8), .B1(KEYINPUT71), .B2(G58), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(new_n295), .A3(G33), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n289), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n289), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G1), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G20), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G50), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT73), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n303), .A2(new_n307), .B1(G50), .B2(new_n302), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT74), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI221_X1 g0110(.A(KEYINPUT74), .B1(G50), .B2(new_n302), .C1(new_n303), .C2(new_n307), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n299), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n281), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n283), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT9), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n312), .B(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n281), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(G200), .B2(new_n281), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n318), .B1(new_n317), .B2(new_n321), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n315), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n261), .A2(G226), .A3(new_n258), .ZN(new_n326));
  INV_X1    g0126(.A(G97), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n261), .A2(G232), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n326), .B1(new_n253), .B2(new_n327), .C1(new_n328), .C2(new_n258), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n251), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n271), .A2(new_n277), .A3(new_n272), .A4(G238), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n332), .A2(new_n279), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n330), .B2(new_n333), .ZN(new_n336));
  OAI21_X1  g0136(.A(G169), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT14), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n330), .A2(new_n333), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT13), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT77), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT77), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n341), .A2(G179), .A3(new_n343), .A4(new_n334), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n334), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(G169), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n338), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n289), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n295), .A2(G33), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n350), .A2(new_n267), .B1(new_n295), .B2(G68), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT78), .ZN(new_n352));
  INV_X1    g0152(.A(new_n297), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n351), .A2(new_n352), .B1(new_n202), .B2(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n351), .A2(new_n352), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT11), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n302), .A2(KEYINPUT12), .A3(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n284), .A2(new_n208), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n302), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n220), .B1(new_n304), .B2(G20), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n360), .A2(new_n361), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n358), .A2(new_n359), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n348), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n345), .B2(G200), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n341), .A2(G190), .A3(new_n343), .A4(new_n334), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n305), .A2(G77), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n364), .A2(new_n373), .B1(G77), .B2(new_n302), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G20), .A2(G77), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT15), .B(G87), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT8), .B(G58), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n375), .B1(new_n376), .B2(new_n350), .C1(new_n353), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n374), .B1(new_n378), .B2(new_n362), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT76), .ZN(new_n380));
  INV_X1    g0180(.A(new_n251), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n262), .A2(new_n263), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT69), .B1(new_n261), .B2(G1698), .ZN(new_n383));
  OAI21_X1  g0183(.A(G238), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G107), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n328), .A2(G1698), .B1(new_n385), .B2(new_n261), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n381), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n273), .A2(G244), .A3(new_n277), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n279), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n380), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n221), .B1(new_n260), .B2(new_n264), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n251), .B1(new_n392), .B2(new_n386), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n389), .A2(new_n279), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(KEYINPUT76), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n379), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n391), .A2(new_n395), .A3(new_n313), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n319), .B1(new_n391), .B2(new_n395), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G200), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n379), .C1(new_n403), .C2(new_n396), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n369), .A2(new_n372), .A3(new_n400), .A4(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n325), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n302), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n291), .B(new_n407), .C1(new_n292), .C2(new_n293), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n294), .A2(new_n305), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n303), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT81), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT81), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n412), .B(new_n408), .C1(new_n303), .C2(new_n409), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n261), .A2(new_n415), .A3(G20), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT7), .B1(new_n257), .B2(new_n295), .ZN(new_n417));
  OAI21_X1  g0217(.A(G68), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT16), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT80), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT79), .ZN(new_n421));
  OR2_X1    g0221(.A1(KEYINPUT71), .A2(G58), .ZN(new_n422));
  NAND2_X1  g0222(.A1(KEYINPUT71), .A2(G58), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n220), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(G20), .B1(new_n424), .B2(new_n201), .ZN(new_n425));
  INV_X1    g0225(.A(G159), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n353), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n421), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(KEYINPUT71), .A2(G58), .ZN(new_n430));
  NOR2_X1   g0230(.A1(KEYINPUT71), .A2(G58), .ZN(new_n431));
  OAI21_X1  g0231(.A(G68), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n295), .B1(new_n432), .B2(new_n206), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n433), .A2(KEYINPUT79), .A3(new_n427), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n420), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT79), .B1(new_n433), .B2(new_n427), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT71), .B(G58), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n201), .B1(new_n437), .B2(G68), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n421), .B(new_n428), .C1(new_n438), .C2(new_n295), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n439), .A3(KEYINPUT80), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n419), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n436), .A2(new_n418), .A3(new_n439), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT16), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n362), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n414), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n254), .A2(new_n256), .A3(G226), .A4(G1698), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n254), .A2(new_n256), .A3(G223), .A4(new_n258), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n448), .B(new_n449), .C1(new_n253), .C2(new_n222), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n251), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n271), .A2(new_n277), .A3(new_n272), .A4(G232), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n279), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n452), .A2(new_n454), .A3(new_n397), .ZN(new_n455));
  INV_X1    g0255(.A(new_n454), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n313), .B1(new_n456), .B2(new_n451), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n446), .A2(new_n447), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n451), .A2(new_n319), .A3(new_n279), .A4(new_n453), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT82), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n403), .B1(new_n452), .B2(new_n454), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n456), .A2(new_n464), .A3(new_n319), .A4(new_n451), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n414), .C1(new_n441), .C2(new_n445), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT17), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n411), .A2(new_n413), .ZN(new_n470));
  INV_X1    g0270(.A(new_n419), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n436), .A2(new_n439), .A3(KEYINPUT80), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT80), .B1(new_n436), .B2(new_n439), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n363), .B1(new_n442), .B2(new_n443), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT18), .B1(new_n476), .B2(new_n458), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(KEYINPUT17), .A3(new_n466), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n460), .A2(new_n469), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n479), .A2(KEYINPUT83), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(KEYINPUT83), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n406), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n254), .A2(new_n256), .A3(G244), .A4(G1698), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT86), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n261), .A2(KEYINPUT86), .A3(G244), .A4(G1698), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n261), .A2(G238), .A3(new_n258), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n304), .A2(G45), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n490), .A2(G274), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n223), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n489), .A2(new_n251), .B1(new_n273), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G190), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n222), .A2(new_n327), .A3(new_n385), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT87), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(new_n222), .A3(new_n327), .A4(new_n385), .ZN(new_n499));
  NAND3_X1  g0299(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n497), .A2(new_n499), .B1(new_n295), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n254), .A2(new_n256), .A3(new_n295), .A4(G68), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n350), .A2(new_n327), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(KEYINPUT19), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n362), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n407), .A2(new_n376), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n304), .A2(G33), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n289), .A2(G87), .A3(new_n302), .A4(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n495), .B(new_n509), .C1(new_n403), .C2(new_n494), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n489), .A2(new_n251), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n493), .A2(new_n273), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n313), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n494), .A2(new_n397), .ZN(new_n515));
  INV_X1    g0315(.A(new_n288), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(new_n302), .A3(new_n286), .A4(new_n507), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n505), .B(new_n506), .C1(new_n376), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n407), .A2(new_n385), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n520), .B(KEYINPUT25), .ZN(new_n521));
  INV_X1    g0321(.A(new_n517), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(G107), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n254), .A2(new_n256), .A3(new_n295), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n261), .A2(new_n526), .A3(new_n295), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT24), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n487), .A2(G20), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT23), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n295), .B2(G107), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n385), .A2(KEYINPUT23), .A3(G20), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n529), .B1(new_n528), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n362), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n523), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n261), .A2(G250), .A3(new_n258), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n261), .A2(G257), .A3(G1698), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n251), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT5), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n274), .ZN(new_n546));
  NAND2_X1  g0346(.A1(KEYINPUT5), .A2(G41), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n490), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(new_n271), .A3(G274), .A4(new_n272), .ZN(new_n549));
  INV_X1    g0349(.A(new_n547), .ZN(new_n550));
  NOR2_X1   g0350(.A1(KEYINPUT5), .A2(G41), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n304), .B(G45), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n273), .A2(G264), .A3(new_n552), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n544), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n397), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G169), .B2(new_n554), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n510), .B(new_n519), .C1(new_n539), .C2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n552), .A2(new_n271), .A3(G270), .A4(new_n272), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n549), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G264), .ZN(new_n561));
  INV_X1    g0361(.A(G303), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n262), .A2(new_n561), .B1(new_n562), .B2(new_n261), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n261), .A2(G257), .A3(new_n258), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT88), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n261), .A2(KEYINPUT88), .A3(G257), .A4(new_n258), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n560), .B1(new_n568), .B2(new_n381), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G200), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n566), .A2(new_n567), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n259), .A2(G264), .B1(G303), .B2(new_n257), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n559), .B1(new_n573), .B2(new_n251), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G190), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G283), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n576), .B(new_n295), .C1(G33), .C2(new_n327), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n577), .B(new_n362), .C1(new_n295), .C2(G116), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT20), .ZN(new_n579));
  INV_X1    g0379(.A(G116), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n301), .A2(G20), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n507), .A2(G116), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n364), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n570), .A2(new_n575), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  OAI21_X1  g0386(.A(G169), .B1(new_n579), .B2(new_n583), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n574), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n584), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n589), .A2(KEYINPUT21), .A3(new_n569), .A4(G169), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n397), .B(new_n559), .C1(new_n573), .C2(new_n251), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n589), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n585), .A2(new_n588), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n552), .A2(new_n271), .A3(new_n272), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n251), .A2(new_n543), .B1(new_n594), .B2(G264), .ZN(new_n595));
  AOI21_X1  g0395(.A(G200), .B1(new_n595), .B2(new_n549), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n319), .A2(new_n544), .A3(new_n549), .A4(new_n553), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n523), .B(new_n537), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n417), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n295), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n385), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n602), .A2(new_n327), .A3(G107), .ZN(new_n603));
  XNOR2_X1  g0403(.A(G97), .B(G107), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n605), .A2(new_n295), .B1(new_n267), .B2(new_n353), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n362), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n301), .A2(G20), .A3(new_n327), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n608), .B(KEYINPUT84), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n517), .A2(new_n327), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n552), .A2(new_n271), .A3(G257), .A4(new_n272), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n549), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n254), .A2(new_n256), .A3(G244), .A4(new_n258), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT4), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n576), .A4(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n613), .B1(new_n251), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n397), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n251), .ZN(new_n622));
  INV_X1    g0422(.A(new_n613), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n313), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n611), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(G190), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n609), .B1(new_n327), .B2(new_n517), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n604), .A2(new_n602), .ZN(new_n629));
  INV_X1    g0429(.A(new_n603), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(G20), .B1(G77), .B2(new_n297), .ZN(new_n632));
  OAI21_X1  g0432(.A(G107), .B1(new_n416), .B2(new_n417), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n628), .B1(new_n634), .B2(new_n362), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n403), .B1(new_n622), .B2(new_n623), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n627), .B(new_n635), .C1(KEYINPUT85), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT85), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n598), .B(new_n626), .C1(new_n637), .C2(new_n639), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n557), .A2(new_n593), .A3(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n482), .A2(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n460), .A2(new_n477), .ZN(new_n643));
  INV_X1    g0443(.A(new_n372), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n369), .B1(new_n644), .B2(new_n400), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n469), .A2(new_n478), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n323), .A2(new_n324), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n315), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT91), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT91), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n651), .B(new_n315), .C1(new_n647), .C2(new_n648), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n482), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT89), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n509), .B(new_n655), .C1(new_n403), .C2(new_n494), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n403), .B1(new_n511), .B2(new_n512), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT89), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n656), .A2(new_n659), .A3(new_n495), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n611), .A2(new_n621), .A3(new_n625), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .A4(new_n519), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n510), .A2(new_n519), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT26), .B1(new_n664), .B2(new_n626), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n665), .A3(new_n519), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n539), .A2(new_n556), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n590), .A2(new_n592), .A3(new_n588), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n660), .A2(new_n519), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n640), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT90), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT90), .B1(new_n640), .B2(new_n670), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n666), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n653), .B1(new_n654), .B2(new_n675), .ZN(G369));
  INV_X1    g0476(.A(new_n301), .ZN(new_n677));
  OR3_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .A3(G20), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT27), .B1(new_n677), .B2(G20), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n584), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT92), .B1(new_n668), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n593), .B2(new_n684), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n668), .A2(KEYINPUT92), .A3(new_n684), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G330), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n667), .A2(new_n683), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n538), .A2(new_n682), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(new_n598), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n694), .B2(new_n667), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n668), .A2(new_n683), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n692), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT93), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(KEYINPUT93), .A3(new_n692), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n697), .A2(new_n704), .ZN(G399));
  NAND3_X1  g0505(.A1(new_n497), .A2(new_n580), .A3(new_n499), .ZN(new_n706));
  INV_X1    g0506(.A(new_n213), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n706), .A2(new_n708), .A3(new_n304), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT94), .ZN(new_n710));
  INV_X1    g0510(.A(new_n207), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n709), .A2(new_n710), .B1(new_n711), .B2(new_n708), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n710), .B2(new_n709), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT26), .B1(new_n670), .B2(new_n626), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n661), .A2(new_n510), .A3(new_n519), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n715), .B(new_n519), .C1(KEYINPUT26), .C2(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n669), .A2(new_n640), .A3(new_n670), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT29), .B(new_n683), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n675), .A2(new_n682), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n641), .A2(new_n683), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n620), .A2(new_n595), .A3(new_n494), .ZN(new_n723));
  OAI211_X1 g0523(.A(G179), .B(new_n560), .C1(new_n568), .C2(new_n381), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n574), .A2(new_n554), .A3(new_n620), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n494), .A2(G179), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n725), .A2(KEYINPUT30), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n723), .B2(new_n724), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n683), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n722), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT95), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT95), .B(new_n729), .C1(new_n723), .C2(new_n724), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n728), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT31), .B1(new_n740), .B2(new_n682), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n735), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n721), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n714), .B1(new_n744), .B2(G1), .ZN(G364));
  NOR2_X1   g0545(.A1(new_n300), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n304), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n708), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n690), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n688), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n751), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n749), .B(KEYINPUT96), .Z(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n208), .B1(G20), .B2(new_n313), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n707), .A2(new_n257), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT97), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(G355), .B(KEYINPUT98), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n767), .A2(new_n768), .B1(G116), .B2(new_n213), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT99), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n244), .A2(new_n275), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n261), .B(new_n707), .C1(new_n711), .C2(new_n275), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n769), .A2(KEYINPUT99), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n764), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n295), .A2(G179), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G87), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n775), .A2(new_n319), .A3(G200), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n778), .B(new_n261), .C1(new_n385), .C2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT100), .Z(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n295), .A2(new_n397), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G200), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n785), .A2(KEYINPUT32), .B1(new_n788), .B2(new_n437), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n787), .A2(new_n403), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n319), .A2(G179), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n295), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n789), .B1(new_n202), .B2(new_n791), .C1(new_n327), .C2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n786), .A2(new_n319), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n786), .A2(new_n782), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n796), .A2(G68), .B1(new_n798), .B2(G77), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(KEYINPUT32), .B2(new_n785), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n781), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n788), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n802), .A2(new_n803), .B1(new_n779), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n793), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(G294), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(KEYINPUT33), .B(G317), .Z(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n795), .A2(new_n808), .B1(new_n797), .B2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n261), .B(new_n810), .C1(G329), .C2(new_n784), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n790), .A2(G326), .B1(new_n777), .B2(G303), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n801), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n761), .B(new_n774), .C1(new_n762), .C2(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n750), .A2(new_n753), .B1(new_n759), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  OAI21_X1  g0618(.A(new_n379), .B1(new_n396), .B2(new_n403), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n819), .A2(new_n401), .B1(new_n379), .B2(new_n683), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n400), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n398), .A2(new_n399), .A3(new_n683), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n720), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n637), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n661), .B1(new_n826), .B2(new_n638), .ZN(new_n827));
  INV_X1    g0627(.A(new_n519), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n509), .B1(new_n403), .B2(new_n494), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(KEYINPUT89), .B1(G190), .B2(new_n494), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n656), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n827), .A2(new_n831), .A3(new_n672), .A4(new_n598), .ZN(new_n832));
  INV_X1    g0632(.A(new_n669), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n832), .A2(new_n674), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n666), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT102), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n404), .A2(new_n400), .A3(new_n683), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT102), .B1(new_n675), .B2(new_n838), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n825), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n743), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n844), .B(new_n845), .C1(new_n708), .C2(new_n748), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n796), .A2(G150), .B1(new_n798), .B2(G159), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n788), .A2(G143), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n791), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  INV_X1    g0654(.A(new_n437), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n261), .B1(new_n783), .B2(new_n854), .C1(new_n793), .C2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n779), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(G68), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n202), .B2(new_n776), .ZN(new_n859));
  NOR4_X1   g0659(.A1(new_n852), .A2(new_n853), .A3(new_n856), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n779), .A2(new_n222), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G303), .B2(new_n790), .ZN(new_n862));
  INV_X1    g0662(.A(G294), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(new_n802), .ZN(new_n864));
  XOR2_X1   g0664(.A(KEYINPUT101), .B(G283), .Z(new_n865));
  OAI21_X1  g0665(.A(new_n257), .B1(new_n795), .B2(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n797), .A2(new_n580), .B1(new_n783), .B2(new_n809), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n793), .A2(new_n327), .B1(new_n776), .B2(new_n385), .ZN(new_n868));
  NOR4_X1   g0668(.A1(new_n864), .A2(new_n866), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n762), .B1(new_n860), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n762), .A2(new_n754), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n761), .B1(new_n267), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n870), .B(new_n872), .C1(new_n824), .C2(new_n755), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n846), .A2(new_n873), .ZN(G384));
  NOR2_X1   g0674(.A1(new_n746), .A2(new_n304), .ZN(new_n875));
  INV_X1    g0675(.A(new_n418), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n435), .B2(new_n440), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n474), .B(new_n349), .C1(new_n877), .C2(KEYINPUT16), .ZN(new_n878));
  INV_X1    g0678(.A(new_n410), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n458), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n467), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT104), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT104), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n441), .A2(new_n289), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n418), .B1(new_n472), .B2(new_n473), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n443), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n410), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n883), .B(new_n467), .C1(new_n887), .C2(new_n458), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n887), .A2(new_n680), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n882), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n446), .A2(new_n459), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n680), .B(KEYINPUT105), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n446), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n892), .A2(new_n894), .A3(new_n895), .A4(new_n467), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n887), .A2(new_n680), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n479), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n896), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n890), .B2(KEYINPUT37), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n905), .B2(new_n900), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n494), .A2(new_n595), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n591), .A2(new_n908), .A3(KEYINPUT30), .A4(new_n620), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n554), .A2(new_n620), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n569), .A3(new_n727), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n737), .B2(new_n738), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT106), .B1(new_n913), .B2(new_n683), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT106), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n740), .A2(new_n915), .A3(new_n682), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(new_n916), .A3(new_n732), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n641), .A2(new_n683), .B1(new_n740), .B2(new_n733), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n368), .A2(new_n682), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n369), .A2(new_n372), .A3(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n368), .B(new_n682), .C1(new_n644), .C2(new_n348), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n823), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT40), .B1(new_n907), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n899), .A2(KEYINPUT38), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n891), .B2(new_n896), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n892), .A2(new_n894), .A3(new_n467), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT37), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n896), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n479), .A2(new_n446), .A3(new_n893), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT107), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n931), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n901), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT107), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n905), .C2(new_n926), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n919), .A2(new_n923), .A3(KEYINPUT40), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n933), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT108), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT108), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n933), .A2(new_n937), .A3(new_n938), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n925), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n482), .A2(new_n919), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n689), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n903), .A2(new_n906), .A3(KEYINPUT39), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n369), .A2(new_n682), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n927), .B2(new_n932), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n837), .B1(new_n836), .B2(new_n839), .ZN(new_n952));
  AOI211_X1 g0752(.A(KEYINPUT102), .B(new_n838), .C1(new_n834), .C2(new_n835), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n822), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n921), .A2(new_n922), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(new_n907), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n893), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n643), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n951), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n482), .B(new_n719), .C1(KEYINPUT29), .C2(new_n720), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n653), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n875), .B1(new_n946), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n962), .B2(new_n946), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n210), .A2(new_n580), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n631), .B(KEYINPUT103), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT35), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n968), .B2(new_n967), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT36), .Z(new_n971));
  NAND3_X1  g0771(.A1(new_n711), .A2(G77), .A3(new_n432), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(G50), .B2(new_n220), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(G1), .A3(new_n300), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n964), .A2(new_n971), .A3(new_n974), .ZN(G367));
  NOR2_X1   g0775(.A1(new_n707), .A2(new_n261), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n240), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n763), .B1(new_n213), .B2(new_n376), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n760), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n791), .A2(new_n809), .B1(new_n779), .B2(new_n327), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n802), .A2(new_n562), .B1(new_n385), .B2(new_n793), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(G317), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n865), .A2(new_n797), .B1(new_n783), .B2(new_n983), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n261), .B(new_n984), .C1(G294), .C2(new_n796), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n777), .A2(KEYINPUT46), .A3(G116), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT46), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n776), .B2(new_n580), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n982), .A2(new_n985), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n261), .B1(new_n779), .B2(new_n267), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT113), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n795), .A2(new_n426), .B1(new_n797), .B2(new_n202), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G137), .B2(new_n784), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G68), .A2(new_n806), .B1(new_n790), .B2(G143), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n788), .A2(G150), .B1(new_n777), .B2(new_n437), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n989), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT47), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n979), .B1(new_n998), .B2(new_n762), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n509), .A2(new_n683), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n828), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n670), .B2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n999), .B1(new_n1002), .B2(new_n757), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT114), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1002), .A2(KEYINPUT109), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(KEYINPUT109), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n699), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n827), .B1(new_n635), .B2(new_n683), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n661), .A2(new_n682), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT42), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT111), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n667), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n626), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1015), .A2(KEYINPUT42), .B1(new_n683), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1010), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1014), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n697), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1021), .A2(new_n1022), .A3(new_n1010), .ZN(new_n1027));
  AND3_X1   g0827(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1026), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n702), .A2(new_n703), .A3(new_n1025), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT44), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n704), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1034));
  AOI21_X1  g0834(.A(KEYINPUT45), .B1(new_n704), .B2(new_n1014), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n696), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n695), .A2(new_n698), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT112), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n690), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n690), .A2(new_n1039), .ZN(new_n1041));
  AND3_X1   g0841(.A1(new_n1040), .A2(new_n1011), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1011), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n744), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n697), .A3(new_n1033), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1037), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n744), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n708), .B(KEYINPUT41), .Z(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n748), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1005), .B1(new_n1030), .B2(new_n1054), .ZN(G387));
  OR2_X1    g0855(.A1(new_n1045), .A2(new_n744), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1056), .A2(new_n708), .A3(new_n1046), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n796), .A2(G311), .B1(new_n798), .B2(G303), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n802), .B2(new_n983), .C1(new_n803), .C2(new_n791), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n793), .A2(new_n865), .B1(new_n776), .B2(new_n863), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT49), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n261), .B1(new_n784), .B2(G326), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n580), .B2(new_n779), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(G150), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n261), .B1(new_n783), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G68), .B2(new_n798), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n788), .A2(G50), .B1(new_n857), .B2(G97), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n294), .A2(new_n796), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n793), .A2(new_n376), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n791), .A2(new_n426), .B1(new_n776), .B2(new_n267), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n762), .B1(new_n1068), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n976), .B1(new_n236), .B2(new_n275), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n706), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n767), .ZN(new_n1081));
  OR3_X1    g0881(.A1(new_n377), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT50), .B1(new_n377), .B2(G50), .ZN(new_n1083));
  AOI21_X1  g0883(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1081), .A2(new_n1085), .B1(new_n385), .B2(new_n707), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1078), .B(new_n760), .C1(new_n764), .C2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n695), .B2(new_n756), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1045), .B2(new_n748), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1057), .A2(new_n1089), .ZN(G393));
  NAND3_X1  g0890(.A1(new_n1037), .A2(new_n748), .A3(new_n1049), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n763), .B1(new_n327), .B2(new_n213), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n247), .B2(new_n976), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n865), .A2(new_n776), .B1(new_n783), .B2(new_n803), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT115), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n257), .B1(new_n385), .B2(new_n779), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1095), .B2(new_n1094), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT116), .Z(new_n1098));
  AOI22_X1  g0898(.A1(G311), .A2(new_n788), .B1(new_n790), .B2(G317), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT52), .Z(new_n1100));
  OAI22_X1  g0900(.A1(new_n795), .A2(new_n562), .B1(new_n797), .B2(new_n863), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G116), .B2(new_n806), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(KEYINPUT117), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G150), .A2(new_n790), .B1(new_n788), .B2(G159), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT51), .Z(new_n1106));
  OAI22_X1  g0906(.A1(new_n795), .A2(new_n202), .B1(new_n797), .B2(new_n377), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n257), .B(new_n1107), .C1(G143), .C2(new_n784), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n793), .A2(new_n267), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n861), .B(new_n1109), .C1(G68), .C2(new_n777), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1103), .A2(KEYINPUT117), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1104), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n761), .B(new_n1093), .C1(new_n1113), .C2(new_n762), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n757), .B2(new_n1014), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1091), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1036), .A2(new_n696), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n697), .B1(new_n1048), .B2(new_n1033), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1046), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n1050), .A3(new_n708), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT118), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1050), .A3(KEYINPUT118), .A4(new_n708), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(G390));
  AOI21_X1  g0925(.A(new_n689), .B1(new_n917), .B2(new_n918), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n923), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n954), .A2(new_n955), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n948), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1129), .A2(new_n1130), .B1(new_n950), .B2(new_n947), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n683), .B(new_n821), .C1(new_n717), .C2(new_n718), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n822), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n948), .B1(new_n1133), .B2(new_n955), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n933), .A3(new_n937), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1128), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(G330), .B(new_n824), .C1(new_n735), .C2(new_n741), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n955), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n947), .A2(new_n950), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n948), .B1(new_n954), .B2(new_n955), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1135), .B(new_n1140), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(new_n747), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1141), .A2(new_n755), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n871), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n760), .B1(new_n294), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(G125), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n795), .A2(new_n849), .B1(new_n783), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n257), .B(new_n1150), .C1(new_n798), .C2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n776), .A2(new_n1069), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G159), .A2(new_n806), .B1(new_n788), .B2(G132), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n790), .A2(G128), .B1(new_n857), .B2(G50), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1153), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G97), .A2(new_n798), .B1(new_n784), .B2(G294), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n261), .B1(new_n796), .B2(G107), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n778), .A4(new_n858), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1109), .B1(G116), .B2(new_n788), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n804), .B2(new_n791), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1158), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1148), .B1(new_n1164), .B2(new_n762), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1145), .B1(new_n1146), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n482), .A2(new_n1126), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n960), .A2(new_n653), .A3(new_n1167), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n954), .B1(new_n1169), .B2(new_n1128), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1133), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1126), .A2(new_n824), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1140), .B(new_n1171), .C1(new_n955), .C2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1168), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1144), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1137), .A2(new_n1174), .A3(new_n1143), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(new_n708), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1166), .A2(new_n1178), .ZN(G378));
  INV_X1    g0979(.A(new_n958), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n841), .A2(new_n840), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1139), .B1(new_n1181), .B2(new_n822), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n1182), .B2(new_n907), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT121), .B1(new_n1183), .B2(new_n951), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n951), .A2(new_n956), .A3(KEYINPUT121), .A4(new_n958), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n940), .A2(new_n942), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n925), .A2(new_n689), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n312), .A2(new_n680), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n325), .B(new_n1191), .Z(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1192), .B(new_n1193), .Z(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1190), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(new_n1189), .A3(new_n1194), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1187), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n959), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1188), .A2(new_n1189), .A3(new_n1194), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1194), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1194), .A2(new_n754), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n749), .B1(new_n1147), .B2(G50), .ZN(new_n1205));
  AOI21_X1  g1005(.A(G50), .B1(new_n253), .B2(new_n274), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n261), .B2(G41), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n855), .A2(new_n779), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G107), .B2(new_n788), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n580), .B2(new_n791), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n274), .B(new_n257), .C1(new_n795), .C2(new_n327), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n797), .A2(new_n376), .B1(new_n783), .B2(new_n804), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n793), .A2(new_n220), .B1(new_n776), .B2(new_n267), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1207), .B1(new_n1214), .B2(KEYINPUT58), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT119), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(KEYINPUT58), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n795), .A2(new_n854), .B1(new_n797), .B2(new_n849), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G150), .B2(new_n806), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n788), .A2(G128), .B1(new_n777), .B2(new_n1152), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT120), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1222), .A2(KEYINPUT120), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1221), .B1(new_n1149), .B2(new_n791), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n857), .A2(G159), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G33), .B(G41), .C1(new_n784), .C2(G124), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1219), .B1(new_n1216), .B2(new_n1215), .C1(new_n1227), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1205), .B1(new_n1232), .B2(new_n762), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1203), .A2(new_n748), .B1(new_n1204), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1168), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1177), .B2(new_n1236), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1200), .A2(new_n1201), .A3(new_n1199), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n959), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n708), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1177), .A2(new_n1236), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1234), .B1(new_n1241), .B2(new_n1243), .ZN(G375));
  AND2_X1   g1044(.A1(new_n1173), .A2(new_n1170), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1168), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1175), .A2(new_n1246), .A3(new_n1053), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n760), .B1(G68), .B2(new_n1147), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n776), .A2(new_n327), .B1(new_n783), .B2(new_n562), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT122), .Z(new_n1250));
  OAI21_X1  g1050(.A(new_n257), .B1(new_n797), .B2(new_n385), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G116), .B2(new_n796), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1075), .B1(G77), .B2(new_n857), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G283), .A2(new_n788), .B1(new_n790), .B2(G294), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1252), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n790), .A2(G132), .B1(new_n796), .B2(new_n1152), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n849), .B2(new_n802), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT123), .Z(new_n1258));
  AOI22_X1  g1058(.A1(new_n777), .A2(G159), .B1(new_n784), .B2(G128), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT124), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n257), .B(new_n1208), .C1(G150), .C2(new_n798), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(new_n202), .C2(new_n793), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1255), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1248), .B1(new_n1263), .B2(new_n762), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n955), .B2(new_n755), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1245), .B2(new_n747), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1247), .A2(new_n1267), .ZN(G381));
  INV_X1    g1068(.A(G387), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1271), .A2(G381), .A3(G384), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1124), .A3(new_n1272), .ZN(new_n1273));
  OR3_X1    g1073(.A1(new_n1273), .A2(G375), .A3(G378), .ZN(G407));
  AND2_X1   g1074(.A1(new_n1166), .A2(new_n1178), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n681), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(G375), .C2(new_n1278), .ZN(G409));
  OAI211_X1 g1079(.A(G378), .B(new_n1234), .C1(new_n1241), .C2(new_n1243), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT121), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n959), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1185), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1200), .A2(new_n1283), .A3(new_n1201), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1053), .B(new_n1242), .C1(new_n1284), .C2(new_n1239), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1204), .A2(new_n1233), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n748), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1275), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1277), .B1(new_n1280), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n846), .A2(new_n1291), .A3(new_n873), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1246), .B1(new_n1293), .B2(new_n1174), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1245), .A2(KEYINPUT60), .A3(new_n1168), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1295), .A2(new_n708), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n1266), .B(new_n1292), .C1(new_n1294), .C2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1266), .B1(new_n1296), .B2(new_n1294), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1291), .B1(new_n846), .B2(new_n873), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1292), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1290), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1280), .A2(new_n1289), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1276), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G2897), .B(new_n1277), .C1(new_n1297), .C2(new_n1301), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1298), .B1(KEYINPUT125), .B2(G384), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1277), .A2(G2897), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1309), .B(new_n1310), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(G387), .A2(new_n1124), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G387), .A2(new_n1124), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G393), .A2(G396), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  OR3_X1    g1119(.A1(new_n1319), .A2(KEYINPUT126), .A3(new_n1270), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT126), .B1(new_n1319), .B2(new_n1270), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1316), .A2(new_n1317), .A3(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(G387), .A2(new_n1124), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1321), .B1(new_n1324), .B2(new_n1315), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1302), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1305), .A2(new_n1314), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1290), .A2(new_n1329), .A3(new_n1302), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1331), .B1(new_n1290), .B2(new_n1312), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1329), .B1(new_n1290), .B2(new_n1302), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1330), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1328), .B1(new_n1334), .B2(new_n1326), .ZN(G405));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1302), .A2(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(KEYINPUT127), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1275), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1339), .B1(new_n1340), .B2(new_n1280), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1339), .A2(new_n1280), .A3(new_n1340), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1342), .A2(new_n1323), .A3(new_n1325), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1343), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1326), .B1(new_n1345), .B2(new_n1341), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(G402));
endmodule


