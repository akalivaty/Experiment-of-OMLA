//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n958, new_n959;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT29), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR3_X1   g015(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT27), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n227));
  OAI211_X1 g026(.A(KEYINPUT67), .B(G183gat), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n224), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n225), .A2(G183gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n230), .A2(new_n234), .A3(KEYINPUT28), .A4(new_n229), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n220), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  INV_X1    g036(.A(G169gat), .ZN(new_n238));
  INV_X1    g037(.A(G176gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n229), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT24), .A3(new_n219), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n219), .A2(KEYINPUT24), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n246), .B(new_n215), .C1(KEYINPUT64), .C2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n242), .A2(new_n244), .A3(new_n215), .A4(new_n245), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n242), .A2(new_n244), .A3(KEYINPUT64), .A4(new_n245), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT25), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n213), .B1(new_n236), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT73), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n253), .A2(KEYINPUT73), .A3(new_n254), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n254), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT25), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n249), .B1(KEYINPUT25), .B2(new_n250), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n251), .A3(KEYINPUT65), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n236), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n266), .A2(KEYINPUT72), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT72), .B1(new_n266), .B2(new_n267), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n260), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n212), .B1(new_n259), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n212), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n260), .A2(KEYINPUT29), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n268), .B2(new_n269), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n236), .A2(new_n254), .A3(new_n252), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n205), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT74), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n281), .B(new_n205), .C1(new_n271), .C2(new_n277), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT75), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n278), .A2(new_n280), .ZN(new_n285));
  INV_X1    g084(.A(new_n258), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT73), .B1(new_n253), .B2(new_n254), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n267), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n236), .B1(new_n264), .B2(new_n265), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT72), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n254), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n272), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n273), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(new_n291), .B2(new_n293), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n212), .B1(new_n297), .B2(new_n275), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(new_n205), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n285), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n279), .A2(new_n302), .A3(new_n280), .A4(new_n282), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT88), .ZN(new_n305));
  INV_X1    g104(.A(G120gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G113gat), .ZN(new_n307));
  INV_X1    g106(.A(G113gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G120gat), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT1), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n311));
  INV_X1    g110(.A(G134gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(G127gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(G127gat), .B(G134gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(new_n311), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT69), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n317), .B(new_n313), .C1(new_n314), .C2(new_n311), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n310), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n307), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n309), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n323), .A2(new_n324), .A3(new_n314), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327));
  INV_X1    g126(.A(G141gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(G148gat), .ZN(new_n329));
  INV_X1    g128(.A(G148gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n329), .B(new_n331), .C1(G141gat), .C2(new_n330), .ZN(new_n332));
  AND2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n332), .B(new_n335), .C1(new_n333), .C2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n333), .A2(new_n336), .ZN(new_n338));
  XNOR2_X1  g137(.A(G141gat), .B(G148gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(KEYINPUT2), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n319), .A2(new_n341), .A3(new_n325), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(KEYINPUT4), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT80), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n326), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n337), .A2(new_n351), .A3(new_n340), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n349), .A2(new_n350), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n353), .B(new_n352), .C1(new_n319), .C2(new_n325), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OR3_X1    g156(.A1(new_n343), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n348), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n326), .A2(new_n342), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n363), .A2(new_n346), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n364), .A2(new_n361), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(KEYINPUT39), .A3(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G57gat), .B(G85gat), .Z(new_n367));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT78), .B(KEYINPUT0), .Z(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT79), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n369), .B(new_n371), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n366), .B(new_n373), .C1(KEYINPUT39), .C2(new_n362), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n305), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n346), .B(new_n344), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n343), .A2(new_n361), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n357), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT5), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n364), .B2(new_n361), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n361), .A2(KEYINPUT5), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n348), .A2(new_n357), .A3(new_n358), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT87), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT87), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(new_n387), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n376), .A2(KEYINPUT40), .B1(new_n372), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n373), .B1(new_n362), .B2(KEYINPUT39), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n362), .A2(new_n365), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(KEYINPUT39), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT88), .B1(new_n393), .B2(KEYINPUT86), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT40), .B1(new_n393), .B2(KEYINPUT88), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n304), .A2(new_n390), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n352), .A2(new_n213), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n212), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT84), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n212), .A2(KEYINPUT29), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n401), .A2(KEYINPUT83), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n351), .B1(new_n401), .B2(KEYINPUT83), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n341), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G228gat), .ZN(new_n406));
  INV_X1    g205(.A(G233gat), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI211_X1 g207(.A(new_n406), .B(new_n407), .C1(new_n401), .C2(new_n341), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n353), .A3(new_n399), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT31), .B(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(G22gat), .ZN(new_n415));
  INV_X1    g214(.A(G22gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(KEYINPUT85), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n411), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n271), .B2(new_n277), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT38), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n259), .A2(new_n270), .A3(new_n212), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n274), .A2(new_n272), .A3(new_n276), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT37), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n422), .A2(new_n423), .A3(new_n204), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(new_n279), .A3(new_n282), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n205), .B1(new_n299), .B2(new_n421), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n295), .A2(KEYINPUT37), .A3(new_n298), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n423), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n382), .A2(new_n373), .A3(new_n384), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n389), .B2(new_n372), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n385), .A2(KEYINPUT6), .A3(new_n372), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n373), .B1(new_n382), .B2(new_n384), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n420), .B1(new_n432), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n397), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT81), .B1(new_n435), .B2(new_n440), .ZN(new_n446));
  INV_X1    g245(.A(new_n440), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n434), .A4(new_n433), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n446), .A2(new_n449), .A3(new_n441), .A4(new_n439), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n284), .A2(new_n450), .A3(new_n301), .A4(new_n303), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  INV_X1    g251(.A(G71gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(KEYINPUT71), .B(G99gat), .Z(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(new_n455), .Z(new_n456));
  INV_X1    g255(.A(G227gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(new_n407), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n289), .A2(new_n349), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n292), .A2(new_n326), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n456), .B1(new_n462), .B2(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n461), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n458), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(KEYINPUT32), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT32), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT34), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n464), .A2(new_n458), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n467), .B2(new_n469), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n467), .A2(new_n469), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n470), .ZN(new_n477));
  INV_X1    g276(.A(new_n463), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n479), .A3(KEYINPUT36), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n473), .A2(new_n474), .A3(new_n463), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n478), .B1(new_n477), .B2(new_n472), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n451), .A2(new_n420), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n482), .A2(new_n483), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n419), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT35), .B1(new_n451), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n284), .A2(new_n301), .A3(new_n303), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n475), .A2(new_n479), .A3(new_n490), .A4(new_n419), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(new_n443), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n445), .A2(new_n485), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G230gat), .A2(G233gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G71gat), .B(G78gat), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n499), .B(new_n500), .Z(new_n501));
  XOR2_X1   g300(.A(G99gat), .B(G106gat), .Z(new_n502));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT98), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT98), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(G99gat), .A3(G106gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n506), .A3(KEYINPUT8), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n510), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT99), .B(new_n502), .C1(new_n508), .C2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n513), .ZN(new_n515));
  INV_X1    g314(.A(new_n502), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n507), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT99), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n502), .B1(new_n508), .B2(new_n513), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT10), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n499), .B(new_n500), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n519), .A3(new_n517), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT101), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT101), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n521), .A2(new_n527), .A3(new_n522), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n520), .A2(new_n514), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(KEYINPUT10), .A3(new_n523), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n496), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n521), .A2(new_n524), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n496), .ZN(new_n535));
  XNOR2_X1  g334(.A(G120gat), .B(G148gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n531), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n526), .B2(new_n528), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n535), .B1(new_n542), .B2(new_n496), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n538), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(G15gat), .B(G22gat), .Z(new_n546));
  INV_X1    g345(.A(G1gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G15gat), .B(G22gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(KEYINPUT16), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G8gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT94), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n549), .B2(new_n550), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n552), .B1(new_n548), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n546), .A2(new_n555), .A3(new_n547), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n557), .A2(KEYINPUT93), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT93), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n556), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(G8gat), .A3(new_n558), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n557), .A2(KEYINPUT93), .A3(new_n558), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n553), .A2(KEYINPUT94), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n553), .A2(KEYINPUT94), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n567), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT95), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT15), .ZN(new_n573));
  INV_X1    g372(.A(G50gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G43gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT89), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT90), .B(G50gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(G43gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n573), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G43gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G50gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n575), .A3(KEYINPUT15), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G29gat), .ZN(new_n585));
  INV_X1    g384(.A(G36gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT14), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT14), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(G29gat), .B2(G36gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(G29gat), .A2(G36gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n583), .ZN(new_n594));
  NAND2_X1  g393(.A1(KEYINPUT91), .A2(KEYINPUT17), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT91), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n591), .B1(new_n580), .B2(new_n583), .ZN(new_n600));
  INV_X1    g399(.A(new_n594), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n596), .B(new_n597), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n563), .A2(new_n572), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n561), .A2(new_n593), .A3(new_n594), .ZN(new_n605));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT96), .Z(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT18), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n594), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n571), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n607), .B(KEYINPUT13), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n604), .A2(KEYINPUT18), .A3(new_n605), .A4(new_n607), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618));
  INV_X1    g417(.A(G197gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT11), .B(G169gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n610), .A2(new_n623), .A3(new_n615), .A4(new_n616), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n523), .A2(KEYINPUT21), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n554), .B(new_n631), .C1(new_n560), .C2(new_n559), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(G183gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n571), .A2(new_n223), .A3(new_n631), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n523), .A2(KEYINPUT21), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n633), .B2(new_n634), .ZN(new_n638));
  INV_X1    g437(.A(G231gat), .ZN(new_n639));
  OAI22_X1  g438(.A1(new_n637), .A2(new_n638), .B1(new_n639), .B2(new_n407), .ZN(new_n640));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G211gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n633), .A2(new_n634), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n635), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n639), .A2(new_n407), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n640), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n643), .B1(new_n640), .B2(new_n648), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n630), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n640), .A2(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n642), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n640), .A2(new_n648), .A3(new_n643), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n629), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G134gat), .B(G162gat), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n599), .B2(new_n602), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT100), .B1(new_n599), .B2(new_n602), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n611), .A2(new_n530), .ZN(new_n663));
  OAI22_X1  g462(.A1(new_n530), .A2(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G190gat), .B(G218gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n664), .B2(new_n667), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n659), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n658), .A3(new_n668), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n651), .A2(new_n655), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR4_X1   g475(.A1(new_n494), .A2(new_n545), .A3(new_n628), .A4(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n450), .B(KEYINPUT102), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n304), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT16), .B(G8gat), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n684), .A2(KEYINPUT104), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(KEYINPUT104), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n682), .B2(G8gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(KEYINPUT42), .ZN(new_n690));
  OAI22_X1  g489(.A1(new_n687), .A2(new_n689), .B1(new_n682), .B2(new_n690), .ZN(G1325gat));
  AOI21_X1  g490(.A(G15gat), .B1(new_n677), .B2(new_n486), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n484), .A2(new_n480), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT105), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n692), .B1(new_n677), .B2(new_n696), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n677), .A2(new_n420), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n651), .A2(new_n655), .ZN(new_n701));
  INV_X1    g500(.A(new_n545), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n627), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n494), .A2(new_n674), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n585), .A3(new_n679), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n445), .A2(new_n485), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n488), .A2(new_n493), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n674), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(KEYINPUT44), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n494), .B2(new_n674), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n703), .B(KEYINPUT106), .Z(new_n714));
  NAND3_X1  g513(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT107), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n711), .A2(new_n713), .A3(new_n717), .A4(new_n714), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n678), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n706), .B1(new_n719), .B2(new_n585), .ZN(G1328gat));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n718), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n304), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT108), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n724), .A3(new_n304), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(G36gat), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n704), .A2(new_n586), .A3(new_n304), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT46), .Z(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(G1329gat));
  OAI21_X1  g528(.A(G43gat), .B1(new_n715), .B2(new_n693), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n704), .A2(new_n581), .A3(new_n486), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(KEYINPUT47), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n731), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n721), .A2(new_n694), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(G43gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n735), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g535(.A(new_n578), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n715), .B2(new_n419), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n704), .A2(new_n578), .A3(new_n420), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(KEYINPUT48), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n739), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n721), .A2(new_n420), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(new_n737), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(G1331gat));
  NOR4_X1   g544(.A1(new_n494), .A2(new_n702), .A3(new_n627), .A4(new_n676), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n679), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n304), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n750), .B(new_n751), .Z(G1333gat));
  NAND3_X1  g551(.A1(new_n746), .A2(new_n453), .A3(new_n486), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n746), .A2(new_n694), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n453), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g555(.A1(new_n746), .A2(new_n420), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n494), .A2(new_n674), .ZN(new_n759));
  INV_X1    g558(.A(new_n701), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n627), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n759), .A2(KEYINPUT51), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT51), .B1(new_n759), .B2(new_n761), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n702), .ZN(new_n765));
  INV_X1    g564(.A(G85gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n766), .A3(new_n679), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n760), .A2(new_n702), .A3(new_n627), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n711), .A2(new_n713), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(new_n679), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n766), .B2(new_n770), .ZN(G1336gat));
  INV_X1    g570(.A(G92gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n304), .A2(new_n772), .A3(new_n545), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n762), .B2(new_n763), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n711), .A2(new_n713), .A3(new_n304), .A4(new_n768), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G92gat), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n773), .B(KEYINPUT110), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n762), .B2(new_n763), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n777), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT111), .B(new_n779), .C1(new_n782), .C2(new_n778), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n778), .B1(new_n781), .B2(new_n777), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(G1337gat));
  XOR2_X1   g587(.A(KEYINPUT112), .B(G99gat), .Z(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n765), .A2(new_n486), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n769), .A2(new_n694), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n790), .ZN(G1338gat));
  NAND4_X1  g592(.A1(new_n711), .A2(new_n713), .A3(new_n420), .A4(new_n768), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n702), .A2(new_n419), .A3(G106gat), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT113), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n764), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n542), .B2(new_n496), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n533), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n539), .B1(new_n532), .B2(new_n800), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT55), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n540), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT115), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n532), .A2(new_n800), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n538), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n495), .B(new_n541), .C1(new_n526), .C2(new_n528), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n532), .A2(new_n810), .A3(new_n800), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n804), .A2(new_n813), .A3(new_n540), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n806), .A2(new_n627), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n607), .B1(new_n604), .B2(new_n605), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n613), .A2(new_n614), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n622), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n626), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n545), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n710), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n812), .A3(new_n814), .A4(new_n819), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n674), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n701), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n675), .A2(KEYINPUT114), .A3(new_n702), .A4(new_n628), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n651), .A2(new_n655), .A3(new_n702), .A4(new_n674), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(new_n627), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n678), .A2(new_n487), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n830), .A2(new_n489), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT116), .ZN(new_n833));
  OAI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n628), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n308), .A3(new_n627), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1340gat));
  OAI21_X1  g635(.A(G120gat), .B1(new_n833), .B2(new_n702), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n832), .A2(new_n306), .A3(new_n545), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1341gat));
  AOI21_X1  g638(.A(G127gat), .B1(new_n832), .B2(new_n760), .ZN(new_n840));
  INV_X1    g639(.A(new_n833), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n760), .A2(G127gat), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(G1342gat));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n833), .B2(new_n674), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n832), .A2(new_n312), .A3(new_n710), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT56), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n844), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n848), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n845), .A3(KEYINPUT117), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(G1343gat));
  AOI21_X1  g651(.A(new_n419), .B1(new_n824), .B2(new_n829), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n678), .A2(new_n694), .A3(new_n304), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n328), .A3(new_n627), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n419), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n804), .A2(new_n813), .A3(new_n540), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n813), .B1(new_n804), .B2(new_n540), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(new_n710), .A3(new_n812), .A4(new_n819), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n809), .B2(new_n811), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n627), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n820), .B1(new_n866), .B2(new_n805), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n674), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n760), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n825), .A2(new_n828), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n859), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(KEYINPUT119), .B(new_n859), .C1(new_n869), .C2(new_n870), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n873), .B(new_n874), .C1(KEYINPUT57), .C2(new_n853), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n875), .A2(KEYINPUT120), .A3(new_n854), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT120), .B1(new_n875), .B2(new_n854), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n627), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n857), .B1(new_n878), .B2(G141gat), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n875), .A2(new_n627), .A3(new_n854), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT58), .B1(new_n881), .B2(G141gat), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(KEYINPUT121), .A3(new_n856), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT121), .B1(new_n882), .B2(new_n856), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n879), .A2(new_n880), .B1(new_n883), .B2(new_n884), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n855), .A2(new_n330), .A3(new_n545), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n873), .A2(new_n874), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n853), .A2(KEYINPUT57), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n854), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n875), .A2(KEYINPUT120), .A3(new_n854), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n702), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(KEYINPUT59), .A3(new_n330), .ZN(new_n894));
  XOR2_X1   g693(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n895));
  NOR2_X1   g694(.A1(new_n827), .A2(new_n627), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n858), .B(new_n420), .C1(new_n869), .C2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n830), .A2(new_n420), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(KEYINPUT57), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n545), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n854), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n895), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n886), .B1(new_n894), .B2(new_n904), .ZN(G1345gat));
  AOI21_X1  g704(.A(G155gat), .B1(new_n855), .B2(new_n760), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n701), .B1(new_n891), .B2(new_n892), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g707(.A(G162gat), .B1(new_n855), .B2(new_n710), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n674), .B1(new_n891), .B2(new_n892), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(G162gat), .ZN(G1347gat));
  AOI21_X1  g710(.A(new_n487), .B1(new_n824), .B2(new_n829), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n679), .A2(new_n489), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n628), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(new_n238), .ZN(G1348gat));
  NOR2_X1   g715(.A1(new_n914), .A2(new_n702), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(new_n239), .ZN(G1349gat));
  NAND2_X1  g717(.A1(new_n230), .A2(new_n234), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n914), .A2(new_n701), .ZN(new_n920));
  MUX2_X1   g719(.A(new_n223), .B(new_n919), .S(new_n920), .Z(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT60), .Z(G1350gat));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n923));
  OAI221_X1 g722(.A(G190gat), .B1(KEYINPUT123), .B2(new_n923), .C1(new_n914), .C2(new_n674), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n912), .A2(new_n229), .A3(new_n710), .A4(new_n913), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n925), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G1351gat));
  NOR3_X1   g728(.A1(new_n679), .A2(new_n489), .A3(new_n694), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n897), .B(new_n930), .C1(new_n853), .C2(new_n858), .ZN(new_n931));
  OR3_X1    g730(.A1(new_n931), .A2(KEYINPUT124), .A3(new_n628), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT124), .B1(new_n931), .B2(new_n628), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(G197gat), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n853), .A2(new_n930), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n619), .A3(new_n627), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT125), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n902), .A2(new_n930), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n902), .A2(new_n945), .A3(new_n930), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(G204gat), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(KEYINPUT126), .ZN(new_n949));
  NOR4_X1   g748(.A1(new_n935), .A2(G204gat), .A3(new_n702), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(KEYINPUT126), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n947), .A2(new_n952), .ZN(G1353gat));
  OAI21_X1  g752(.A(G211gat), .B1(new_n931), .B2(new_n701), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT63), .Z(new_n955));
  NAND3_X1  g754(.A1(new_n936), .A2(new_n207), .A3(new_n760), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1354gat));
  OAI21_X1  g756(.A(G218gat), .B1(new_n931), .B2(new_n674), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n936), .A2(new_n208), .A3(new_n710), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1355gat));
endmodule


