

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  XNOR2_X1 U323 ( .A(n433), .B(KEYINPUT48), .ZN(n527) );
  INV_X1 U324 ( .A(n527), .ZN(n529) );
  XOR2_X1 U325 ( .A(n394), .B(n393), .Z(n291) );
  INV_X1 U326 ( .A(KEYINPUT99), .ZN(n391) );
  INV_X1 U327 ( .A(KEYINPUT11), .ZN(n378) );
  XNOR2_X1 U328 ( .A(n391), .B(KEYINPUT36), .ZN(n392) );
  XNOR2_X1 U329 ( .A(n379), .B(n378), .ZN(n388) );
  XNOR2_X1 U330 ( .A(n544), .B(n392), .ZN(n586) );
  XNOR2_X1 U331 ( .A(n388), .B(n387), .ZN(n389) );
  NOR2_X1 U332 ( .A1(n530), .A2(n455), .ZN(n566) );
  XOR2_X1 U333 ( .A(n469), .B(KEYINPUT28), .Z(n532) );
  XOR2_X1 U334 ( .A(n447), .B(n309), .Z(n530) );
  XNOR2_X1 U335 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U336 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT17), .B(KEYINPUT79), .Z(n293) );
  XNOR2_X1 U338 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n292) );
  XNOR2_X1 U339 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U340 ( .A(KEYINPUT19), .B(n294), .Z(n447) );
  XOR2_X1 U341 ( .A(KEYINPUT78), .B(G113GAT), .Z(n296) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(G15GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n308) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G71GAT), .Z(n412) );
  XOR2_X1 U345 ( .A(G176GAT), .B(G99GAT), .Z(n298) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(G190GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U348 ( .A(n412), .B(n299), .Z(n301) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U351 ( .A(n302), .B(KEYINPUT80), .Z(n306) );
  XOR2_X1 U352 ( .A(G127GAT), .B(KEYINPUT0), .Z(n304) );
  XNOR2_X1 U353 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n346) );
  XNOR2_X1 U355 ( .A(n346), .B(KEYINPUT20), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U357 ( .A(n308), .B(n307), .Z(n309) );
  XOR2_X1 U358 ( .A(KEYINPUT82), .B(KEYINPUT23), .Z(n311) );
  XNOR2_X1 U359 ( .A(KEYINPUT22), .B(KEYINPUT83), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U361 ( .A(KEYINPUT87), .B(n312), .Z(n314) );
  NAND2_X1 U362 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U364 ( .A(n315), .B(KEYINPUT24), .Z(n322) );
  XOR2_X1 U365 ( .A(G211GAT), .B(KEYINPUT85), .Z(n317) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n446) );
  XOR2_X1 U368 ( .A(n446), .B(KEYINPUT86), .Z(n319) );
  XOR2_X1 U369 ( .A(G141GAT), .B(G22GAT), .Z(n397) );
  XNOR2_X1 U370 ( .A(n397), .B(KEYINPUT81), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n320), .B(KEYINPUT84), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n324) );
  XNOR2_X1 U374 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n323), .B(KEYINPUT2), .ZN(n345) );
  XOR2_X1 U376 ( .A(n324), .B(n345), .Z(n332) );
  XNOR2_X1 U377 ( .A(G148GAT), .B(KEYINPUT71), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n325), .B(KEYINPUT72), .ZN(n326) );
  XOR2_X1 U379 ( .A(n326), .B(G204GAT), .Z(n328) );
  XNOR2_X1 U380 ( .A(G78GAT), .B(G106GAT), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n422) );
  XOR2_X1 U382 ( .A(G162GAT), .B(KEYINPUT74), .Z(n330) );
  XNOR2_X1 U383 ( .A(G50GAT), .B(G218GAT), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n377) );
  XNOR2_X1 U385 ( .A(n422), .B(n377), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n469) );
  XOR2_X1 U387 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n334) );
  XNOR2_X1 U388 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n341) );
  XOR2_X1 U390 ( .A(G85GAT), .B(G148GAT), .Z(n336) );
  XNOR2_X1 U391 ( .A(G141GAT), .B(G120GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(n337), .B(G162GAT), .Z(n339) );
  XOR2_X1 U394 ( .A(G113GAT), .B(G1GAT), .Z(n399) );
  XNOR2_X1 U395 ( .A(G29GAT), .B(n399), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n350) );
  XOR2_X1 U398 ( .A(KEYINPUT89), .B(KEYINPUT1), .Z(n343) );
  NAND2_X1 U399 ( .A1(G225GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U401 ( .A(n344), .B(KEYINPUT88), .Z(n348) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U404 ( .A(n350), .B(n349), .Z(n468) );
  INV_X1 U405 ( .A(n468), .ZN(n518) );
  XOR2_X1 U406 ( .A(KEYINPUT110), .B(KEYINPUT45), .Z(n351) );
  XNOR2_X1 U407 ( .A(KEYINPUT64), .B(n351), .ZN(n394) );
  XOR2_X1 U408 ( .A(G57GAT), .B(KEYINPUT13), .Z(n411) );
  XOR2_X1 U409 ( .A(G71GAT), .B(G127GAT), .Z(n353) );
  XNOR2_X1 U410 ( .A(G15GAT), .B(G183GAT), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U412 ( .A(n411), .B(n354), .Z(n356) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U415 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n358) );
  XNOR2_X1 U416 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U418 ( .A(n360), .B(n359), .Z(n368) );
  XOR2_X1 U419 ( .A(G211GAT), .B(G155GAT), .Z(n362) );
  XNOR2_X1 U420 ( .A(G22GAT), .B(G78GAT), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U422 ( .A(KEYINPUT76), .B(G64GAT), .Z(n364) );
  XNOR2_X1 U423 ( .A(G8GAT), .B(G1GAT), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U426 ( .A(n368), .B(n367), .Z(n581) );
  INV_X1 U427 ( .A(n581), .ZN(n540) );
  XOR2_X1 U428 ( .A(G29GAT), .B(KEYINPUT66), .Z(n370) );
  XNOR2_X1 U429 ( .A(KEYINPUT8), .B(G43GAT), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n372) );
  XOR2_X1 U431 ( .A(KEYINPUT65), .B(KEYINPUT7), .Z(n371) );
  XOR2_X1 U432 ( .A(n372), .B(n371), .Z(n407) );
  INV_X1 U433 ( .A(n407), .ZN(n376) );
  XOR2_X1 U434 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n374) );
  XNOR2_X1 U435 ( .A(G106GAT), .B(G92GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U437 ( .A(n376), .B(n375), .Z(n390) );
  XNOR2_X1 U438 ( .A(G134GAT), .B(n377), .ZN(n379) );
  XNOR2_X1 U439 ( .A(G99GAT), .B(G85GAT), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n380), .B(KEYINPUT73), .ZN(n419) );
  XOR2_X1 U441 ( .A(G36GAT), .B(G190GAT), .Z(n436) );
  NAND2_X1 U442 ( .A1(n419), .A2(n436), .ZN(n384) );
  INV_X1 U443 ( .A(n419), .ZN(n382) );
  INV_X1 U444 ( .A(n436), .ZN(n381) );
  NAND2_X1 U445 ( .A1(n382), .A2(n381), .ZN(n383) );
  NAND2_X1 U446 ( .A1(n384), .A2(n383), .ZN(n386) );
  AND2_X1 U447 ( .A1(G232GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U449 ( .A(n390), .B(n389), .Z(n544) );
  NOR2_X1 U450 ( .A1(n540), .A2(n586), .ZN(n393) );
  XOR2_X1 U451 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n396) );
  XNOR2_X1 U452 ( .A(G15GAT), .B(G197GAT), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n403) );
  XOR2_X1 U455 ( .A(n399), .B(KEYINPUT29), .Z(n401) );
  NAND2_X1 U456 ( .A1(G229GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U459 ( .A(G169GAT), .B(G8GAT), .Z(n437) );
  XOR2_X1 U460 ( .A(n404), .B(n437), .Z(n406) );
  XNOR2_X1 U461 ( .A(G50GAT), .B(G36GAT), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U463 ( .A(n408), .B(n407), .Z(n533) );
  INV_X1 U464 ( .A(n533), .ZN(n571) );
  XOR2_X1 U465 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n410) );
  XNOR2_X1 U466 ( .A(KEYINPUT68), .B(KEYINPUT70), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n416) );
  XOR2_X1 U468 ( .A(KEYINPUT69), .B(KEYINPUT31), .Z(n414) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U471 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U472 ( .A1(G230GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U474 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U475 ( .A(G176GAT), .B(G92GAT), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n421), .B(G64GAT), .ZN(n444) );
  XNOR2_X1 U477 ( .A(n422), .B(n444), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n576) );
  NOR2_X1 U479 ( .A1(n571), .A2(n576), .ZN(n425) );
  AND2_X1 U480 ( .A1(n291), .A2(n425), .ZN(n426) );
  XOR2_X1 U481 ( .A(n426), .B(KEYINPUT111), .Z(n432) );
  INV_X1 U482 ( .A(n544), .ZN(n557) );
  XNOR2_X1 U483 ( .A(KEYINPUT41), .B(n576), .ZN(n535) );
  INV_X1 U484 ( .A(n535), .ZN(n561) );
  NAND2_X1 U485 ( .A1(n561), .A2(n571), .ZN(n427) );
  XNOR2_X1 U486 ( .A(KEYINPUT46), .B(n427), .ZN(n428) );
  NAND2_X1 U487 ( .A1(n428), .A2(n540), .ZN(n429) );
  NOR2_X1 U488 ( .A1(n557), .A2(n429), .ZN(n430) );
  XOR2_X1 U489 ( .A(KEYINPUT47), .B(n430), .Z(n431) );
  NOR2_X1 U490 ( .A1(n432), .A2(n431), .ZN(n433) );
  XOR2_X1 U491 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n435) );
  XNOR2_X1 U492 ( .A(KEYINPUT92), .B(KEYINPUT90), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U494 ( .A(n436), .B(G218GAT), .Z(n439) );
  XNOR2_X1 U495 ( .A(n437), .B(G204GAT), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U497 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U498 ( .A1(G226GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U500 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n520) );
  NOR2_X1 U503 ( .A1(n527), .A2(n520), .ZN(n452) );
  XOR2_X1 U504 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n450) );
  XNOR2_X1 U505 ( .A(KEYINPUT118), .B(n450), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U507 ( .A1(n518), .A2(n453), .ZN(n569) );
  NOR2_X1 U508 ( .A1(n469), .A2(n569), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n454), .B(KEYINPUT55), .ZN(n455) );
  NAND2_X1 U510 ( .A1(n566), .A2(n557), .ZN(n459) );
  XOR2_X1 U511 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n457) );
  INV_X1 U512 ( .A(G190GAT), .ZN(n456) );
  NOR2_X1 U513 ( .A1(n533), .A2(n576), .ZN(n490) );
  NOR2_X1 U514 ( .A1(n530), .A2(n520), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n469), .A2(n460), .ZN(n461) );
  XOR2_X1 U516 ( .A(KEYINPUT25), .B(n461), .Z(n466) );
  XNOR2_X1 U517 ( .A(n520), .B(KEYINPUT94), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT27), .ZN(n470) );
  XOR2_X1 U519 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n464) );
  NAND2_X1 U520 ( .A1(n469), .A2(n530), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n464), .B(n463), .ZN(n570) );
  NOR2_X1 U522 ( .A1(n470), .A2(n570), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n474) );
  INV_X1 U525 ( .A(n532), .ZN(n472) );
  NOR2_X1 U526 ( .A1(n518), .A2(n470), .ZN(n528) );
  NAND2_X1 U527 ( .A1(n530), .A2(n528), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n487) );
  NOR2_X1 U530 ( .A1(n557), .A2(n540), .ZN(n475) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  NOR2_X1 U532 ( .A1(n487), .A2(n476), .ZN(n503) );
  NAND2_X1 U533 ( .A1(n490), .A2(n503), .ZN(n484) );
  NOR2_X1 U534 ( .A1(n518), .A2(n484), .ZN(n478) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(KEYINPUT96), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n479), .Z(G1324GAT) );
  NOR2_X1 U538 ( .A1(n520), .A2(n484), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(G1325GAT) );
  NOR2_X1 U541 ( .A1(n530), .A2(n484), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U544 ( .A1(n532), .A2(n484), .ZN(n485) );
  XOR2_X1 U545 ( .A(KEYINPUT98), .B(n485), .Z(n486) );
  XNOR2_X1 U546 ( .A(G22GAT), .B(n486), .ZN(G1327GAT) );
  NOR2_X1 U547 ( .A1(n586), .A2(n487), .ZN(n488) );
  NAND2_X1 U548 ( .A1(n540), .A2(n488), .ZN(n489) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n489), .ZN(n517) );
  NAND2_X1 U550 ( .A1(n517), .A2(n490), .ZN(n492) );
  XNOR2_X1 U551 ( .A(KEYINPUT100), .B(KEYINPUT38), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n500) );
  NOR2_X1 U553 ( .A1(n518), .A2(n500), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n520), .A2(n500), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT101), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1329GAT) );
  NOR2_X1 U559 ( .A1(n530), .A2(n500), .ZN(n498) );
  XNOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U562 ( .A(G43GAT), .B(n499), .Z(G1330GAT) );
  NOR2_X1 U563 ( .A1(n532), .A2(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(G1331GAT) );
  NOR2_X1 U566 ( .A1(n571), .A2(n535), .ZN(n516) );
  NAND2_X1 U567 ( .A1(n503), .A2(n516), .ZN(n504) );
  XOR2_X1 U568 ( .A(KEYINPUT105), .B(n504), .Z(n511) );
  NOR2_X1 U569 ( .A1(n518), .A2(n511), .ZN(n506) );
  XNOR2_X1 U570 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n507), .Z(G1332GAT) );
  NOR2_X1 U573 ( .A1(n520), .A2(n511), .ZN(n508) );
  XOR2_X1 U574 ( .A(G64GAT), .B(n508), .Z(G1333GAT) );
  NOR2_X1 U575 ( .A1(n530), .A2(n511), .ZN(n509) );
  XOR2_X1 U576 ( .A(KEYINPUT106), .B(n509), .Z(n510) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U578 ( .A1(n511), .A2(n532), .ZN(n515) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n513) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT108), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n523) );
  NOR2_X1 U584 ( .A1(n518), .A2(n523), .ZN(n519) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n519), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n520), .A2(n523), .ZN(n521) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U588 ( .A1(n530), .A2(n523), .ZN(n522) );
  XOR2_X1 U589 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  NOR2_X1 U590 ( .A1(n532), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NAND2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n547) );
  NOR2_X1 U595 ( .A1(n530), .A2(n547), .ZN(n531) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n543) );
  NOR2_X1 U597 ( .A1(n533), .A2(n543), .ZN(n534) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n534), .Z(G1340GAT) );
  NOR2_X1 U599 ( .A1(n535), .A2(n543), .ZN(n537) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n539) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n542) );
  NOR2_X1 U605 ( .A1(n540), .A2(n543), .ZN(n541) );
  XOR2_X1 U606 ( .A(n542), .B(n541), .Z(G1342GAT) );
  NOR2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U610 ( .A1(n570), .A2(n547), .ZN(n548) );
  XNOR2_X1 U611 ( .A(KEYINPUT114), .B(n548), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n558), .A2(n571), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n551) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U617 ( .A(KEYINPUT115), .B(n552), .Z(n554) );
  NAND2_X1 U618 ( .A1(n561), .A2(n558), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  XOR2_X1 U620 ( .A(G155GAT), .B(KEYINPUT117), .Z(n556) );
  NAND2_X1 U621 ( .A1(n558), .A2(n581), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n571), .A2(n566), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n566), .A2(n561), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  XOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT121), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n581), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT60), .Z(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n584) );
  NAND2_X1 U637 ( .A1(n584), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n578) );
  NAND2_X1 U642 ( .A1(n584), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n580) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT124), .Z(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  INV_X1 U649 ( .A(n584), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(G218GAT), .ZN(G1355GAT) );
endmodule

