

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601;

  XNOR2_X1 U324 ( .A(n364), .B(n363), .ZN(n365) );
  INV_X1 U325 ( .A(KEYINPUT48), .ZN(n412) );
  XNOR2_X1 U326 ( .A(n482), .B(n481), .ZN(n490) );
  XNOR2_X1 U327 ( .A(n480), .B(KEYINPUT37), .ZN(n481) );
  XNOR2_X1 U328 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U329 ( .A(n383), .B(n382), .ZN(n589) );
  AND2_X1 U330 ( .A1(n456), .A2(n455), .ZN(n571) );
  XNOR2_X1 U331 ( .A(n567), .B(n404), .ZN(n576) );
  XNOR2_X1 U332 ( .A(KEYINPUT90), .B(n466), .ZN(n580) );
  NOR2_X1 U333 ( .A1(n471), .A2(n348), .ZN(n292) );
  XOR2_X1 U334 ( .A(n392), .B(n391), .Z(n293) );
  XOR2_X1 U335 ( .A(n387), .B(n386), .Z(n294) );
  NOR2_X1 U336 ( .A1(n585), .A2(n408), .ZN(n409) );
  NOR2_X1 U337 ( .A1(n557), .A2(n433), .ZN(n434) );
  INV_X1 U338 ( .A(KEYINPUT101), .ZN(n480) );
  OR2_X1 U339 ( .A1(n411), .A2(n410), .ZN(n413) );
  XNOR2_X1 U340 ( .A(n362), .B(n370), .ZN(n363) );
  XNOR2_X1 U341 ( .A(n413), .B(n412), .ZN(n557) );
  XNOR2_X1 U342 ( .A(n427), .B(n426), .ZN(n430) );
  XNOR2_X1 U343 ( .A(n436), .B(n435), .ZN(n456) );
  XOR2_X1 U344 ( .A(KEYINPUT41), .B(n589), .Z(n545) );
  NOR2_X1 U345 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U346 ( .A1(n576), .A2(n575), .ZN(n578) );
  XOR2_X1 U347 ( .A(n398), .B(n397), .Z(n585) );
  XNOR2_X1 U348 ( .A(n432), .B(n431), .ZN(n533) );
  XNOR2_X1 U349 ( .A(n457), .B(G183GAT), .ZN(n458) );
  XNOR2_X1 U350 ( .A(n486), .B(KEYINPUT112), .ZN(n487) );
  XNOR2_X1 U351 ( .A(n459), .B(n458), .ZN(G1350GAT) );
  XNOR2_X1 U352 ( .A(n488), .B(n487), .ZN(G1338GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT15), .B(G64GAT), .Z(n296) );
  XNOR2_X1 U354 ( .A(G155GAT), .B(G57GAT), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n296), .B(n295), .ZN(n299) );
  XNOR2_X1 U356 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n297), .B(KEYINPUT12), .ZN(n298) );
  XOR2_X1 U358 ( .A(n299), .B(n298), .Z(n301) );
  NAND2_X1 U359 ( .A1(G231GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n307) );
  XNOR2_X1 U361 ( .A(G8GAT), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n302), .B(G211GAT), .ZN(n419) );
  XNOR2_X1 U363 ( .A(G71GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n303), .B(KEYINPUT13), .ZN(n380) );
  XOR2_X1 U365 ( .A(n419), .B(n380), .Z(n305) );
  XOR2_X1 U366 ( .A(G15GAT), .B(G22GAT), .Z(n387) );
  XOR2_X1 U367 ( .A(G1GAT), .B(G127GAT), .Z(n338) );
  XNOR2_X1 U368 ( .A(n387), .B(n338), .ZN(n304) );
  XNOR2_X1 U369 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n405) );
  INV_X1 U371 ( .A(n405), .ZN(n593) );
  XNOR2_X1 U372 ( .A(KEYINPUT113), .B(n593), .ZN(n549) );
  XOR2_X1 U373 ( .A(KEYINPUT24), .B(G148GAT), .Z(n309) );
  XNOR2_X1 U374 ( .A(G22GAT), .B(KEYINPUT70), .ZN(n308) );
  XNOR2_X1 U375 ( .A(n309), .B(n308), .ZN(n322) );
  XOR2_X1 U376 ( .A(G50GAT), .B(G162GAT), .Z(n361) );
  XOR2_X1 U377 ( .A(KEYINPUT22), .B(G78GAT), .Z(n311) );
  XNOR2_X1 U378 ( .A(G218GAT), .B(G106GAT), .ZN(n310) );
  XNOR2_X1 U379 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U380 ( .A(n361), .B(n312), .ZN(n314) );
  AND2_X1 U381 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U382 ( .A(n314), .B(n313), .ZN(n316) );
  INV_X1 U383 ( .A(G211GAT), .ZN(n315) );
  XNOR2_X1 U384 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U385 ( .A(G155GAT), .B(KEYINPUT2), .Z(n318) );
  XNOR2_X1 U386 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n317) );
  XNOR2_X1 U387 ( .A(n318), .B(n317), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n332), .B(KEYINPUT23), .ZN(n319) );
  XNOR2_X1 U389 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U390 ( .A(n322), .B(n321), .ZN(n327) );
  XNOR2_X1 U391 ( .A(KEYINPUT21), .B(KEYINPUT84), .ZN(n323) );
  XNOR2_X1 U392 ( .A(n323), .B(KEYINPUT85), .ZN(n324) );
  XNOR2_X1 U393 ( .A(n324), .B(KEYINPUT83), .ZN(n326) );
  XNOR2_X1 U394 ( .A(G197GAT), .B(G204GAT), .ZN(n325) );
  XNOR2_X1 U395 ( .A(n326), .B(n325), .ZN(n417) );
  XNOR2_X1 U396 ( .A(n327), .B(n417), .ZN(n471) );
  XOR2_X1 U397 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n329) );
  NAND2_X1 U398 ( .A1(G225GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U399 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U400 ( .A(n330), .B(KEYINPUT88), .Z(n334) );
  XNOR2_X1 U401 ( .A(G120GAT), .B(G148GAT), .ZN(n331) );
  XNOR2_X1 U402 ( .A(n331), .B(G57GAT), .ZN(n381) );
  XNOR2_X1 U403 ( .A(n332), .B(n381), .ZN(n333) );
  XNOR2_X1 U404 ( .A(n334), .B(n333), .ZN(n342) );
  XOR2_X1 U405 ( .A(KEYINPUT87), .B(KEYINPUT6), .Z(n336) );
  XNOR2_X1 U406 ( .A(KEYINPUT86), .B(KEYINPUT5), .ZN(n335) );
  XNOR2_X1 U407 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U408 ( .A(n337), .B(KEYINPUT1), .Z(n340) );
  XNOR2_X1 U409 ( .A(G162GAT), .B(n338), .ZN(n339) );
  XNOR2_X1 U410 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U411 ( .A(n342), .B(n341), .Z(n347) );
  XOR2_X1 U412 ( .A(KEYINPUT79), .B(KEYINPUT0), .Z(n344) );
  XNOR2_X1 U413 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n343) );
  XNOR2_X1 U414 ( .A(n344), .B(n343), .ZN(n446) );
  XNOR2_X1 U415 ( .A(G29GAT), .B(G134GAT), .ZN(n345) );
  XNOR2_X1 U416 ( .A(n345), .B(G85GAT), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n446), .B(n360), .ZN(n346) );
  XNOR2_X1 U418 ( .A(n347), .B(n346), .ZN(n466) );
  INV_X1 U419 ( .A(n580), .ZN(n348) );
  XOR2_X1 U420 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n350) );
  XNOR2_X1 U421 ( .A(KEYINPUT65), .B(KEYINPUT75), .ZN(n349) );
  XNOR2_X1 U422 ( .A(n350), .B(n349), .ZN(n366) );
  XOR2_X1 U423 ( .A(G43GAT), .B(KEYINPUT7), .Z(n352) );
  XNOR2_X1 U424 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n351) );
  XNOR2_X1 U425 ( .A(n352), .B(n351), .ZN(n386) );
  XOR2_X1 U426 ( .A(G92GAT), .B(G218GAT), .Z(n354) );
  XNOR2_X1 U427 ( .A(G36GAT), .B(G190GAT), .ZN(n353) );
  XNOR2_X1 U428 ( .A(n354), .B(n353), .ZN(n428) );
  XNOR2_X1 U429 ( .A(n386), .B(n428), .ZN(n359) );
  XOR2_X1 U430 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n356) );
  NAND2_X1 U431 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U432 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U433 ( .A(n357), .B(KEYINPUT11), .ZN(n358) );
  XNOR2_X1 U434 ( .A(n359), .B(n358), .ZN(n364) );
  XNOR2_X1 U435 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U436 ( .A(G99GAT), .B(G106GAT), .Z(n370) );
  XNOR2_X1 U437 ( .A(n366), .B(n365), .ZN(n567) );
  XOR2_X1 U438 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n368) );
  XNOR2_X1 U439 ( .A(KEYINPUT72), .B(KEYINPUT69), .ZN(n367) );
  XOR2_X1 U440 ( .A(n368), .B(n367), .Z(n373) );
  XOR2_X1 U441 ( .A(G176GAT), .B(G64GAT), .Z(n420) );
  XOR2_X1 U442 ( .A(G85GAT), .B(G92GAT), .Z(n369) );
  XNOR2_X1 U443 ( .A(n420), .B(n369), .ZN(n371) );
  XNOR2_X1 U444 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U445 ( .A(n373), .B(n372), .ZN(n375) );
  NAND2_X1 U446 ( .A1(G230GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U447 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U448 ( .A(KEYINPUT71), .B(KEYINPUT31), .Z(n377) );
  XNOR2_X1 U449 ( .A(G204GAT), .B(KEYINPUT70), .ZN(n376) );
  XOR2_X1 U450 ( .A(n377), .B(n376), .Z(n378) );
  XNOR2_X1 U451 ( .A(n379), .B(n378), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n381), .B(n380), .ZN(n382) );
  INV_X1 U453 ( .A(n545), .ZN(n570) );
  XOR2_X1 U454 ( .A(G197GAT), .B(G113GAT), .Z(n385) );
  XNOR2_X1 U455 ( .A(G169GAT), .B(G29GAT), .ZN(n384) );
  XNOR2_X1 U456 ( .A(n385), .B(n384), .ZN(n398) );
  XNOR2_X1 U457 ( .A(G36GAT), .B(G50GAT), .ZN(n388) );
  XNOR2_X1 U458 ( .A(n294), .B(n388), .ZN(n392) );
  XOR2_X1 U459 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n390) );
  NAND2_X1 U460 ( .A1(G229GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U461 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U462 ( .A(KEYINPUT66), .B(G8GAT), .Z(n394) );
  XNOR2_X1 U463 ( .A(G141GAT), .B(G1GAT), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U465 ( .A(n395), .B(KEYINPUT30), .ZN(n396) );
  XNOR2_X1 U466 ( .A(n293), .B(n396), .ZN(n397) );
  NAND2_X1 U467 ( .A1(n570), .A2(n585), .ZN(n400) );
  XNOR2_X1 U468 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n401) );
  NAND2_X1 U470 ( .A1(n401), .A2(n549), .ZN(n402) );
  NOR2_X1 U471 ( .A1(n567), .A2(n402), .ZN(n403) );
  XOR2_X1 U472 ( .A(KEYINPUT47), .B(n403), .Z(n411) );
  INV_X1 U473 ( .A(KEYINPUT76), .ZN(n404) );
  XNOR2_X1 U474 ( .A(KEYINPUT36), .B(n576), .ZN(n598) );
  NOR2_X1 U475 ( .A1(n598), .A2(n405), .ZN(n406) );
  XNOR2_X1 U476 ( .A(n406), .B(KEYINPUT45), .ZN(n407) );
  NAND2_X1 U477 ( .A1(n407), .A2(n589), .ZN(n408) );
  XOR2_X1 U478 ( .A(KEYINPUT115), .B(n409), .Z(n410) );
  XOR2_X1 U479 ( .A(KEYINPUT81), .B(KEYINPUT17), .Z(n415) );
  XNOR2_X1 U480 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U482 ( .A(G169GAT), .B(n416), .Z(n450) );
  XOR2_X1 U483 ( .A(n450), .B(n417), .Z(n432) );
  INV_X1 U484 ( .A(n420), .ZN(n418) );
  NAND2_X1 U485 ( .A1(n419), .A2(n418), .ZN(n423) );
  INV_X1 U486 ( .A(n419), .ZN(n421) );
  NAND2_X1 U487 ( .A1(n421), .A2(n420), .ZN(n422) );
  NAND2_X1 U488 ( .A1(n423), .A2(n422), .ZN(n427) );
  NAND2_X1 U489 ( .A1(G226GAT), .A2(G233GAT), .ZN(n425) );
  INV_X1 U490 ( .A(KEYINPUT91), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n428), .B(KEYINPUT92), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n533), .B(KEYINPUT120), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(KEYINPUT54), .ZN(n581) );
  AND2_X1 U495 ( .A1(n292), .A2(n581), .ZN(n436) );
  XNOR2_X1 U496 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n435) );
  XOR2_X1 U497 ( .A(KEYINPUT20), .B(G183GAT), .Z(n438) );
  XNOR2_X1 U498 ( .A(KEYINPUT82), .B(G127GAT), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n454) );
  XOR2_X1 U500 ( .A(G134GAT), .B(G99GAT), .Z(n440) );
  XNOR2_X1 U501 ( .A(G43GAT), .B(G190GAT), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U503 ( .A(KEYINPUT80), .B(G71GAT), .Z(n442) );
  XNOR2_X1 U504 ( .A(G15GAT), .B(G120GAT), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U506 ( .A(n444), .B(n443), .Z(n452) );
  INV_X1 U507 ( .A(G176GAT), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n448) );
  NAND2_X1 U509 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n454), .B(n453), .ZN(n540) );
  INV_X1 U514 ( .A(n540), .ZN(n455) );
  INV_X1 U515 ( .A(n571), .ZN(n575) );
  NOR2_X1 U516 ( .A1(n549), .A2(n575), .ZN(n459) );
  INV_X1 U517 ( .A(KEYINPUT122), .ZN(n457) );
  INV_X1 U518 ( .A(KEYINPUT110), .ZN(n485) );
  INV_X1 U519 ( .A(KEYINPUT100), .ZN(n478) );
  NAND2_X1 U520 ( .A1(n471), .A2(n540), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT26), .ZN(n582) );
  XOR2_X1 U522 ( .A(n533), .B(KEYINPUT93), .Z(n461) );
  XNOR2_X1 U523 ( .A(KEYINPUT27), .B(n461), .ZN(n470) );
  NOR2_X1 U524 ( .A1(n582), .A2(n470), .ZN(n559) );
  NOR2_X1 U525 ( .A1(n533), .A2(n540), .ZN(n462) );
  NOR2_X1 U526 ( .A1(n471), .A2(n462), .ZN(n463) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(n463), .Z(n464) );
  NOR2_X1 U528 ( .A1(n559), .A2(n464), .ZN(n465) );
  XNOR2_X1 U529 ( .A(n465), .B(KEYINPUT95), .ZN(n467) );
  NAND2_X1 U530 ( .A1(n467), .A2(n466), .ZN(n469) );
  INV_X1 U531 ( .A(KEYINPUT96), .ZN(n468) );
  XNOR2_X1 U532 ( .A(n469), .B(n468), .ZN(n476) );
  INV_X1 U533 ( .A(n470), .ZN(n472) );
  XOR2_X1 U534 ( .A(KEYINPUT28), .B(n471), .Z(n536) );
  NAND2_X1 U535 ( .A1(n472), .A2(n536), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n580), .A2(n473), .ZN(n542) );
  NAND2_X1 U537 ( .A1(n542), .A2(n540), .ZN(n474) );
  XOR2_X1 U538 ( .A(n474), .B(KEYINPUT94), .Z(n475) );
  NOR2_X2 U539 ( .A1(n476), .A2(n475), .ZN(n499) );
  NOR2_X1 U540 ( .A1(n593), .A2(n499), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n478), .B(n477), .ZN(n479) );
  NOR2_X1 U542 ( .A1(n598), .A2(n479), .ZN(n482) );
  INV_X1 U543 ( .A(n585), .ZN(n543) );
  NAND2_X1 U544 ( .A1(n570), .A2(n543), .ZN(n483) );
  XOR2_X1 U545 ( .A(KEYINPUT107), .B(n483), .Z(n520) );
  NOR2_X1 U546 ( .A1(n490), .A2(n520), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(n537) );
  NOR2_X1 U548 ( .A1(n537), .A2(n540), .ZN(n488) );
  INV_X1 U549 ( .A(G99GAT), .ZN(n486) );
  INV_X1 U550 ( .A(G50GAT), .ZN(n495) );
  NAND2_X1 U551 ( .A1(n589), .A2(n585), .ZN(n489) );
  XOR2_X1 U552 ( .A(KEYINPUT73), .B(n489), .Z(n496) );
  NOR2_X1 U553 ( .A1(n496), .A2(n490), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n514) );
  NOR2_X1 U556 ( .A1(n536), .A2(n514), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(KEYINPUT106), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(G1331GAT) );
  INV_X1 U559 ( .A(n496), .ZN(n500) );
  NAND2_X1 U560 ( .A1(n593), .A2(n576), .ZN(n497) );
  XNOR2_X1 U561 ( .A(KEYINPUT16), .B(n497), .ZN(n498) );
  NOR2_X1 U562 ( .A1(n499), .A2(n498), .ZN(n521) );
  NAND2_X1 U563 ( .A1(n500), .A2(n521), .ZN(n509) );
  NOR2_X1 U564 ( .A1(n580), .A2(n509), .ZN(n502) );
  XNOR2_X1 U565 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U567 ( .A(G1GAT), .B(n503), .ZN(G1324GAT) );
  NOR2_X1 U568 ( .A1(n533), .A2(n509), .ZN(n504) );
  XOR2_X1 U569 ( .A(KEYINPUT98), .B(n504), .Z(n505) );
  XNOR2_X1 U570 ( .A(G8GAT), .B(n505), .ZN(G1325GAT) );
  NOR2_X1 U571 ( .A1(n540), .A2(n509), .ZN(n507) );
  XNOR2_X1 U572 ( .A(KEYINPUT99), .B(KEYINPUT35), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U574 ( .A(G15GAT), .B(n508), .Z(G1326GAT) );
  NOR2_X1 U575 ( .A1(n536), .A2(n509), .ZN(n510) );
  XOR2_X1 U576 ( .A(G22GAT), .B(n510), .Z(G1327GAT) );
  NOR2_X1 U577 ( .A1(n580), .A2(n514), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1328GAT) );
  NOR2_X1 U580 ( .A1(n533), .A2(n514), .ZN(n513) );
  XOR2_X1 U581 ( .A(G36GAT), .B(n513), .Z(G1329GAT) );
  NOR2_X1 U582 ( .A1(n540), .A2(n514), .ZN(n519) );
  XOR2_X1 U583 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n516) );
  XNOR2_X1 U584 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n515) );
  XNOR2_X1 U585 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U586 ( .A(KEYINPUT103), .B(n517), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(G1330GAT) );
  INV_X1 U588 ( .A(n520), .ZN(n522) );
  NAND2_X1 U589 ( .A1(n522), .A2(n521), .ZN(n529) );
  NOR2_X1 U590 ( .A1(n580), .A2(n529), .ZN(n524) );
  XNOR2_X1 U591 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U593 ( .A(G57GAT), .B(n525), .Z(G1332GAT) );
  NOR2_X1 U594 ( .A1(n533), .A2(n529), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n527), .B(n526), .ZN(G1333GAT) );
  NOR2_X1 U597 ( .A1(n540), .A2(n529), .ZN(n528) );
  XOR2_X1 U598 ( .A(G71GAT), .B(n528), .Z(G1334GAT) );
  NOR2_X1 U599 ( .A1(n536), .A2(n529), .ZN(n531) );
  XNOR2_X1 U600 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n530) );
  XNOR2_X1 U601 ( .A(n531), .B(n530), .ZN(G1335GAT) );
  NOR2_X1 U602 ( .A1(n537), .A2(n580), .ZN(n532) );
  XOR2_X1 U603 ( .A(G85GAT), .B(n532), .Z(G1336GAT) );
  XNOR2_X1 U604 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n535) );
  NOR2_X1 U605 ( .A1(n533), .A2(n537), .ZN(n534) );
  XNOR2_X1 U606 ( .A(n535), .B(n534), .ZN(G1337GAT) );
  NOR2_X1 U607 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U608 ( .A(KEYINPUT44), .B(n538), .Z(n539) );
  XNOR2_X1 U609 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NOR2_X1 U610 ( .A1(n540), .A2(n557), .ZN(n541) );
  NAND2_X1 U611 ( .A1(n542), .A2(n541), .ZN(n552) );
  NOR2_X1 U612 ( .A1(n543), .A2(n552), .ZN(n544) );
  XOR2_X1 U613 ( .A(G113GAT), .B(n544), .Z(G1340GAT) );
  NOR2_X1 U614 ( .A1(n545), .A2(n552), .ZN(n547) );
  XNOR2_X1 U615 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U617 ( .A(G120GAT), .B(n548), .ZN(G1341GAT) );
  NOR2_X1 U618 ( .A1(n549), .A2(n552), .ZN(n550) );
  XOR2_X1 U619 ( .A(KEYINPUT50), .B(n550), .Z(n551) );
  XNOR2_X1 U620 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  NOR2_X1 U621 ( .A1(n552), .A2(n576), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n554) );
  XNOR2_X1 U623 ( .A(G134GAT), .B(KEYINPUT118), .ZN(n553) );
  XNOR2_X1 U624 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n556), .B(n555), .ZN(G1343GAT) );
  NOR2_X1 U626 ( .A1(n580), .A2(n557), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(KEYINPUT119), .B(n560), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n566), .A2(n585), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n561), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n563) );
  NAND2_X1 U632 ( .A1(n566), .A2(n570), .ZN(n562) );
  XNOR2_X1 U633 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U634 ( .A(G148GAT), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U635 ( .A1(n566), .A2(n593), .ZN(n565) );
  XNOR2_X1 U636 ( .A(n565), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U638 ( .A(n568), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U639 ( .A1(n585), .A2(n571), .ZN(n569) );
  XNOR2_X1 U640 ( .A(G169GAT), .B(n569), .ZN(G1348GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n573) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U643 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U644 ( .A(G176GAT), .B(n574), .ZN(G1349GAT) );
  XNOR2_X1 U645 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U647 ( .A(G190GAT), .B(n579), .ZN(G1351GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n587) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n583) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n584), .B(KEYINPUT124), .ZN(n592) );
  NAND2_X1 U652 ( .A1(n585), .A2(n592), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(G197GAT), .B(n588), .ZN(G1352GAT) );
  XOR2_X1 U655 ( .A(G204GAT), .B(KEYINPUT61), .Z(n591) );
  INV_X1 U656 ( .A(n592), .ZN(n597) );
  OR2_X1 U657 ( .A1(n597), .A2(n589), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n591), .B(n590), .ZN(G1353GAT) );
  XOR2_X1 U659 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n595) );
  NAND2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U662 ( .A(G211GAT), .B(n596), .ZN(G1354GAT) );
  XNOR2_X1 U663 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n600) );
  XNOR2_X1 U664 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U665 ( .A(G218GAT), .B(n601), .ZN(G1355GAT) );
endmodule

