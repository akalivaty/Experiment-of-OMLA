//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(new_n192), .ZN(new_n198));
  AND4_X1   g012(.A1(new_n196), .A2(new_n188), .A3(new_n190), .A4(new_n192), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT67), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n204), .A2(new_n207), .A3(new_n210), .A4(new_n205), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n213), .B(new_n195), .C1(new_n198), .C2(new_n199), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n201), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n203), .A2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n206), .A2(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n211), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  OR2_X1    g036(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n190), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(new_n188), .B2(new_n190), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n223), .A2(G128), .A3(new_n224), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(new_n197), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n220), .B(new_n222), .C1(new_n225), .C2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n215), .A2(KEYINPUT30), .A3(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(G116), .B(G119), .Z(new_n232));
  OR2_X1    g046(.A1(KEYINPUT2), .A2(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT2), .A2(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G116), .B(G119), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n233), .A3(new_n234), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(KEYINPUT66), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n240), .A3(new_n235), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n209), .A2(new_n211), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n228), .A2(new_n197), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n191), .A2(G128), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n225), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI22_X1  g060(.A1(new_n243), .A2(new_n200), .B1(new_n246), .B2(new_n219), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n242), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n231), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT31), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT27), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT26), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT27), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n253), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT26), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n255), .A2(new_n259), .A3(G101), .ZN(new_n260));
  AOI21_X1  g074(.A(G101), .B1(new_n255), .B2(new_n259), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n215), .A2(new_n242), .A3(new_n230), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n250), .A2(new_n251), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT70), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n263), .A2(new_n262), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n251), .A4(new_n250), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n231), .A2(new_n249), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n263), .A2(new_n262), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n266), .A2(KEYINPUT69), .A3(new_n250), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(KEYINPUT31), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n276));
  INV_X1    g090(.A(new_n242), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n247), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n263), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n262), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n263), .A2(new_n276), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT71), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n281), .B(new_n282), .C1(new_n279), .C2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n269), .A2(new_n275), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G472), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n269), .A2(new_n275), .A3(KEYINPUT72), .A4(new_n285), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n288), .A2(new_n289), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n286), .B2(new_n287), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n295), .A2(KEYINPUT32), .A3(new_n289), .A4(new_n291), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n250), .A2(new_n263), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT29), .B1(new_n298), .B2(new_n282), .ZN(new_n299));
  MUX2_X1   g113(.A(new_n284), .B(KEYINPUT71), .S(new_n279), .Z(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(new_n299), .C1(new_n300), .C2(new_n282), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n263), .A2(new_n278), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT71), .B(new_n283), .C1(new_n302), .C2(new_n276), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n282), .B1(new_n303), .B2(new_n281), .ZN(new_n304));
  INV_X1    g118(.A(new_n299), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT73), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n215), .A2(new_n230), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n277), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT74), .A3(new_n263), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n310), .A3(new_n277), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(KEYINPUT28), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n312), .A2(KEYINPUT29), .A3(new_n262), .A4(new_n283), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n301), .A2(new_n306), .A3(new_n290), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G472), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n294), .A2(new_n296), .A3(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT75), .B(G217), .Z(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G234), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(G902), .ZN(new_n320));
  XOR2_X1   g134(.A(G119), .B(G128), .Z(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT24), .B(G110), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(G128), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n226), .A2(KEYINPUT23), .A3(G119), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(G119), .C2(new_n226), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n323), .B1(G110), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT77), .B(G125), .ZN(new_n331));
  NOR2_X1   g145(.A1(KEYINPUT16), .A2(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT79), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT76), .A3(G125), .ZN(new_n339));
  AND3_X1   g153(.A1(KEYINPUT76), .A2(KEYINPUT77), .A3(G125), .ZN(new_n340));
  OAI21_X1  g154(.A(G140), .B1(KEYINPUT77), .B2(G125), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT16), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n337), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n187), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n337), .A2(new_n344), .A3(G146), .A4(new_n345), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n330), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  XOR2_X1   g163(.A(G125), .B(G140), .Z(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(G146), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n328), .A2(G110), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n321), .A2(new_n322), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G137), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT80), .ZN(new_n359));
  INV_X1    g173(.A(G953), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n360), .A2(G221), .A3(G234), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n359), .B(new_n361), .Z(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n349), .B2(new_n356), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n365), .A3(new_n290), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n320), .B1(new_n366), .B2(KEYINPUT25), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n365), .A3(new_n368), .A4(new_n290), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n320), .A2(new_n290), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n363), .A2(new_n365), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  OAI21_X1  g190(.A(G221), .B1(new_n376), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G469), .ZN(new_n379));
  XNOR2_X1  g193(.A(G110), .B(G140), .ZN(new_n380));
  INV_X1    g194(.A(G227), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G953), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n380), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G107), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(KEYINPUT81), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n386), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G101), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n385), .A2(G107), .ZN(new_n393));
  INV_X1    g207(.A(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G104), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(KEYINPUT81), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n391), .A2(new_n392), .A3(new_n393), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n392), .B1(new_n395), .B2(new_n393), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n189), .A2(KEYINPUT1), .A3(G146), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n398), .B(new_n400), .C1(new_n229), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT10), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n244), .A2(new_n245), .ZN(new_n404));
  INV_X1    g218(.A(new_n225), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n393), .B1(new_n386), .B2(new_n388), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n395), .B1(new_n396), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n399), .B1(new_n410), .B2(new_n392), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n402), .A2(new_n403), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n410), .B2(new_n392), .ZN(new_n414));
  OAI21_X1  g228(.A(G101), .B1(new_n407), .B2(new_n409), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT82), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n397), .B(new_n393), .C1(new_n417), .C2(new_n395), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(G101), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n413), .B(G101), .C1(new_n407), .C2(new_n409), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n201), .A2(new_n214), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n412), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT84), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n412), .B(new_n427), .C1(new_n422), .C2(new_n424), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n212), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n212), .B(KEYINPUT83), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n412), .B(new_n430), .C1(new_n422), .C2(new_n424), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n384), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n384), .ZN(new_n433));
  INV_X1    g247(.A(new_n246), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n402), .B1(new_n434), .B2(new_n411), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n435), .A2(KEYINPUT12), .A3(new_n212), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT12), .B1(new_n435), .B2(new_n212), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n379), .B(new_n290), .C1(new_n432), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n433), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n431), .B1(new_n436), .B2(new_n437), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n429), .A2(new_n441), .B1(new_n383), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G469), .B1(new_n443), .B2(G902), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n378), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G237), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n360), .A3(G214), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT89), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n189), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n252), .B(G214), .C1(KEYINPUT89), .C2(G143), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G131), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT91), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n454), .A3(G131), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT17), .ZN(new_n457));
  INV_X1    g271(.A(new_n451), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n210), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT17), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n453), .A2(new_n459), .A3(new_n460), .A4(new_n455), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n457), .A2(new_n347), .A3(new_n461), .A4(new_n348), .ZN(new_n462));
  XNOR2_X1  g276(.A(G113), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n385), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n451), .A2(KEYINPUT18), .A3(G131), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT90), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT18), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n458), .B1(new_n467), .B2(new_n210), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n340), .A2(new_n341), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n339), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G146), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(G146), .B2(new_n350), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n466), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n462), .A2(new_n464), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n464), .B1(new_n462), .B2(new_n473), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n290), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G475), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n453), .A2(new_n455), .A3(new_n459), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n350), .A2(KEYINPUT19), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n470), .B2(KEYINPUT19), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n479), .B(new_n348), .C1(G146), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n464), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n462), .A2(new_n473), .A3(new_n464), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(G475), .A2(G902), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n478), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n489), .ZN(new_n491));
  AOI211_X1 g305(.A(KEYINPUT20), .B(new_n491), .C1(new_n486), .C2(new_n487), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n477), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n317), .A2(G953), .A3(new_n376), .ZN(new_n494));
  XNOR2_X1  g308(.A(G128), .B(G143), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n203), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n495), .A2(KEYINPUT13), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n189), .A2(G128), .ZN(new_n498));
  OAI21_X1  g312(.A(G134), .B1(new_n498), .B2(KEYINPUT13), .ZN(new_n499));
  INV_X1    g313(.A(G122), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G116), .ZN(new_n501));
  INV_X1    g315(.A(G116), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G122), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G107), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n503), .A3(new_n394), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n505), .A2(KEYINPUT92), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT92), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  OAI221_X1 g322(.A(new_n496), .B1(new_n497), .B2(new_n499), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT93), .B1(new_n503), .B2(KEYINPUT14), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n503), .A2(KEYINPUT14), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n501), .A3(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n503), .A2(KEYINPUT93), .A3(KEYINPUT14), .ZN(new_n513));
  OAI21_X1  g327(.A(G107), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n496), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n495), .A2(new_n203), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n514), .B(new_n506), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n494), .B1(new_n509), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n509), .A2(new_n517), .A3(new_n494), .ZN(new_n520));
  AOI21_X1  g334(.A(G902), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n522));
  INV_X1    g336(.A(G478), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n521), .A2(new_n522), .B1(KEYINPUT15), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n525));
  INV_X1    g339(.A(new_n520), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(new_n518), .ZN(new_n527));
  OAI211_X1 g341(.A(KEYINPUT94), .B(new_n525), .C1(new_n527), .C2(G902), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n521), .A2(new_n522), .ZN(new_n529));
  NAND2_X1  g343(.A1(G234), .A2(G237), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(G952), .A3(new_n360), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT21), .B(G898), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(G902), .A3(G953), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n524), .A2(new_n528), .A3(new_n529), .A4(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n493), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n445), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT6), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n237), .A2(KEYINPUT5), .ZN(new_n540));
  INV_X1    g354(.A(G113), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n325), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n233), .A2(new_n234), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n540), .A2(new_n543), .B1(new_n544), .B2(new_n237), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n545), .A2(new_n398), .A3(new_n400), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n239), .A2(new_n423), .A3(new_n241), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n546), .B1(new_n421), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G122), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n539), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n549), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n239), .A2(new_n423), .A3(new_n241), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n419), .B1(new_n418), .B2(G101), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n552), .B1(new_n555), .B2(new_n420), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n551), .B1(new_n556), .B2(new_n546), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n200), .A2(new_n331), .ZN(new_n559));
  INV_X1    g373(.A(new_n331), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n246), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G224), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G953), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(KEYINPUT85), .Z(new_n565));
  XNOR2_X1  g379(.A(new_n562), .B(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n539), .B(new_n551), .C1(new_n556), .C2(new_n546), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n558), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT7), .B1(new_n563), .B2(G953), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT64), .B1(new_n191), .B2(new_n193), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n197), .A2(new_n196), .A3(new_n192), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n560), .B1(new_n572), .B2(new_n195), .ZN(new_n573));
  AOI211_X1 g387(.A(new_n331), .B(new_n225), .C1(new_n244), .C2(new_n245), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n569), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n559), .A2(new_n561), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n548), .B2(new_n549), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n549), .B(KEYINPUT8), .Z(new_n580));
  NAND2_X1  g394(.A1(new_n398), .A2(new_n400), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n545), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n542), .A2(new_n325), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G113), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n584), .A2(KEYINPUT86), .B1(new_n237), .B2(KEYINPUT5), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT86), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n543), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n585), .A2(new_n587), .B1(new_n544), .B2(new_n237), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n582), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT87), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n582), .B(KEYINPUT87), .C1(new_n581), .C2(new_n588), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n579), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n568), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(G210), .B1(G237), .B2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n568), .A2(new_n596), .A3(new_n594), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(KEYINPUT88), .A3(new_n599), .ZN(new_n600));
  AOI211_X1 g414(.A(KEYINPUT88), .B(new_n596), .C1(new_n568), .C2(new_n594), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G214), .B1(G237), .B2(G902), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n538), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n316), .A2(new_n375), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT95), .B(G101), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  INV_X1    g422(.A(new_n292), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT96), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n295), .A2(new_n612), .A3(new_n291), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(G472), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n611), .A2(KEYINPUT97), .A3(G472), .A4(new_n613), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n440), .A2(new_n444), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n377), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n374), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n603), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n598), .B2(new_n599), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n535), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n527), .B(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n290), .A2(G478), .ZN(new_n627));
  OAI22_X1  g441(.A1(new_n626), .A2(new_n627), .B1(G478), .B2(new_n521), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n493), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND3_X1  g447(.A1(new_n488), .A2(new_n478), .A3(new_n489), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT98), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n464), .B1(new_n473), .B2(new_n483), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n474), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT20), .B1(new_n637), .B2(new_n491), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n488), .A2(new_n639), .A3(new_n478), .A4(new_n489), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n635), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n477), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n625), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n622), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  OR2_X1    g461(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n357), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n372), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n370), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n605), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n616), .A2(new_n652), .A3(new_n617), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND2_X1  g469(.A1(new_n651), .A2(new_n624), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n534), .A2(G900), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(KEYINPUT99), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(KEYINPUT99), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n531), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n620), .A2(new_n643), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n316), .A2(new_n657), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT100), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n226), .ZN(G30));
  XNOR2_X1  g480(.A(new_n661), .B(KEYINPUT39), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n445), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT40), .Z(new_n669));
  AND2_X1   g483(.A1(new_n273), .A2(new_n274), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n309), .A2(new_n282), .A3(new_n311), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n672), .B2(G902), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n294), .A2(new_n296), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n600), .A2(new_n602), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT38), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n493), .A2(new_n642), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n678), .A2(new_n651), .A3(new_n623), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n669), .A2(new_n674), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  AND2_X1   g495(.A1(new_n493), .A2(new_n628), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n661), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n620), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n316), .A2(new_n657), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  OAI21_X1  g500(.A(new_n290), .B1(new_n432), .B2(new_n439), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n377), .A3(new_n440), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n316), .A2(new_n375), .A3(new_n690), .A4(new_n630), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n316), .A2(new_n375), .A3(new_n690), .A4(new_n644), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  NAND2_X1  g509(.A1(new_n537), .A2(new_n651), .ZN(new_n696));
  INV_X1    g510(.A(new_n599), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n596), .B1(new_n568), .B2(new_n594), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n603), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n696), .A2(new_n689), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n316), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  NOR3_X1   g516(.A1(new_n689), .A2(new_n625), .A3(new_n678), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n289), .A2(new_n290), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n269), .A2(new_n275), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n312), .A2(new_n283), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n282), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n704), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n610), .B2(G472), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n703), .A2(new_n375), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT101), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  INV_X1    g526(.A(new_n683), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n689), .A2(new_n699), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n709), .A3(new_n714), .A4(new_n651), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  XOR2_X1   g530(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n717));
  AOI21_X1  g531(.A(new_n623), .B1(new_n600), .B2(new_n602), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n718), .A2(KEYINPUT102), .A3(new_n445), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT102), .B1(new_n718), .B2(new_n445), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n713), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n316), .A2(new_n375), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n717), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n599), .A2(KEYINPUT88), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n698), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n603), .B1(new_n726), .B2(new_n601), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n724), .B1(new_n727), .B2(new_n620), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n718), .A2(KEYINPUT102), .A3(new_n445), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n683), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n316), .A4(new_n375), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n723), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  NOR2_X1   g547(.A1(new_n643), .A2(new_n662), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n719), .B2(new_n720), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n722), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n203), .ZN(G36));
  INV_X1    g551(.A(new_n493), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n628), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT43), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n741), .A3(new_n628), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n651), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n618), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT44), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n443), .A2(KEYINPUT45), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n443), .A2(KEYINPUT45), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(G469), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(G469), .A2(G902), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT104), .B1(new_n751), .B2(KEYINPUT46), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT46), .B1(new_n749), .B2(new_n750), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT104), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(KEYINPUT46), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n752), .A2(new_n440), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n377), .ZN(new_n758));
  INV_X1    g572(.A(new_n667), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n758), .A2(new_n759), .A3(new_n727), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n745), .A2(new_n746), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n757), .A2(new_n763), .A3(new_n377), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n763), .B1(new_n757), .B2(new_n377), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT105), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n316), .A2(new_n375), .A3(new_n683), .A4(new_n727), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n758), .A2(KEYINPUT47), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n764), .A3(new_n769), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT105), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NAND2_X1  g589(.A1(new_n690), .A2(new_n718), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT116), .ZN(new_n777));
  INV_X1    g591(.A(new_n674), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n374), .A2(new_n531), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n629), .ZN(new_n781));
  INV_X1    g595(.A(G952), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n781), .A2(new_n782), .A3(G953), .ZN(new_n783));
  INV_X1    g597(.A(new_n531), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n740), .A2(new_n784), .A3(new_n742), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n709), .A2(new_n375), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n714), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n783), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n722), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n793), .A3(new_n777), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT48), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n690), .A2(new_n623), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n677), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n677), .B2(new_n797), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n787), .A2(new_n798), .A3(new_n788), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT50), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n787), .A2(new_n651), .A3(new_n777), .A4(new_n709), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n493), .A2(new_n628), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n780), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT50), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n787), .A2(new_n788), .A3(new_n718), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n688), .A2(new_n440), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n378), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n809), .B1(new_n767), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT51), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n792), .B(new_n795), .C1(new_n808), .C2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n765), .B2(new_n766), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n771), .A2(KEYINPUT112), .A3(new_n764), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n811), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n809), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT113), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n822), .A3(new_n809), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n823), .A3(new_n807), .A4(new_n806), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n815), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n827));
  AND3_X1   g641(.A1(new_n616), .A2(new_n617), .A3(new_n652), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n691), .A2(new_n694), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n606), .A2(new_n701), .A3(new_n710), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n600), .A2(new_n602), .A3(new_n603), .A4(new_n535), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT108), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n682), .A2(new_n833), .B1(new_n738), .B2(new_n642), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n629), .A2(KEYINPUT108), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n616), .A2(new_n836), .A3(new_n617), .A4(new_n621), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n713), .B(new_n709), .C1(new_n719), .C2(new_n720), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n641), .A2(new_n477), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n642), .A2(new_n662), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n445), .A2(new_n718), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n316), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n651), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n736), .B1(new_n723), .B2(new_n731), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n831), .A2(new_n837), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n664), .A2(new_n715), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n678), .A2(new_n699), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n651), .A2(new_n662), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n849), .A2(new_n850), .A3(new_n445), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n674), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n847), .A2(new_n848), .A3(new_n685), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n664), .A2(new_n685), .A3(new_n715), .A4(new_n852), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n827), .B1(new_n846), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n858));
  INV_X1    g672(.A(new_n736), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n732), .A2(new_n859), .A3(new_n844), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n854), .B(new_n848), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n691), .A2(new_n694), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n606), .A2(new_n701), .A3(new_n710), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n653), .A2(new_n862), .A3(new_n863), .A4(new_n837), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n860), .A2(new_n861), .A3(new_n864), .A4(KEYINPUT53), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n857), .A2(new_n858), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n732), .A2(new_n859), .A3(new_n844), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n862), .A2(new_n863), .A3(new_n653), .A4(new_n837), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n856), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n827), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n846), .B2(new_n856), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n867), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n866), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n826), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(G952), .B2(G953), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n375), .A2(new_n603), .A3(new_n377), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT106), .ZN(new_n880));
  INV_X1    g694(.A(new_n739), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT49), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n880), .B(new_n881), .C1(new_n882), .C2(new_n810), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT107), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n677), .B1(new_n882), .B2(new_n810), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n778), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n878), .A2(new_n886), .ZN(G75));
  NOR2_X1   g701(.A1(new_n360), .A2(G952), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n889), .B(new_n290), .C1(new_n857), .C2(new_n865), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT120), .B1(new_n891), .B2(G902), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n597), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n558), .A2(new_n567), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n566), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT118), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(KEYINPUT56), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n888), .B1(new_n893), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n290), .B1(new_n857), .B2(new_n865), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(KEYINPUT119), .A3(G210), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT119), .B1(new_n900), .B2(G210), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n897), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n899), .A2(new_n905), .ZN(G51));
  INV_X1    g720(.A(new_n749), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n890), .B2(new_n892), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n432), .A2(new_n439), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n750), .B(KEYINPUT121), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT57), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n858), .B1(new_n857), .B2(new_n865), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n866), .B2(new_n913), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n908), .A2(new_n909), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(KEYINPUT122), .B(new_n907), .C1(new_n890), .C2(new_n892), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n888), .B1(new_n915), .B2(new_n916), .ZN(G54));
  AND2_X1   g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n890), .B2(new_n892), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n888), .B1(new_n919), .B2(new_n637), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n488), .B(new_n918), .C1(new_n890), .C2(new_n892), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(G60));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n923));
  INV_X1    g737(.A(new_n626), .ZN(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n858), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n891), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n857), .A2(new_n858), .A3(new_n865), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n923), .B1(new_n931), .B2(new_n888), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n926), .B1(new_n866), .B2(new_n875), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n626), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n931), .A2(new_n923), .A3(new_n888), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(G63));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n363), .A2(new_n365), .ZN(new_n939));
  INV_X1    g753(.A(new_n891), .ZN(new_n940));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n888), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n942), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n649), .B(KEYINPUT124), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n891), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n938), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n948), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n943), .A4(new_n944), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(G66));
  NAND3_X1  g766(.A1(new_n533), .A2(G224), .A3(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n869), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n894), .B1(G898), .B2(new_n360), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n954), .B(new_n955), .Z(G69));
  NOR2_X1   g770(.A1(new_n360), .A2(G900), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n381), .B2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT127), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n247), .A2(new_n248), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n231), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n482), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n680), .A2(new_n847), .A3(new_n685), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT62), .Z(new_n965));
  NAND3_X1  g779(.A1(new_n718), .A2(new_n445), .A3(new_n667), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n835), .B2(new_n834), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n793), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT125), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n965), .A2(new_n774), .A3(new_n761), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n963), .B1(new_n970), .B2(new_n360), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n793), .A2(new_n849), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n973), .A2(new_n758), .A3(new_n759), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n847), .A2(new_n685), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n774), .A2(new_n761), .A3(new_n845), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n957), .B1(new_n977), .B2(new_n360), .ZN(new_n978));
  INV_X1    g792(.A(new_n963), .ZN(new_n979));
  OAI22_X1  g793(.A1(new_n971), .A2(new_n972), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n971), .A2(new_n972), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n960), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n978), .A2(new_n979), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n970), .A2(new_n360), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT126), .B1(new_n985), .B2(new_n963), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n984), .A2(new_n986), .A3(new_n981), .A4(new_n959), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n983), .A2(new_n987), .ZN(G72));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n977), .B2(new_n869), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n298), .A2(new_n262), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n888), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n990), .B1(new_n970), .B2(new_n869), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n262), .A3(new_n298), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n872), .A2(new_n874), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n298), .A2(new_n282), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n670), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n996), .A2(new_n990), .A3(new_n998), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n993), .A2(new_n995), .A3(new_n999), .ZN(G57));
endmodule


