

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U558 ( .A1(n642), .A2(n548), .ZN(n662) );
  NOR2_X4 U559 ( .A1(n564), .A2(n563), .ZN(G160) );
  XOR2_X2 U560 ( .A(KEYINPUT17), .B(n531), .Z(n571) );
  NOR2_X1 U561 ( .A1(n723), .A2(n722), .ZN(n724) );
  BUF_X2 U562 ( .A(n556), .Z(n889) );
  AND2_X1 U563 ( .A1(n534), .A2(G2104), .ZN(n556) );
  NOR2_X2 U564 ( .A1(G2104), .A2(n534), .ZN(n895) );
  INV_X1 U565 ( .A(KEYINPUT101), .ZN(n718) );
  INV_X2 U566 ( .A(G2105), .ZN(n534) );
  XNOR2_X1 U567 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n557) );
  NOR2_X1 U568 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U569 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U570 ( .A1(n818), .A2(n826), .ZN(n526) );
  AND2_X1 U571 ( .A1(n526), .A2(n819), .ZN(n527) );
  OR2_X1 U572 ( .A1(n785), .A2(n784), .ZN(n528) );
  OR2_X1 U573 ( .A1(n771), .A2(n785), .ZN(n529) );
  NOR2_X1 U574 ( .A1(n785), .A2(n766), .ZN(n530) );
  NOR2_X1 U575 ( .A1(n710), .A2(n955), .ZN(n711) );
  AND2_X1 U576 ( .A1(n735), .A2(n745), .ZN(n736) );
  INV_X1 U577 ( .A(G168), .ZN(n737) );
  AND2_X1 U578 ( .A1(n738), .A2(n737), .ZN(n741) );
  NOR2_X1 U579 ( .A1(G1966), .A2(n785), .ZN(n733) );
  AND2_X1 U580 ( .A1(n751), .A2(n745), .ZN(n746) );
  INV_X1 U581 ( .A(KEYINPUT32), .ZN(n759) );
  XNOR2_X1 U582 ( .A(n760), .B(n759), .ZN(n761) );
  INV_X1 U583 ( .A(KEYINPUT64), .ZN(n768) );
  NAND2_X1 U584 ( .A1(n960), .A2(n529), .ZN(n772) );
  NAND2_X1 U585 ( .A1(n807), .A2(n697), .ZN(n752) );
  NAND2_X1 U586 ( .A1(G8), .A2(n752), .ZN(n785) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n642) );
  NOR2_X1 U588 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n549), .Z(n656) );
  XNOR2_X1 U590 ( .A(n558), .B(n557), .ZN(n560) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  INV_X1 U592 ( .A(KEYINPUT90), .ZN(n541) );
  NOR2_X2 U593 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  NAND2_X1 U594 ( .A1(n571), .A2(G138), .ZN(n533) );
  NAND2_X1 U595 ( .A1(G126), .A2(n895), .ZN(n532) );
  AND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n556), .A2(G102), .ZN(n535) );
  XNOR2_X1 U598 ( .A(KEYINPUT89), .B(n535), .ZN(n537) );
  AND2_X1 U599 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  AND2_X1 U600 ( .A1(n894), .A2(G114), .ZN(n536) );
  XNOR2_X2 U601 ( .A(n541), .B(n540), .ZN(G164) );
  XOR2_X1 U602 ( .A(KEYINPUT4), .B(KEYINPUT75), .Z(n543) );
  NOR2_X1 U603 ( .A1(G651), .A2(G543), .ZN(n660) );
  NAND2_X1 U604 ( .A1(G89), .A2(n660), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U606 ( .A(KEYINPUT74), .B(n544), .ZN(n546) );
  INV_X1 U607 ( .A(G651), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n662), .A2(G76), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT5), .ZN(n554) );
  NOR2_X1 U611 ( .A1(G543), .A2(n548), .ZN(n549) );
  NAND2_X1 U612 ( .A1(G63), .A2(n656), .ZN(n551) );
  NOR2_X2 U613 ( .A1(G651), .A2(n642), .ZN(n657) );
  NAND2_X1 U614 ( .A1(G51), .A2(n657), .ZN(n550) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U619 ( .A1(G101), .A2(n889), .ZN(n558) );
  NAND2_X1 U620 ( .A1(G113), .A2(n894), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G137), .A2(n571), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G125), .A2(n895), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U625 ( .A1(G85), .A2(n660), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G72), .A2(n662), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G60), .A2(n656), .ZN(n568) );
  NAND2_X1 U629 ( .A1(G47), .A2(n657), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n569) );
  OR2_X1 U631 ( .A1(n570), .A2(n569), .ZN(G290) );
  AND2_X1 U632 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U633 ( .A1(G111), .A2(n894), .ZN(n573) );
  BUF_X1 U634 ( .A(n571), .Z(n890) );
  NAND2_X1 U635 ( .A1(G135), .A2(n890), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n895), .A2(G123), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT18), .B(n574), .Z(n575) );
  NOR2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n889), .A2(G99), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n1007) );
  XNOR2_X1 U642 ( .A(G2096), .B(n1007), .ZN(n579) );
  OR2_X1 U643 ( .A1(G2100), .A2(n579), .ZN(G156) );
  INV_X1 U644 ( .A(G132), .ZN(G219) );
  INV_X1 U645 ( .A(G108), .ZN(G238) );
  NAND2_X1 U646 ( .A1(G64), .A2(n656), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G52), .A2(n657), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n588) );
  NAND2_X1 U649 ( .A1(n662), .A2(G77), .ZN(n582) );
  XNOR2_X1 U650 ( .A(KEYINPUT67), .B(n582), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n660), .A2(G90), .ZN(n583) );
  XOR2_X1 U652 ( .A(KEYINPUT66), .B(n583), .Z(n584) );
  NOR2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U654 ( .A(n586), .B(KEYINPUT9), .ZN(n587) );
  NOR2_X1 U655 ( .A1(n588), .A2(n587), .ZN(G171) );
  XOR2_X1 U656 ( .A(G168), .B(KEYINPUT8), .Z(n589) );
  XNOR2_X1 U657 ( .A(KEYINPUT76), .B(n589), .ZN(G286) );
  NAND2_X1 U658 ( .A1(G7), .A2(G661), .ZN(n590) );
  XNOR2_X1 U659 ( .A(n590), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U660 ( .A(G223), .B(KEYINPUT71), .ZN(n836) );
  NAND2_X1 U661 ( .A1(n836), .A2(G567), .ZN(n591) );
  XOR2_X1 U662 ( .A(KEYINPUT11), .B(n591), .Z(G234) );
  NAND2_X1 U663 ( .A1(n660), .A2(G81), .ZN(n592) );
  XNOR2_X1 U664 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U665 ( .A1(G68), .A2(n662), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U667 ( .A(KEYINPUT13), .B(n595), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G56), .A2(n656), .ZN(n596) );
  XOR2_X1 U669 ( .A(KEYINPUT14), .B(n596), .Z(n599) );
  NAND2_X1 U670 ( .A1(n657), .A2(G43), .ZN(n597) );
  XOR2_X1 U671 ( .A(KEYINPUT72), .B(n597), .Z(n598) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n955) );
  INV_X1 U673 ( .A(G860), .ZN(n630) );
  OR2_X1 U674 ( .A1(n955), .A2(n630), .ZN(G153) );
  INV_X1 U675 ( .A(G171), .ZN(G301) );
  NAND2_X1 U676 ( .A1(G868), .A2(G301), .ZN(n611) );
  NAND2_X1 U677 ( .A1(G92), .A2(n660), .ZN(n603) );
  NAND2_X1 U678 ( .A1(G66), .A2(n656), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G79), .A2(n662), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G54), .A2(n657), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U683 ( .A(KEYINPUT73), .B(n606), .Z(n607) );
  XNOR2_X2 U684 ( .A(KEYINPUT15), .B(n609), .ZN(n949) );
  INV_X1 U685 ( .A(G868), .ZN(n678) );
  NAND2_X1 U686 ( .A1(n949), .A2(n678), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(G284) );
  NAND2_X1 U688 ( .A1(G91), .A2(n660), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G78), .A2(n662), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U691 ( .A(KEYINPUT68), .B(n614), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G65), .A2(n656), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G53), .A2(n657), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n952) );
  XNOR2_X1 U696 ( .A(n952), .B(KEYINPUT69), .ZN(G299) );
  NOR2_X1 U697 ( .A1(G868), .A2(G299), .ZN(n619) );
  XOR2_X1 U698 ( .A(KEYINPUT77), .B(n619), .Z(n621) );
  NOR2_X1 U699 ( .A1(G286), .A2(n678), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(G297) );
  NAND2_X1 U701 ( .A1(n630), .A2(G559), .ZN(n622) );
  INV_X1 U702 ( .A(n949), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n622), .A2(n628), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n623), .B(KEYINPUT78), .ZN(n624) );
  XNOR2_X1 U705 ( .A(KEYINPUT16), .B(n624), .ZN(G148) );
  NOR2_X1 U706 ( .A1(G868), .A2(n955), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G868), .A2(n628), .ZN(n625) );
  NOR2_X1 U708 ( .A1(G559), .A2(n625), .ZN(n626) );
  NOR2_X1 U709 ( .A1(n627), .A2(n626), .ZN(G282) );
  NAND2_X1 U710 ( .A1(G559), .A2(n628), .ZN(n629) );
  XOR2_X1 U711 ( .A(n955), .B(n629), .Z(n675) );
  NAND2_X1 U712 ( .A1(n630), .A2(n675), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G93), .A2(n660), .ZN(n631) );
  XNOR2_X1 U714 ( .A(n631), .B(KEYINPUT79), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G80), .A2(n662), .ZN(n632) );
  XOR2_X1 U716 ( .A(KEYINPUT80), .B(n632), .Z(n633) );
  NOR2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n657), .A2(G55), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U720 ( .A1(G67), .A2(n656), .ZN(n637) );
  XNOR2_X1 U721 ( .A(KEYINPUT81), .B(n637), .ZN(n638) );
  NOR2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n677) );
  XOR2_X1 U723 ( .A(n640), .B(n677), .Z(G145) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n641) );
  XNOR2_X1 U725 ( .A(n641), .B(KEYINPUT82), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G49), .A2(n657), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G87), .A2(n642), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U729 ( .A1(n656), .A2(n645), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U731 ( .A1(n657), .A2(G48), .ZN(n654) );
  NAND2_X1 U732 ( .A1(G86), .A2(n660), .ZN(n649) );
  NAND2_X1 U733 ( .A1(G61), .A2(n656), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U735 ( .A1(n662), .A2(G73), .ZN(n650) );
  XOR2_X1 U736 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U737 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U738 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U739 ( .A(KEYINPUT83), .B(n655), .Z(G305) );
  NAND2_X1 U740 ( .A1(G62), .A2(n656), .ZN(n659) );
  NAND2_X1 U741 ( .A1(G50), .A2(n657), .ZN(n658) );
  NAND2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n660), .A2(G88), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n661), .B(KEYINPUT84), .ZN(n664) );
  NAND2_X1 U745 ( .A1(G75), .A2(n662), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U747 ( .A(KEYINPUT85), .B(n665), .Z(n666) );
  NOR2_X1 U748 ( .A1(n667), .A2(n666), .ZN(G166) );
  XNOR2_X1 U749 ( .A(KEYINPUT86), .B(KEYINPUT19), .ZN(n669) );
  XNOR2_X1 U750 ( .A(G288), .B(KEYINPUT87), .ZN(n668) );
  XNOR2_X1 U751 ( .A(n669), .B(n668), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n677), .B(G290), .ZN(n670) );
  XNOR2_X1 U753 ( .A(n670), .B(G299), .ZN(n671) );
  XNOR2_X1 U754 ( .A(n672), .B(n671), .ZN(n674) );
  XNOR2_X1 U755 ( .A(G305), .B(G166), .ZN(n673) );
  XNOR2_X1 U756 ( .A(n674), .B(n673), .ZN(n908) );
  XOR2_X1 U757 ( .A(n908), .B(n675), .Z(n676) );
  NOR2_X1 U758 ( .A1(n678), .A2(n676), .ZN(n680) );
  AND2_X1 U759 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U760 ( .A1(n680), .A2(n679), .ZN(G295) );
  NAND2_X1 U761 ( .A1(G2084), .A2(G2078), .ZN(n681) );
  XOR2_X1 U762 ( .A(KEYINPUT20), .B(n681), .Z(n682) );
  NAND2_X1 U763 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U764 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U766 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U767 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NAND2_X1 U768 ( .A1(G120), .A2(G69), .ZN(n685) );
  XNOR2_X1 U769 ( .A(KEYINPUT88), .B(n685), .ZN(n686) );
  NOR2_X1 U770 ( .A1(G238), .A2(n686), .ZN(n687) );
  NAND2_X1 U771 ( .A1(G57), .A2(n687), .ZN(n840) );
  NAND2_X1 U772 ( .A1(n840), .A2(G567), .ZN(n692) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n688) );
  XOR2_X1 U774 ( .A(KEYINPUT22), .B(n688), .Z(n689) );
  NOR2_X1 U775 ( .A1(G218), .A2(n689), .ZN(n690) );
  NAND2_X1 U776 ( .A1(G96), .A2(n690), .ZN(n841) );
  NAND2_X1 U777 ( .A1(n841), .A2(G2106), .ZN(n691) );
  NAND2_X1 U778 ( .A1(n692), .A2(n691), .ZN(n842) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n693) );
  NOR2_X1 U780 ( .A1(n842), .A2(n693), .ZN(n839) );
  NAND2_X1 U781 ( .A1(n839), .A2(G36), .ZN(G176) );
  XNOR2_X1 U782 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  NOR2_X2 U783 ( .A1(G1384), .A2(G164), .ZN(n807) );
  NAND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n806) );
  INV_X1 U785 ( .A(n806), .ZN(n697) );
  AND2_X2 U786 ( .A1(n807), .A2(n697), .ZN(n725) );
  NAND2_X1 U787 ( .A1(n725), .A2(G2072), .ZN(n694) );
  XNOR2_X1 U788 ( .A(n694), .B(KEYINPUT27), .ZN(n696) );
  INV_X1 U789 ( .A(G1956), .ZN(n976) );
  NOR2_X1 U790 ( .A1(n976), .A2(n725), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n720) );
  NAND2_X1 U792 ( .A1(n720), .A2(n952), .ZN(n714) );
  NAND2_X1 U793 ( .A1(G1348), .A2(n752), .ZN(n699) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n725), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n715) );
  NAND2_X1 U796 ( .A1(n715), .A2(n949), .ZN(n712) );
  INV_X1 U797 ( .A(KEYINPUT99), .ZN(n701) );
  NAND2_X1 U798 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n700) );
  AND2_X1 U799 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U800 ( .A1(n725), .A2(n702), .ZN(n706) );
  XNOR2_X1 U801 ( .A(KEYINPUT99), .B(G1341), .ZN(n703) );
  AND2_X1 U802 ( .A1(n703), .A2(KEYINPUT26), .ZN(n704) );
  NAND2_X1 U803 ( .A1(n752), .A2(n704), .ZN(n705) );
  NAND2_X1 U804 ( .A1(n706), .A2(n705), .ZN(n708) );
  OR2_X1 U805 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n707) );
  NAND2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U807 ( .A(KEYINPUT100), .B(n709), .ZN(n710) );
  NAND2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n717) );
  NOR2_X1 U810 ( .A1(n949), .A2(n715), .ZN(n716) );
  NOR2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U812 ( .A(n719), .B(n718), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n952), .A2(n720), .ZN(n721) );
  XNOR2_X1 U814 ( .A(KEYINPUT28), .B(n721), .ZN(n722) );
  XNOR2_X1 U815 ( .A(n724), .B(KEYINPUT29), .ZN(n729) );
  OR2_X1 U816 ( .A1(n725), .A2(G1961), .ZN(n727) );
  XNOR2_X1 U817 ( .A(G2078), .B(KEYINPUT25), .ZN(n930) );
  NAND2_X1 U818 ( .A1(n725), .A2(n930), .ZN(n726) );
  NAND2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n739) );
  NAND2_X1 U820 ( .A1(n739), .A2(G171), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n744) );
  INV_X1 U822 ( .A(G8), .ZN(n732) );
  INV_X1 U823 ( .A(KEYINPUT97), .ZN(n731) );
  NOR2_X1 U824 ( .A1(G2084), .A2(n752), .ZN(n730) );
  XNOR2_X1 U825 ( .A(n731), .B(n730), .ZN(n747) );
  NOR2_X1 U826 ( .A1(n732), .A2(n747), .ZN(n735) );
  INV_X1 U827 ( .A(KEYINPUT98), .ZN(n734) );
  XNOR2_X1 U828 ( .A(n734), .B(n733), .ZN(n745) );
  XNOR2_X1 U829 ( .A(n736), .B(KEYINPUT30), .ZN(n738) );
  NOR2_X1 U830 ( .A1(G171), .A2(n739), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U832 ( .A(KEYINPUT31), .B(n742), .Z(n743) );
  NAND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n751) );
  XNOR2_X1 U834 ( .A(n746), .B(KEYINPUT102), .ZN(n749) );
  NAND2_X1 U835 ( .A1(n747), .A2(G8), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n762) );
  AND2_X1 U837 ( .A1(G286), .A2(G8), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n758) );
  NOR2_X1 U839 ( .A1(G1971), .A2(n785), .ZN(n754) );
  NOR2_X1 U840 ( .A1(G2090), .A2(n752), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n755), .A2(G303), .ZN(n756) );
  OR2_X1 U843 ( .A1(n732), .A2(n756), .ZN(n757) );
  NAND2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n760) );
  NAND2_X1 U845 ( .A1(n762), .A2(n761), .ZN(n777) );
  NOR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n967) );
  NOR2_X1 U848 ( .A1(n965), .A2(n967), .ZN(n763) );
  XOR2_X1 U849 ( .A(KEYINPUT103), .B(n763), .Z(n764) );
  NAND2_X1 U850 ( .A1(n777), .A2(n764), .ZN(n765) );
  XNOR2_X1 U851 ( .A(n765), .B(KEYINPUT104), .ZN(n767) );
  NAND2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n968) );
  INV_X1 U853 ( .A(n968), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n767), .A2(n530), .ZN(n769) );
  XNOR2_X1 U855 ( .A(n769), .B(n768), .ZN(n770) );
  NOR2_X1 U856 ( .A1(KEYINPUT33), .A2(n770), .ZN(n773) );
  XOR2_X1 U857 ( .A(G1981), .B(G305), .Z(n960) );
  NAND2_X1 U858 ( .A1(n965), .A2(KEYINPUT33), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U860 ( .A(n774), .B(KEYINPUT105), .ZN(n781) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n775) );
  XNOR2_X1 U862 ( .A(KEYINPUT106), .B(n775), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n776), .A2(G8), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n779), .A2(n785), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U867 ( .A(n782), .B(KEYINPUT107), .ZN(n786) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n783) );
  XOR2_X1 U869 ( .A(n783), .B(KEYINPUT24), .Z(n784) );
  NAND2_X1 U870 ( .A1(n786), .A2(n528), .ZN(n820) );
  NAND2_X1 U871 ( .A1(G107), .A2(n894), .ZN(n788) );
  NAND2_X1 U872 ( .A1(G131), .A2(n890), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G95), .A2(n889), .ZN(n790) );
  NAND2_X1 U875 ( .A1(G119), .A2(n895), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U878 ( .A(KEYINPUT92), .B(n793), .Z(n881) );
  NAND2_X1 U879 ( .A1(G1991), .A2(n881), .ZN(n805) );
  NAND2_X1 U880 ( .A1(G105), .A2(n889), .ZN(n794) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(n794), .Z(n801) );
  NAND2_X1 U882 ( .A1(n895), .A2(G129), .ZN(n795) );
  XNOR2_X1 U883 ( .A(KEYINPUT93), .B(n795), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n894), .A2(G117), .ZN(n796) );
  XOR2_X1 U885 ( .A(KEYINPUT94), .B(n796), .Z(n797) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U887 ( .A(n799), .B(KEYINPUT95), .ZN(n800) );
  NOR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n890), .A2(G141), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n883) );
  NAND2_X1 U891 ( .A1(G1996), .A2(n883), .ZN(n804) );
  NAND2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n1005) );
  NOR2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n830) );
  NAND2_X1 U894 ( .A1(n1005), .A2(n830), .ZN(n808) );
  XOR2_X1 U895 ( .A(KEYINPUT96), .B(n808), .Z(n823) );
  INV_X1 U896 ( .A(n823), .ZN(n818) );
  NAND2_X1 U897 ( .A1(G104), .A2(n889), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G140), .A2(n890), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U900 ( .A(KEYINPUT34), .B(n811), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G116), .A2(n894), .ZN(n813) );
  NAND2_X1 U902 ( .A1(G128), .A2(n895), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U904 ( .A(KEYINPUT35), .B(n814), .Z(n815) );
  NOR2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U906 ( .A(KEYINPUT36), .B(n817), .ZN(n886) );
  XNOR2_X1 U907 ( .A(KEYINPUT37), .B(G2067), .ZN(n828) );
  NOR2_X1 U908 ( .A1(n886), .A2(n828), .ZN(n1013) );
  NAND2_X1 U909 ( .A1(n830), .A2(n1013), .ZN(n826) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n971) );
  NAND2_X1 U911 ( .A1(n971), .A2(n830), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n820), .A2(n527), .ZN(n833) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n883), .ZN(n1021) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n881), .A2(G1991), .ZN(n1010) );
  NOR2_X1 U916 ( .A1(n821), .A2(n1010), .ZN(n822) );
  NOR2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U918 ( .A1(n1021), .A2(n824), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n886), .A2(n828), .ZN(n1004) );
  NAND2_X1 U922 ( .A1(n829), .A2(n1004), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(n835) );
  XNOR2_X1 U925 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n834) );
  XNOR2_X1 U926 ( .A(n835), .B(n834), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U929 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U931 ( .A1(n839), .A2(n838), .ZN(G188) );
  XOR2_X1 U932 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  NOR2_X1 U936 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  INV_X1 U938 ( .A(n842), .ZN(G319) );
  XNOR2_X1 U939 ( .A(G1991), .B(KEYINPUT114), .ZN(n852) );
  XOR2_X1 U940 ( .A(G1976), .B(G1956), .Z(n844) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1986), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U943 ( .A(G1971), .B(G1961), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1981), .B(G1966), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2474), .B(KEYINPUT41), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G229) );
  XNOR2_X1 U950 ( .A(G2084), .B(G2090), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n853), .B(G2678), .ZN(n863) );
  XOR2_X1 U952 ( .A(KEYINPUT42), .B(KEYINPUT111), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT43), .B(G2096), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U955 ( .A(G2100), .B(G2072), .Z(n857) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2078), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U959 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(G227) );
  NAND2_X1 U962 ( .A1(G124), .A2(n895), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U964 ( .A1(n894), .A2(G112), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U966 ( .A1(G100), .A2(n889), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G136), .A2(n890), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U969 ( .A1(n870), .A2(n869), .ZN(G162) );
  XNOR2_X1 U970 ( .A(KEYINPUT48), .B(G164), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n871), .B(n1007), .ZN(n885) );
  XNOR2_X1 U972 ( .A(KEYINPUT47), .B(KEYINPUT117), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G115), .A2(n894), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G127), .A2(n895), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n880) );
  NAND2_X1 U977 ( .A1(n889), .A2(G103), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT116), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G139), .A2(n890), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n1016) );
  XOR2_X1 U982 ( .A(n881), .B(n1016), .Z(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n886), .B(KEYINPUT46), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n904) );
  NAND2_X1 U987 ( .A1(G106), .A2(n889), .ZN(n892) );
  NAND2_X1 U988 ( .A1(G142), .A2(n890), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n893), .B(KEYINPUT45), .ZN(n900) );
  NAND2_X1 U991 ( .A1(G118), .A2(n894), .ZN(n897) );
  NAND2_X1 U992 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(KEYINPUT115), .B(n898), .ZN(n899) );
  NAND2_X1 U995 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n901), .B(G162), .ZN(n902) );
  XOR2_X1 U997 ( .A(G160), .B(n902), .Z(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U999 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(G171), .B(n949), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n906), .B(G286), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(KEYINPUT118), .B(n907), .ZN(n910) );
  XNOR2_X1 U1003 ( .A(n955), .B(n908), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n911), .ZN(G397) );
  XOR2_X1 U1006 ( .A(G2430), .B(G2451), .Z(n913) );
  XNOR2_X1 U1007 ( .A(G2446), .B(G2427), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n920) );
  XOR2_X1 U1009 ( .A(G2438), .B(KEYINPUT109), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G2443), .B(G2454), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1012 ( .A(n916), .B(G2435), .Z(n918) );
  XNOR2_X1 U1013 ( .A(G1348), .B(G1341), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n920), .B(n919), .ZN(n921) );
  NAND2_X1 U1016 ( .A1(n921), .A2(G14), .ZN(n927) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G57), .ZN(G237) );
  INV_X1 U1025 ( .A(n927), .ZN(G401) );
  XNOR2_X1 U1026 ( .A(G2067), .B(G26), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(G32), .B(G1996), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n934) );
  XOR2_X1 U1029 ( .A(n930), .B(G27), .Z(n932) );
  XNOR2_X1 U1030 ( .A(G2072), .B(G33), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n938) );
  XOR2_X1 U1033 ( .A(G1991), .B(G25), .Z(n935) );
  NAND2_X1 U1034 ( .A1(n935), .A2(G28), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(KEYINPUT120), .B(n936), .ZN(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1037 ( .A(KEYINPUT53), .B(n939), .Z(n942) );
  XOR2_X1 U1038 ( .A(G34), .B(KEYINPUT54), .Z(n940) );
  XNOR2_X1 U1039 ( .A(G2084), .B(n940), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G35), .B(G2090), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n945), .A2(KEYINPUT55), .ZN(n1036) );
  INV_X1 U1044 ( .A(n945), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(G29), .A2(KEYINPUT55), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(G11), .A2(n948), .ZN(n1034) );
  XNOR2_X1 U1048 ( .A(KEYINPUT56), .B(G16), .ZN(n975) );
  XNOR2_X1 U1049 ( .A(G301), .B(G1961), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(n949), .B(G1348), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n952), .B(G1956), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(G1971), .A2(G303), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(G1341), .B(n955), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1060 ( .A(KEYINPUT57), .B(n962), .Z(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n973) );
  XOR2_X1 U1062 ( .A(n965), .B(KEYINPUT121), .Z(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n1002) );
  XNOR2_X1 U1068 ( .A(G20), .B(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(G1341), .B(G19), .Z(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(G6), .B(G1981), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1073 ( .A(KEYINPUT122), .B(n981), .Z(n985) );
  XNOR2_X1 U1074 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(G4), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(G1348), .B(n983), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(KEYINPUT60), .B(n986), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G21), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(G1961), .B(G5), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(G1971), .B(G22), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(G23), .B(G1976), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n994) );
  XOR2_X1 U1086 ( .A(G1986), .B(G24), .Z(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(KEYINPUT58), .B(n995), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1090 ( .A(KEYINPUT61), .B(n998), .Z(n999) );
  NOR2_X1 U1091 ( .A1(G16), .A2(n999), .ZN(n1000) );
  XOR2_X1 U1092 ( .A(KEYINPUT124), .B(n1000), .Z(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(n1003), .B(KEYINPUT125), .ZN(n1032) );
  INV_X1 U1095 ( .A(n1004), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1015) );
  XNOR2_X1 U1097 ( .A(G160), .B(G2084), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT119), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1026) );
  XOR2_X1 U1103 ( .A(G2072), .B(n1016), .Z(n1018) );
  XOR2_X1 U1104 ( .A(G164), .B(G2078), .Z(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT50), .B(n1019), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(G2090), .B(G162), .Z(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(KEYINPUT51), .B(n1022), .Z(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(KEYINPUT52), .B(n1027), .ZN(n1029) );
  INV_X1 U1113 ( .A(KEYINPUT55), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(G29), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1119 ( .A(n1037), .B(KEYINPUT62), .ZN(n1038) );
  XOR2_X1 U1120 ( .A(KEYINPUT126), .B(n1038), .Z(G311) );
  XNOR2_X1 U1121 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

