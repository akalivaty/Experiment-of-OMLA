//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n595, new_n596,
    new_n597, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n467), .B1(new_n470), .B2(G137), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n464), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n471), .B1(new_n476), .B2(KEYINPUT66), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n478));
  AOI211_X1 g053(.A(new_n478), .B(new_n464), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT67), .Z(G160));
  NAND2_X1  g056(.A1(new_n470), .A2(G136), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n472), .B2(new_n473), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(KEYINPUT68), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n464), .A2(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n468), .B2(new_n469), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n490), .B(new_n501), .C1(new_n473), .C2(new_n472), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n493), .B(new_n498), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT69), .A3(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT69), .A2(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n510), .A2(G50), .A3(new_n514), .A4(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT6), .B1(KEYINPUT69), .B2(G651), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n520), .A2(KEYINPUT71), .A3(G50), .A4(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT69), .B(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n523), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n531), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n510), .A2(G88), .A3(new_n514), .A4(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n522), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(G166));
  NAND2_X1  g113(.A1(new_n520), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n510), .A2(new_n514), .A3(new_n534), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G89), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n547));
  AND2_X1   g122(.A1(G63), .A2(G651), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n546), .A2(new_n547), .B1(new_n534), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n541), .A2(new_n544), .A3(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  NAND2_X1  g126(.A1(new_n540), .A2(G52), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n543), .A2(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n534), .ZN(new_n555));
  INV_X1    g130(.A(G64), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(new_n523), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n552), .A2(new_n553), .A3(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n555), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(G81), .A2(new_n543), .B1(new_n563), .B2(new_n523), .ZN(new_n564));
  INV_X1    g139(.A(G43), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n565), .B2(new_n539), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g146(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n572));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  NAND3_X1  g150(.A1(new_n520), .A2(G53), .A3(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n543), .A2(G91), .ZN(new_n578));
  AND2_X1   g153(.A1(KEYINPUT5), .A2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(KEYINPUT5), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT75), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n530), .A2(new_n582), .A3(new_n531), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G65), .ZN(new_n585));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT76), .B1(new_n587), .B2(G651), .ZN(new_n588));
  INV_X1    g163(.A(G65), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n581), .B2(new_n583), .ZN(new_n590));
  INV_X1    g165(.A(new_n586), .ZN(new_n591));
  OAI211_X1 g166(.A(KEYINPUT76), .B(G651), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n577), .B(new_n578), .C1(new_n588), .C2(new_n593), .ZN(G299));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n537), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n522), .A2(new_n536), .A3(KEYINPUT77), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(G303));
  NAND3_X1  g173(.A1(new_n520), .A2(G87), .A3(new_n534), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n600));
  INV_X1    g175(.A(G49), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n539), .C2(new_n601), .ZN(G288));
  INV_X1    g177(.A(G61), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n530), .B2(new_n531), .ZN(new_n604));
  AND2_X1   g179(.A1(G73), .A2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n523), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n510), .A2(G48), .A3(new_n514), .A4(G543), .ZN(new_n607));
  INV_X1    g182(.A(G86), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(new_n542), .C2(new_n608), .ZN(G305));
  AOI22_X1  g184(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(KEYINPUT78), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(KEYINPUT78), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n611), .A2(new_n523), .A3(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n540), .A2(G47), .B1(new_n543), .B2(G85), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT79), .Z(new_n617));
  NAND2_X1  g192(.A1(new_n543), .A2(G92), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT10), .Z(new_n619));
  INV_X1    g194(.A(G54), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n620), .B1(new_n539), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(new_n539), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n584), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(new_n511), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n619), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n617), .B1(G868), .B2(new_n627), .ZN(G284));
  OAI21_X1  g203(.A(new_n617), .B1(G868), .B2(new_n627), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n627), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n627), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n483), .A2(G123), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT81), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(G111), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(G2105), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(G135), .B2(new_n470), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n651), .A2(G2100), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(G2100), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n646), .A2(G2096), .ZN(new_n654));
  NAND4_X1  g229(.A1(new_n647), .A2(new_n652), .A3(new_n653), .A4(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT82), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2430), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XOR2_X1   g239(.A(G1341), .B(G1348), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2443), .B(G2446), .Z(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT84), .Z(new_n674));
  XOR2_X1   g249(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2084), .B(G2090), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n674), .B2(new_n677), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n676), .B2(new_n677), .ZN(new_n681));
  INV_X1    g256(.A(new_n677), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n682), .A2(new_n678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n679), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT20), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n691), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n691), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(G229));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NOR2_X1   g283(.A1(G168), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n708), .B2(G21), .ZN(new_n710));
  INV_X1    g285(.A(G1966), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(G5), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G171), .B2(new_n708), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n710), .A2(new_n711), .B1(new_n714), .B2(G1961), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n641), .A2(G29), .A3(new_n645), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(KEYINPUT93), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(KEYINPUT93), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT31), .B(G11), .Z(new_n719));
  XOR2_X1   g294(.A(KEYINPUT30), .B(G28), .Z(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(G29), .ZN(new_n721));
  NOR4_X1   g296(.A1(new_n717), .A2(new_n718), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n712), .A2(new_n715), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n726), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT29), .Z(new_n729));
  INV_X1    g304(.A(G2090), .ZN(new_n730));
  OAI22_X1  g305(.A1(new_n729), .A2(new_n730), .B1(G1961), .B2(new_n714), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(new_n729), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n726), .A2(G32), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n470), .A2(G141), .ZN(new_n734));
  INV_X1    g309(.A(G105), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n465), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT26), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n483), .A2(G129), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n733), .B1(new_n742), .B2(new_n726), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT27), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1996), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT25), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n470), .A2(G139), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT3), .B(G2104), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n749), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n748), .C1(new_n750), .C2(new_n464), .ZN(new_n751));
  MUX2_X1   g326(.A(G33), .B(new_n751), .S(G29), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2072), .ZN(new_n753));
  NOR2_X1   g328(.A1(G27), .A2(G29), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G164), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2078), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n726), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT90), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n470), .A2(G140), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n483), .A2(G128), .ZN(new_n761));
  OR2_X1    g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n763));
  AND3_X1   g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n759), .B1(new_n726), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2067), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n753), .A2(new_n756), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n725), .A2(new_n732), .A3(new_n745), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(G160), .A2(G29), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n770), .B2(G34), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G34), .B2(new_n770), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT92), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2084), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n723), .B2(new_n724), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n768), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n708), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n631), .B2(new_n708), .ZN(new_n780));
  INV_X1    g355(.A(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n708), .A2(G19), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n569), .B2(new_n708), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1341), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n708), .A2(G4), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n627), .B2(new_n708), .ZN(new_n787));
  INV_X1    g362(.A(G1348), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n777), .A2(new_n782), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT34), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n708), .A2(G22), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n537), .B2(G16), .ZN(new_n793));
  INV_X1    g368(.A(G1971), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT88), .ZN(new_n796));
  MUX2_X1   g371(.A(G6), .B(G305), .S(G16), .Z(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT32), .B(G1981), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n708), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(G288), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n708), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT33), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT33), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G1976), .ZN(new_n806));
  INV_X1    g381(.A(G1976), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n803), .A2(new_n807), .A3(new_n804), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n799), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n796), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n810), .A2(KEYINPUT89), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(KEYINPUT89), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n791), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n810), .A2(KEYINPUT89), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(KEYINPUT89), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n814), .A2(KEYINPUT34), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n726), .A2(G25), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G107), .B2(new_n464), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT87), .ZN(new_n821));
  AOI22_X1  g396(.A1(G119), .A2(new_n483), .B1(new_n470), .B2(G131), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n817), .B1(new_n823), .B2(new_n726), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G1986), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n708), .A2(G24), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G290), .B2(G16), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n813), .A2(new_n816), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n813), .A2(new_n816), .A3(new_n834), .A4(new_n831), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n790), .B1(new_n833), .B2(new_n835), .ZN(G311));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  XNOR2_X1  g412(.A(G311), .B(new_n837), .ZN(G150));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n555), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n543), .A2(G93), .B1(new_n841), .B2(new_n523), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT96), .B(G55), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n539), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n568), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n844), .A2(new_n566), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT38), .Z(new_n848));
  NOR2_X1   g423(.A1(new_n626), .A2(new_n634), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  AOI21_X1  g426(.A(G860), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n844), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(G145));
  NAND2_X1  g431(.A1(new_n470), .A2(G142), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n483), .A2(G130), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n464), .A2(G118), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT97), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n649), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n823), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT98), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n505), .B(new_n764), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n751), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n741), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n865), .A2(new_n868), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n865), .A2(KEYINPUT99), .A3(new_n868), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G160), .B(new_n487), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n646), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n868), .A2(KEYINPUT101), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n868), .A2(KEYINPUT101), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n864), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n871), .A3(new_n876), .ZN(new_n882));
  XNOR2_X1  g457(.A(KEYINPUT100), .B(G37), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT40), .B1(new_n877), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n874), .A2(new_n876), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n887), .A2(new_n888), .A3(new_n884), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n886), .A2(new_n889), .ZN(G395));
  XNOR2_X1  g465(.A(new_n626), .B(new_n631), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n847), .B(new_n636), .Z(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n891), .B2(new_n895), .ZN(new_n897));
  XNOR2_X1  g472(.A(G290), .B(new_n801), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n537), .B(G305), .Z(new_n899));
  OR2_X1    g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n904), .A2(new_n905), .B1(KEYINPUT42), .B2(new_n902), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n897), .B(new_n907), .ZN(new_n908));
  MUX2_X1   g483(.A(new_n844), .B(new_n908), .S(G868), .Z(G295));
  MUX2_X1   g484(.A(new_n844), .B(new_n908), .S(G868), .Z(G331));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  XNOR2_X1  g486(.A(G301), .B(G286), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n847), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n893), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n912), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n847), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n891), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n902), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n920), .A2(new_n883), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n914), .A2(new_n902), .A3(new_n917), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n911), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n911), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n920), .A2(KEYINPUT104), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n902), .B1(new_n914), .B2(new_n917), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(G37), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n924), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n923), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n920), .A2(new_n883), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n933), .A2(new_n924), .ZN(new_n934));
  INV_X1    g509(.A(new_n922), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n926), .B2(new_n929), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n932), .B(new_n934), .C1(new_n936), .C2(new_n911), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n931), .A2(new_n937), .ZN(G397));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n940), .A2(KEYINPUT4), .A3(new_n503), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n493), .A2(new_n497), .A3(new_n494), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n749), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n478), .B1(new_n946), .B2(new_n464), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n476), .A2(KEYINPUT66), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(new_n948), .A3(G40), .A4(new_n471), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n764), .B(G2067), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT106), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n945), .A2(new_n949), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT107), .ZN(new_n954));
  INV_X1    g529(.A(G1996), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT105), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n742), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n952), .A2(G1996), .A3(new_n741), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n823), .A2(new_n825), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT127), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G2067), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n764), .A2(new_n964), .ZN(new_n965));
  AOI211_X1 g540(.A(new_n945), .B(new_n949), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n952), .B1(new_n951), .B2(new_n741), .ZN(new_n967));
  INV_X1    g542(.A(new_n957), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n968), .A2(KEYINPUT46), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(KEYINPUT46), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT47), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n823), .B(new_n825), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n952), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n960), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(G290), .A2(G1986), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n952), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT48), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n966), .B(new_n972), .C1(new_n975), .C2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT126), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n827), .B1(new_n613), .B2(new_n614), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n952), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n975), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n596), .A2(G8), .A3(new_n597), .ZN(new_n985));
  NAND2_X1  g560(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n596), .A2(G8), .A3(new_n597), .A4(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n991));
  INV_X1    g566(.A(G40), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n477), .A2(new_n992), .A3(new_n479), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n945), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT108), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n945), .A2(new_n996), .A3(new_n991), .A4(new_n993), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n794), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n949), .B1(new_n943), .B2(KEYINPUT50), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n505), .A2(new_n1000), .A3(new_n939), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n730), .A3(new_n1001), .ZN(new_n1002));
  AOI221_X4 g577(.A(new_n984), .B1(new_n987), .B2(new_n990), .C1(new_n998), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n987), .A2(new_n990), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n998), .A2(new_n1002), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(G8), .B1(new_n943), .B2(new_n949), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT110), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1010), .B(G8), .C1(new_n943), .C2(new_n949), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G288), .A2(new_n807), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n807), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n606), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n520), .A2(G86), .A3(new_n534), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(new_n606), .A3(new_n607), .A4(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1021), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1024), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1012), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT112), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n494), .A2(new_n497), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n501), .B1(new_n749), .B2(new_n490), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n492), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n940), .A2(KEYINPUT4), .A3(new_n503), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1384), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n993), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1010), .B1(new_n1039), .B2(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1011), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1030), .B(new_n1033), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1032), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1020), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1042), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1033), .B1(new_n1012), .B2(new_n1030), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1017), .A2(new_n1015), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n994), .A2(new_n711), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n943), .A2(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g628(.A(G2084), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n993), .A4(new_n1001), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n984), .B(G286), .C1(new_n1052), .C2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1007), .A2(new_n1045), .A3(new_n1051), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1056), .A2(KEYINPUT63), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1048), .A2(new_n1050), .A3(KEYINPUT113), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n1020), .B2(new_n1043), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1007), .B(new_n1060), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n993), .B1(new_n1038), .B2(new_n1000), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1001), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1961), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n999), .A2(KEYINPUT116), .A3(new_n1001), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT45), .B1(new_n505), .B2(new_n939), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n949), .ZN(new_n1076));
  INV_X1    g651(.A(G2078), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1073), .A2(KEYINPUT120), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT120), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n995), .A2(new_n997), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT53), .B1(new_n1083), .B2(new_n1077), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1066), .B(G171), .C1(new_n1082), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1084), .B1(new_n1088), .B2(new_n1079), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT121), .B1(new_n1089), .B2(G301), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1007), .A2(new_n1045), .A3(new_n1051), .ZN(new_n1092));
  OAI211_X1 g667(.A(G168), .B(new_n1055), .C1(new_n1076), .C2(G1966), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G8), .ZN(new_n1094));
  AOI21_X1  g669(.A(G168), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1097), .A3(G8), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT62), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(KEYINPUT62), .A3(new_n1098), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1091), .A2(new_n1092), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1003), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1048), .A2(G1976), .A3(G288), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G305), .A2(G1981), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1012), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1065), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1007), .A2(new_n1045), .A3(new_n1051), .A4(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n946), .A2(KEYINPUT123), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n946), .A2(KEYINPUT123), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(G2105), .ZN(new_n1116));
  INV_X1    g691(.A(new_n471), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1117), .A2(KEYINPUT122), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1077), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1117), .B2(KEYINPUT122), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1113), .A2(new_n1116), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1073), .A2(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1084), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT125), .B1(new_n1123), .B2(G171), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT125), .B(G171), .C1(new_n1084), .C2(new_n1122), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1089), .B2(G301), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1112), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT124), .B1(new_n1123), .B2(G171), .ZN(new_n1131));
  OR4_X1    g706(.A1(KEYINPUT124), .A2(new_n1084), .A3(new_n1122), .A4(G171), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1128), .B1(new_n1091), .B2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1053), .A2(new_n993), .A3(new_n1001), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1076), .A2(new_n1135), .B1(new_n1136), .B2(new_n781), .ZN(new_n1137));
  OAI211_X1 g712(.A(KEYINPUT115), .B(new_n578), .C1(new_n588), .C2(new_n593), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n1139));
  NAND3_X1  g714(.A1(G299), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT76), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n591), .B1(new_n584), .B2(G65), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n511), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1143), .A2(new_n592), .B1(G91), .B2(new_n543), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1144), .B(new_n577), .C1(KEYINPUT115), .C2(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1137), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1070), .A2(new_n788), .A3(new_n1072), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1039), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n964), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n626), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1137), .A2(new_n1146), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1147), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT117), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n1150), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n627), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n626), .A4(new_n1150), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n1164));
  AND4_X1   g739(.A1(new_n945), .A2(new_n991), .A3(new_n993), .A4(new_n1135), .ZN(new_n1165));
  AOI21_X1  g740(.A(G1956), .B1(new_n999), .B2(new_n1001), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1145), .B(new_n1140), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1164), .B1(new_n1167), .B2(KEYINPUT119), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1147), .A2(new_n1167), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1147), .B(new_n1167), .C1(KEYINPUT119), .C2(new_n1164), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(KEYINPUT58), .B(G1341), .ZN(new_n1173));
  OAI22_X1  g748(.A1(new_n994), .A2(G1996), .B1(new_n1149), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n569), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1176), .A2(KEYINPUT118), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1175), .B(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1163), .A2(new_n1172), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1155), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1130), .A2(new_n1134), .A3(new_n1180), .ZN(new_n1181));
  AOI211_X1 g756(.A(new_n980), .B(new_n983), .C1(new_n1110), .C2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1096), .A2(KEYINPUT62), .A3(new_n1098), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1183), .A2(new_n1099), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1007), .A2(new_n1045), .A3(new_n1051), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1108), .B1(new_n1186), .B2(new_n1091), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1133), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT54), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1129), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1112), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1180), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1187), .B(new_n1065), .C1(new_n1190), .C2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n983), .ZN(new_n1195));
  AOI21_X1  g770(.A(KEYINPUT126), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n979), .B1(new_n1182), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g772(.A(new_n671), .ZN(new_n1199));
  NOR4_X1   g773(.A1(G229), .A2(new_n462), .A3(new_n1199), .A4(G227), .ZN(new_n1200));
  OAI21_X1  g774(.A(new_n1200), .B1(new_n887), .B2(new_n884), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n936), .A2(new_n911), .ZN(new_n1202));
  INV_X1    g776(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1201), .B1(new_n1203), .B2(new_n934), .ZN(G308));
  INV_X1    g778(.A(new_n934), .ZN(new_n1205));
  OAI221_X1 g779(.A(new_n1200), .B1(new_n887), .B2(new_n884), .C1(new_n1202), .C2(new_n1205), .ZN(G225));
endmodule


