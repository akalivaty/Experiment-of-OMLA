//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NOR2_X1   g0010(.A1(G58), .A2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT67), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n227), .B1(new_n223), .B2(new_n224), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n210), .B(new_n218), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT69), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT71), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(KEYINPUT70), .B(G50), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  NAND2_X1  g0051(.A1(new_n203), .A2(G20), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT76), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n247), .A2(KEYINPUT8), .ZN(new_n254));
  XOR2_X1   g0054(.A(KEYINPUT74), .B(G58), .Z(new_n255));
  AOI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(KEYINPUT8), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n216), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT75), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n262), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n253), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT73), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(new_n267), .A3(new_n215), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n266), .B2(new_n215), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G13), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n273), .A2(new_n216), .A3(G1), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n266), .A2(new_n215), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT73), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n268), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G1), .B2(new_n216), .ZN(new_n279));
  MUX2_X1   g0079(.A(new_n275), .B(new_n279), .S(G50), .Z(new_n280));
  NAND2_X1  g0080(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n286), .B1(new_n290), .B2(G226), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G222), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G77), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(G1698), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT72), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n296), .B1(new_n298), .B2(G223), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n291), .B1(new_n299), .B2(new_n288), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n300), .A2(G179), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n282), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(KEYINPUT78), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n272), .A2(new_n306), .A3(new_n280), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT78), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n300), .A2(new_n308), .B1(new_n309), .B2(KEYINPUT9), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  XOR2_X1   g0111(.A(KEYINPUT77), .B(G200), .Z(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n300), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n307), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n306), .B1(new_n272), .B2(new_n280), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT10), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n316), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n310), .B1(new_n300), .B2(new_n313), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .A4(new_n307), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n304), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G50), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n260), .A2(new_n323), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n257), .A2(new_n295), .B1(new_n216), .B2(G68), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n271), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G68), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n274), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT12), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n329), .B2(new_n279), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT80), .ZN(new_n334));
  INV_X1    g0134(.A(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G33), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n336), .A2(new_n338), .A3(G232), .A4(G1698), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n336), .A2(new_n338), .A3(G226), .A4(new_n293), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n288), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n286), .B1(new_n290), .B2(G238), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n345), .B1(new_n344), .B2(new_n346), .ZN(new_n348));
  OAI21_X1  g0148(.A(G169), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n349), .A2(KEYINPUT14), .B1(new_n350), .B2(G179), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT14), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(G169), .C1(new_n347), .C2(new_n348), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n334), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(KEYINPUT14), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n350), .A2(G179), .ZN(new_n356));
  AND4_X1   g0156(.A1(new_n334), .A2(new_n355), .A3(new_n353), .A4(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n333), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n333), .B1(G190), .B2(new_n350), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(new_n350), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n286), .B1(new_n290), .B2(G244), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n292), .A2(G232), .A3(new_n293), .ZN(new_n364));
  INV_X1    g0164(.A(G107), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n292), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n298), .B2(G238), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n363), .B1(new_n367), .B2(new_n288), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n308), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G20), .A2(G77), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT8), .B(G58), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n370), .B1(new_n371), .B2(new_n257), .C1(new_n260), .C2(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n271), .B1(new_n295), .B2(new_n274), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n295), .B2(new_n279), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n368), .A2(new_n313), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n368), .A2(new_n301), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n379), .A2(new_n375), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n368), .A2(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n322), .A2(new_n362), .A3(new_n378), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n336), .A2(new_n338), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n384), .A2(KEYINPUT81), .A3(KEYINPUT7), .A4(new_n216), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n292), .B2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(G20), .B1(new_n336), .B2(new_n338), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT81), .B1(new_n389), .B2(KEYINPUT7), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT74), .B(G58), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n211), .B1(new_n392), .B2(G68), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT82), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n260), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n259), .A2(KEYINPUT82), .A3(G159), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n394), .A2(G20), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n391), .A2(KEYINPUT16), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT83), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(new_n337), .A3(G33), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n386), .A2(G20), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n384), .C2(new_n402), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n329), .B1(new_n405), .B2(new_n387), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n397), .A2(new_n398), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n393), .B2(new_n216), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n401), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n400), .A2(new_n409), .A3(new_n271), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n256), .B1(new_n283), .B2(G20), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n274), .B1(new_n277), .B2(new_n268), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n411), .A2(new_n412), .B1(new_n274), .B2(new_n256), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT84), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT84), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n410), .A2(new_n416), .A3(new_n413), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G223), .A2(G1698), .ZN(new_n418));
  INV_X1    g0218(.A(G226), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n418), .B1(new_n419), .B2(G1698), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n292), .B1(G33), .B2(G87), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n288), .ZN(new_n422));
  INV_X1    g0222(.A(G179), .ZN(new_n423));
  INV_X1    g0223(.A(G232), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n289), .A2(new_n424), .B1(new_n285), .B2(new_n284), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n422), .A2(new_n425), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(G169), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n415), .A2(new_n417), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT18), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n360), .B1(new_n422), .B2(new_n425), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n427), .B2(G190), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n410), .A2(new_n433), .A3(new_n413), .A4(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n436), .A2(KEYINPUT86), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n410), .A2(new_n433), .A3(new_n413), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n436), .A2(KEYINPUT86), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n415), .A2(new_n443), .A3(new_n417), .A4(new_n429), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n431), .A2(new_n440), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n383), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n336), .A2(new_n338), .A3(G264), .A4(G1698), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n336), .A2(new_n338), .A3(G257), .A4(new_n293), .ZN(new_n448));
  INV_X1    g0248(.A(G303), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(new_n448), .C1(new_n449), .C2(new_n292), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n450), .A2(new_n343), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT90), .ZN(new_n452));
  INV_X1    g0252(.A(G41), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT5), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(KEYINPUT90), .B2(G41), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n454), .A2(new_n456), .A3(new_n283), .A4(G45), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(G270), .A3(new_n288), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n459), .A2(new_n285), .A3(G1), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n460), .A2(new_n288), .A3(new_n454), .A4(new_n456), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(G200), .B1(new_n451), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT95), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n283), .A2(G33), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n275), .B(new_n465), .C1(new_n269), .C2(new_n270), .ZN(new_n466));
  INV_X1    g0266(.A(G116), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n412), .A2(KEYINPUT95), .A3(G116), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n458), .A2(new_n461), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n450), .A2(new_n343), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(G190), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT20), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n216), .A2(G116), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n215), .B2(new_n266), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n216), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT88), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(KEYINPUT88), .A2(G97), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n479), .B1(new_n484), .B2(new_n335), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n474), .B1(new_n477), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT88), .A2(G97), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT88), .A2(G97), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G33), .ZN(new_n490));
  OAI211_X1 g0290(.A(KEYINPUT20), .B(new_n476), .C1(new_n490), .C2(new_n479), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n273), .A2(G1), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n486), .A2(new_n491), .B1(new_n492), .B2(new_n475), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n463), .A2(new_n470), .A3(new_n473), .A4(new_n493), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n494), .B(KEYINPUT96), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n470), .A2(new_n493), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n301), .B1(new_n471), .B2(new_n472), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT21), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n496), .A2(KEYINPUT21), .A3(new_n497), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n451), .A2(new_n423), .A3(new_n462), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  AND2_X1   g0306(.A1(G97), .A2(G107), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n365), .A2(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n489), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G20), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n259), .A2(G77), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT87), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT87), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n259), .A2(new_n515), .A3(G77), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n365), .B1(new_n405), .B2(new_n387), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n271), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n466), .A2(new_n481), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n274), .A2(new_n481), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT89), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n521), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n336), .A2(new_n338), .A3(G244), .A4(new_n293), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n478), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n343), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n457), .A2(G257), .A3(new_n288), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n461), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n301), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n533), .B2(new_n343), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n423), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n527), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n534), .A2(new_n537), .A3(new_n308), .ZN(new_n544));
  AOI21_X1  g0344(.A(G200), .B1(new_n534), .B2(new_n537), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT91), .B1(new_n546), .B2(new_n527), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n534), .A2(new_n537), .A3(new_n308), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G200), .B2(new_n540), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT83), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n403), .A2(new_n404), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n550), .A2(new_n551), .B1(new_n389), .B2(KEYINPUT7), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n517), .B1(new_n511), .B2(G20), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n278), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n555), .A2(new_n522), .A3(new_n525), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT91), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n549), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n543), .B1(new_n547), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n336), .A2(new_n338), .A3(new_n216), .A4(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT22), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT22), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n292), .A2(new_n562), .A3(new_n216), .A4(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT24), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G116), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(G20), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n216), .B2(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n365), .A2(KEYINPUT23), .A3(G20), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n565), .B1(new_n564), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n271), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n274), .A2(new_n365), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT25), .ZN(new_n576));
  INV_X1    g0376(.A(new_n466), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(G107), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n336), .A2(new_n338), .A3(G250), .A4(new_n293), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n336), .A2(new_n338), .A3(G257), .A4(G1698), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G294), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT97), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n288), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT97), .A4(new_n582), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n457), .A2(G264), .A3(new_n288), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n461), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n301), .ZN(new_n590));
  INV_X1    g0390(.A(new_n588), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n585), .B2(new_n586), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n423), .A3(new_n461), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n579), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n589), .A2(G200), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(G190), .A3(new_n461), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n574), .A3(new_n578), .A4(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n336), .A2(new_n338), .A3(G238), .A4(new_n293), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n336), .A2(new_n338), .A3(G244), .A4(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n566), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n343), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT92), .B1(new_n459), .B2(G1), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT92), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n283), .A3(G45), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n288), .A2(new_n602), .A3(new_n604), .A4(G250), .ZN(new_n605));
  INV_X1    g0405(.A(new_n460), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n312), .B1(new_n601), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n371), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(new_n275), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n335), .A2(G20), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n487), .B2(new_n488), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G87), .A2(G107), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n482), .A2(new_n483), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n216), .B1(new_n341), .B2(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n336), .A2(new_n338), .A3(new_n216), .A4(G68), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n615), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n611), .B1(new_n621), .B2(new_n271), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n412), .A2(G87), .A3(new_n465), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n609), .A2(KEYINPUT94), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT94), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n257), .B1(new_n482), .B2(new_n483), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n620), .B1(new_n626), .B2(KEYINPUT19), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n617), .A2(new_n618), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n271), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n611), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n623), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n625), .B1(new_n631), .B2(new_n608), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n601), .A2(G190), .A3(new_n607), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n624), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n601), .A2(new_n423), .A3(new_n607), .ZN(new_n635));
  AOI21_X1  g0435(.A(G169), .B1(new_n601), .B2(new_n607), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n412), .A2(new_n610), .A3(new_n465), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n622), .A2(KEYINPUT93), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT93), .B1(new_n622), .B2(new_n638), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n594), .A2(new_n597), .A3(new_n634), .A4(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n446), .A2(new_n505), .A3(new_n559), .A4(new_n642), .ZN(G372));
  AOI21_X1  g0443(.A(new_n428), .B1(new_n410), .B2(new_n413), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT18), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n351), .A2(new_n353), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT80), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n351), .A2(new_n334), .A3(new_n353), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n380), .A2(new_n381), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n649), .A2(new_n333), .B1(new_n650), .B2(new_n361), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n441), .B1(new_n437), .B2(new_n439), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n645), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(KEYINPUT102), .B1(new_n317), .B2(new_n321), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT102), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n656), .B(new_n645), .C1(new_n651), .C2(new_n653), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n304), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n601), .A2(G190), .A3(new_n607), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n608), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT98), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n661), .A2(new_n629), .A3(new_n630), .A4(new_n623), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(new_n622), .B2(new_n623), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n641), .A2(new_n664), .A3(KEYINPUT99), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT99), .B1(new_n641), .B2(new_n664), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n543), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(KEYINPUT101), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT101), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT99), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n601), .A2(new_n423), .A3(new_n607), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n605), .A2(new_n606), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n343), .B2(new_n600), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(G169), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n629), .A2(new_n630), .A3(new_n638), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT93), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n622), .A2(KEYINPUT93), .A3(new_n638), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n633), .B1(new_n312), .B2(new_n674), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n631), .A2(KEYINPUT98), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n622), .A2(new_n661), .A3(new_n623), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n671), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n641), .A2(new_n664), .A3(KEYINPUT99), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n542), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n670), .B1(new_n687), .B2(KEYINPUT26), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n543), .A2(KEYINPUT26), .A3(new_n641), .A4(new_n634), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n669), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n665), .A2(new_n666), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n549), .A2(new_n556), .A3(new_n557), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n557), .B1(new_n549), .B2(new_n556), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n542), .B(new_n597), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n504), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT100), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n594), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n594), .A2(new_n697), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n680), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n690), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n446), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n658), .A2(new_n703), .ZN(G369));
  NAND2_X1  g0504(.A1(new_n492), .A2(new_n216), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n496), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n505), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n696), .B2(new_n711), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n597), .A2(new_n594), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n579), .A2(new_n710), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n710), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n594), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n696), .A2(new_n710), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n715), .ZN(new_n722));
  OR3_X1    g0522(.A1(new_n698), .A2(new_n699), .A3(new_n710), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n720), .A2(new_n725), .ZN(G399));
  INV_X1    g0526(.A(new_n207), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G1), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n489), .A2(new_n467), .A3(new_n616), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(new_n213), .B2(new_n729), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  AOI211_X1 g0533(.A(KEYINPUT29), .B(new_n710), .C1(new_n690), .C2(new_n701), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT29), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n685), .A2(new_n686), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n594), .A2(new_n501), .A3(new_n500), .A4(new_n503), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n559), .A2(new_n736), .A3(new_n597), .A4(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT104), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n543), .A2(new_n634), .A3(new_n668), .A4(new_n641), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT103), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n641), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n747));
  INV_X1    g0547(.A(new_n694), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(KEYINPUT104), .A3(new_n736), .A4(new_n737), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n740), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n735), .B1(new_n750), .B2(new_n718), .ZN(new_n751));
  INV_X1    g0551(.A(G330), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n502), .A2(new_n592), .A3(new_n540), .A4(new_n674), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AND4_X1   g0555(.A1(G179), .A2(new_n674), .A3(new_n472), .A4(new_n471), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n756), .A2(KEYINPUT30), .A3(new_n540), .A4(new_n592), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n601), .A2(new_n607), .ZN(new_n758));
  AOI21_X1  g0558(.A(G179), .B1(new_n471), .B2(new_n472), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n589), .A2(new_n538), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n755), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n710), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT31), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT31), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n761), .A2(new_n764), .A3(new_n710), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n505), .A2(new_n642), .A3(new_n559), .A4(new_n718), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n752), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n734), .A2(new_n751), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n733), .B1(new_n769), .B2(G1), .ZN(G364));
  NOR2_X1   g0570(.A1(new_n713), .A2(G330), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n273), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n283), .B1(new_n772), .B2(G45), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n771), .B(new_n714), .C1(new_n729), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n773), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n728), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n292), .A2(G355), .A3(new_n207), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G116), .B2(new_n207), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n250), .A2(new_n459), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n727), .A2(new_n292), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n459), .B2(new_n214), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n778), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n215), .B1(G20), .B2(new_n301), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n776), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n216), .A2(G190), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G179), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n292), .B1(new_n794), .B2(G329), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n216), .B1(new_n792), .B2(G190), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n216), .A2(new_n308), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n423), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n791), .A2(new_n800), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n801), .A2(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n423), .A2(new_n360), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n808), .A2(G326), .ZN(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT33), .B(G317), .Z(new_n810));
  NAND2_X1  g0610(.A1(new_n806), .A2(new_n791), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR4_X1   g0612(.A1(new_n798), .A2(new_n805), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G283), .ZN(new_n814));
  INV_X1    g0614(.A(new_n791), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n312), .A2(G179), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n313), .A2(new_n423), .A3(new_n799), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT105), .Z(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n813), .B1(new_n814), .B2(new_n817), .C1(new_n820), .C2(new_n449), .ZN(new_n821));
  INV_X1    g0621(.A(new_n803), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G77), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n823), .B1(new_n329), .B2(new_n811), .C1(new_n255), .C2(new_n801), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G107), .B2(new_n816), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n794), .A2(G159), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT32), .ZN(new_n827));
  INV_X1    g0627(.A(new_n797), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G97), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(new_n292), .C1(new_n323), .C2(new_n807), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G87), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n825), .B(new_n831), .C1(new_n832), .C2(new_n818), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n821), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n790), .B1(new_n787), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n786), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n713), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT106), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n774), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  AOI21_X1  g0640(.A(new_n710), .B1(new_n690), .B2(new_n701), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n382), .A2(new_n710), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n375), .A2(new_n710), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n378), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n842), .B1(new_n844), .B2(new_n382), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n841), .B(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n768), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n776), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n292), .B1(new_n819), .B2(G107), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT108), .Z(new_n851));
  NOR2_X1   g0651(.A1(new_n817), .A2(new_n832), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n794), .A2(G311), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n853), .B1(new_n796), .B2(new_n801), .C1(new_n449), .C2(new_n807), .ZN(new_n854));
  XOR2_X1   g0654(.A(KEYINPUT107), .B(G283), .Z(new_n855));
  OAI221_X1 g0655(.A(new_n829), .B1(new_n467), .B2(new_n803), .C1(new_n811), .C2(new_n855), .ZN(new_n856));
  NOR4_X1   g0656(.A1(new_n851), .A2(new_n852), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n816), .A2(G68), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n292), .B1(new_n793), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n392), .B2(new_n828), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n858), .B(new_n861), .C1(new_n820), .C2(new_n323), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT110), .ZN(new_n863));
  INV_X1    g0663(.A(new_n811), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G137), .A2(new_n808), .B1(new_n864), .B2(G150), .ZN(new_n865));
  XNOR2_X1  g0665(.A(KEYINPUT109), .B(G143), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n865), .B1(new_n396), .B2(new_n803), .C1(new_n801), .C2(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT34), .Z(new_n868));
  NOR2_X1   g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n787), .B1(new_n857), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n787), .A2(new_n784), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n775), .B(new_n728), .C1(new_n295), .C2(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n870), .B(new_n872), .C1(new_n845), .C2(new_n785), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n849), .A2(new_n873), .ZN(G384));
  OR2_X1    g0674(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(G116), .A3(new_n217), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT36), .Z(new_n878));
  OAI211_X1 g0678(.A(new_n214), .B(G77), .C1(new_n255), .C2(new_n329), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n323), .A2(G68), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT111), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n283), .B(G13), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n333), .A2(new_n710), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n358), .A2(new_n361), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n649), .A2(new_n333), .A3(new_n710), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n766), .A2(new_n767), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n845), .ZN(new_n889));
  INV_X1    g0689(.A(new_n413), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n400), .A2(new_n271), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n391), .A2(new_n399), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n401), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(new_n708), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n445), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n438), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n410), .A2(new_n416), .A3(new_n413), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n416), .B1(new_n410), .B2(new_n413), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n901), .B2(new_n429), .ZN(new_n902));
  INV_X1    g0702(.A(new_n708), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n415), .A2(new_n417), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n438), .B1(new_n894), .B2(new_n708), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n894), .A2(new_n428), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT37), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n410), .A2(new_n433), .A3(new_n413), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n644), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n904), .A2(new_n902), .B1(new_n914), .B2(KEYINPUT37), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n904), .B1(new_n652), .B2(new_n645), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n889), .B1(new_n910), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n909), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n896), .B2(new_n909), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n887), .A2(new_n888), .A3(new_n919), .A4(new_n845), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n918), .A2(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n924), .A2(new_n446), .A3(new_n888), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n446), .B2(new_n888), .ZN(new_n926));
  OR3_X1    g0726(.A1(new_n925), .A2(new_n926), .A3(new_n752), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n844), .A2(new_n382), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n650), .A2(new_n718), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n710), .B(new_n930), .C1(new_n690), .C2(new_n701), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n887), .B1(new_n920), .B2(new_n921), .C1(new_n931), .C2(new_n842), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n645), .A2(new_n903), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT39), .B1(new_n910), .B2(new_n917), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n896), .A2(new_n909), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n911), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n358), .A2(new_n710), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n932), .B(new_n934), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n446), .B1(new_n734), .B2(new_n751), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n658), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n943), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n927), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n283), .B2(new_n772), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n927), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n883), .B1(new_n948), .B2(new_n949), .ZN(G367));
  NAND3_X1  g0750(.A1(new_n682), .A2(new_n683), .A3(new_n710), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n736), .A2(KEYINPUT112), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n641), .B2(new_n951), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT112), .B1(new_n736), .B2(new_n951), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n836), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n292), .B1(new_n797), .B2(new_n329), .C1(new_n396), .C2(new_n811), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n807), .A2(new_n866), .B1(new_n801), .B2(new_n258), .ZN(new_n959));
  INV_X1    g0759(.A(G137), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n803), .A2(new_n323), .B1(new_n793), .B2(new_n960), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n816), .A2(G77), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(new_n255), .C2(new_n818), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G311), .A2(new_n808), .B1(new_n864), .B2(G294), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n449), .B2(new_n801), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n292), .B(new_n966), .C1(G317), .C2(new_n794), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n855), .A2(new_n803), .B1(new_n797), .B2(new_n365), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT114), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n967), .B(new_n969), .C1(new_n489), .C2(new_n817), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n818), .A2(KEYINPUT46), .A3(new_n467), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n819), .A2(G116), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n971), .B1(new_n972), .B2(KEYINPUT46), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n964), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT47), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n787), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n240), .A2(new_n780), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n977), .B(new_n788), .C1(new_n207), .C2(new_n371), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n776), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n957), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n527), .A2(new_n710), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n559), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT113), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n543), .A2(new_n710), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT113), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n559), .A2(new_n987), .A3(new_n983), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n982), .B1(new_n990), .B2(new_n724), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n725), .A2(new_n989), .A3(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n725), .B2(new_n989), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n990), .A2(KEYINPUT44), .A3(new_n724), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(new_n714), .A3(new_n719), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n993), .A2(new_n997), .A3(new_n720), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n722), .B1(new_n719), .B2(new_n721), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n714), .B(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n999), .A2(new_n769), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n769), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n728), .B(KEYINPUT41), .Z(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n775), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n989), .A2(new_n715), .A3(new_n721), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT42), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n594), .B1(new_n985), .B2(new_n988), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n718), .B1(new_n1010), .B2(new_n543), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(KEYINPUT42), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1015), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1017), .A2(new_n1018), .B1(new_n720), .B2(new_n990), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1018), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n720), .A2(new_n990), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n1021), .A3(new_n1016), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n981), .B1(new_n1007), .B2(new_n1023), .ZN(G387));
  NAND2_X1  g0824(.A1(new_n1002), .A2(new_n775), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n719), .A2(new_n836), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n807), .A2(new_n396), .B1(new_n801), .B2(new_n323), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n292), .B1(new_n793), .B2(new_n258), .C1(new_n371), .C2(new_n797), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G68), .C2(new_n822), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n818), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n256), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1030), .A2(G77), .B1(new_n1031), .B2(new_n864), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1029), .B(new_n1032), .C1(new_n481), .C2(new_n817), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n292), .B1(new_n794), .B2(G326), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n818), .A2(new_n796), .B1(new_n797), .B2(new_n855), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n807), .A2(new_n802), .B1(new_n811), .B2(new_n804), .ZN(new_n1036));
  INV_X1    g0836(.A(G317), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n801), .A2(new_n1037), .B1(new_n803), .B2(new_n449), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1035), .B1(new_n1039), .B2(KEYINPUT48), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(KEYINPUT48), .B2(new_n1039), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT49), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1034), .B1(new_n467), .B2(new_n817), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n787), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n236), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n780), .B1(new_n1047), .B2(new_n459), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n731), .A2(new_n207), .A3(new_n292), .ZN(new_n1049));
  AOI211_X1 g0849(.A(G45), .B(new_n731), .C1(G68), .C2(G77), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n372), .A2(G50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1048), .A2(new_n1049), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n207), .A2(G107), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n788), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1046), .A2(new_n776), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n769), .A2(new_n1002), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n728), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n769), .A2(new_n1002), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1025), .B1(new_n1026), .B2(new_n1056), .C1(new_n1058), .C2(new_n1059), .ZN(G393));
  NAND2_X1  g0860(.A1(new_n999), .A2(new_n1000), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n1057), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(new_n728), .A3(new_n1003), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(KEYINPUT115), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT115), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n999), .A2(new_n1065), .A3(new_n1000), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n775), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n245), .A2(new_n781), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n788), .B1(new_n207), .B2(new_n489), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n776), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n797), .A2(new_n295), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n292), .B1(new_n811), .B2(new_n323), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n803), .A2(new_n372), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n793), .A2(new_n866), .ZN(new_n1074));
  OR4_X1    g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT51), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n807), .A2(new_n258), .B1(new_n801), .B2(new_n396), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1030), .A2(G68), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n1076), .B2(new_n1077), .C1(new_n832), .C2(new_n817), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n807), .A2(new_n1037), .B1(new_n801), .B2(new_n804), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n365), .B2(new_n817), .C1(new_n818), .C2(new_n855), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G303), .A2(new_n864), .B1(new_n822), .B2(G294), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n292), .B1(new_n794), .B2(G322), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n467), .C2(new_n797), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1075), .A2(new_n1079), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1070), .B1(new_n1087), .B2(new_n787), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n989), .B2(new_n836), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1063), .A2(new_n1067), .A3(new_n1089), .ZN(G390));
  NAND3_X1  g0890(.A1(new_n888), .A2(new_n845), .A3(G330), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n887), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n750), .A2(new_n718), .A3(new_n928), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n768), .A2(new_n845), .A3(new_n887), .ZN(new_n1095));
  AND4_X1   g0895(.A1(new_n929), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n702), .A2(new_n718), .A3(new_n845), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1097), .A2(new_n929), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n446), .A2(new_n768), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n658), .A2(new_n944), .A3(new_n1100), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n887), .B1(new_n931), .B2(new_n842), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1103), .A2(new_n942), .B1(new_n936), .B2(new_n939), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n910), .A2(new_n917), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n942), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1094), .A2(new_n929), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n887), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1095), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1104), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n842), .B1(new_n841), .B2(new_n845), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n942), .B1(new_n1111), .B2(new_n1092), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n940), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1107), .A2(new_n887), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n942), .A3(new_n1105), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1095), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1102), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1109), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1113), .A2(new_n1115), .A3(new_n1095), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n728), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1118), .A2(new_n775), .A3(new_n1119), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n871), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n776), .B1(new_n1031), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n818), .A2(new_n258), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n807), .A2(new_n1129), .B1(new_n801), .B2(new_n859), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT117), .Z(new_n1131));
  NAND2_X1  g0931(.A1(new_n816), .A2(G50), .ZN(new_n1132));
  INV_X1    g0932(.A(G125), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n292), .B1(new_n793), .B2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n811), .A2(new_n960), .B1(new_n803), .B2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(G159), .C2(new_n828), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n820), .A2(new_n832), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n292), .B(new_n1071), .C1(G283), .C2(new_n808), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n811), .A2(new_n365), .B1(new_n803), .B2(new_n489), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n801), .A2(new_n467), .B1(new_n793), .B2(new_n796), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n858), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1138), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1125), .B1(new_n1145), .B2(new_n787), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n935), .B1(new_n922), .B2(KEYINPUT39), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n785), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1123), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1122), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT119), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1122), .A2(new_n1149), .A3(KEYINPUT119), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(G378));
  OAI21_X1  g0955(.A(new_n776), .B1(new_n1124), .B2(G50), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1030), .A2(G77), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n453), .B(new_n384), .C1(new_n807), .C2(new_n467), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G68), .B2(new_n828), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n801), .A2(new_n365), .B1(new_n803), .B2(new_n371), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n811), .A2(new_n481), .B1(new_n793), .B2(new_n814), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n816), .A2(new_n392), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1157), .A2(new_n1159), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT58), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n453), .B1(new_n337), .B2(new_n335), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1164), .A2(new_n1165), .B1(new_n323), .B2(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n811), .A2(new_n859), .B1(new_n803), .B2(new_n960), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n807), .A2(new_n1133), .B1(new_n801), .B2(new_n1129), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(G150), .C2(new_n828), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n818), .B2(new_n1135), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n816), .A2(G159), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G33), .B(G41), .C1(new_n794), .C2(G124), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1167), .B1(new_n1165), .B2(new_n1164), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1156), .B1(new_n1177), .B2(new_n787), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n317), .A2(new_n321), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n304), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n281), .A2(new_n903), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT120), .Z(new_n1185));
  INV_X1    g0985(.A(new_n1182), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n322), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1183), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1185), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n322), .A2(new_n1186), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1182), .B(new_n304), .C1(new_n317), .C2(new_n321), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1178), .B1(new_n1193), .B2(new_n785), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1193), .B1(new_n924), .B2(G330), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n887), .A2(new_n888), .A3(new_n845), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n919), .B1(new_n1105), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n923), .B1(new_n938), .B2(new_n910), .ZN(new_n1199));
  OAI211_X1 g0999(.A(G330), .B(new_n1193), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n943), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(G330), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1193), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n933), .B1(new_n1147), .B2(new_n941), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n932), .A4(new_n1200), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1195), .B1(new_n1208), .B2(new_n775), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1101), .B(KEYINPUT121), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1121), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT122), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1202), .A2(new_n1212), .A3(new_n1207), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n943), .B(KEYINPUT122), .C1(new_n1196), .C2(new_n1201), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1213), .A3(KEYINPUT57), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n728), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT57), .B1(new_n1211), .B2(new_n1208), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1209), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT123), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1102), .A2(new_n1006), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1099), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1092), .A2(new_n784), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n776), .B1(new_n1124), .B2(G68), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n819), .A2(G97), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n467), .A2(new_n811), .B1(new_n801), .B2(new_n814), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n807), .A2(new_n796), .B1(new_n803), .B2(new_n365), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n384), .B1(new_n793), .B2(new_n449), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n610), .B2(new_n828), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1226), .A2(new_n963), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n807), .A2(new_n859), .B1(new_n801), .B2(new_n960), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1135), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n864), .B2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT124), .Z(new_n1236));
  OAI221_X1 g1036(.A(new_n292), .B1(new_n793), .B2(new_n1129), .C1(new_n258), .C2(new_n803), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G50), .B2(new_n828), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1163), .A3(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n820), .A2(new_n396), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1232), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1225), .B1(new_n1241), .B2(new_n787), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1223), .A2(new_n775), .B1(new_n1224), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1222), .A2(new_n1243), .ZN(G381));
  INV_X1    g1044(.A(new_n1150), .ZN(new_n1245));
  OR4_X1    g1045(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1246), .A2(G387), .A3(G381), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1219), .A2(new_n1245), .A3(new_n1247), .ZN(G407));
  NAND2_X1  g1048(.A1(new_n1219), .A2(new_n1245), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(new_n1249), .C2(G343), .ZN(G409));
  INV_X1    g1050(.A(G390), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G387), .A2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G390), .B(new_n981), .C1(new_n1007), .C2(new_n1023), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT126), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n773), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1023), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n980), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1255), .B1(new_n1259), .B2(G390), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(G393), .B(new_n839), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1254), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1261), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1252), .A2(new_n1253), .A3(new_n1263), .A4(new_n1255), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1211), .A2(new_n1006), .A3(new_n1208), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1213), .A2(new_n775), .A3(new_n1214), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1194), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1245), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1218), .B2(new_n1154), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n709), .A2(G213), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1102), .A2(KEYINPUT60), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1273), .A2(new_n1221), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n728), .B1(new_n1273), .B2(new_n1221), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1243), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G384), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G384), .B(new_n1243), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1271), .A2(new_n1272), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT125), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT125), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1271), .A2(new_n1283), .A3(new_n1272), .A4(new_n1280), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT62), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n709), .A2(G213), .A3(G2897), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1278), .A2(new_n1279), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT61), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1281), .A2(KEYINPUT62), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1266), .B1(new_n1285), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1282), .A2(new_n1295), .A3(new_n1284), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1265), .B2(new_n1298), .ZN(new_n1299));
  AOI211_X1 g1099(.A(KEYINPUT127), .B(KEYINPUT61), .C1(new_n1262), .C2(new_n1264), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1281), .A2(new_n1295), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1296), .A2(new_n1301), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1294), .A2(new_n1304), .ZN(G405));
  NOR2_X1   g1105(.A1(new_n1218), .A2(KEYINPUT123), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT123), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1217), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n728), .A3(new_n1215), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1307), .B1(new_n1309), .B2(new_n1209), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1306), .A2(new_n1310), .A3(new_n1150), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1218), .A2(new_n1154), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1266), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1312), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1265), .B(new_n1314), .C1(new_n1219), .C2(new_n1150), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1313), .A2(new_n1315), .A3(new_n1280), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1280), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(G402));
endmodule


