//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT64), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G137), .A4(new_n461), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n462), .A2(new_n461), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT65), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n462), .A2(new_n476), .A3(new_n461), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n462), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n467), .A2(new_n469), .A3(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(KEYINPUT66), .ZN(new_n484));
  OAI21_X1  g059(.A(G124), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n479), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n479), .A2(new_n485), .A3(KEYINPUT67), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n461), .B2(G114), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G102), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n461), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n494), .A2(new_n496), .A3(G2104), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n503), .A2(new_n494), .A3(KEYINPUT69), .A4(new_n496), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n483), .A2(G126), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n461), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n505), .A2(new_n506), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n501), .A2(new_n504), .B1(G126), .B2(new_n483), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n507), .B(KEYINPUT4), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(KEYINPUT70), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(G164));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G62), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G651), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n527), .A2(new_n529), .A3(G50), .A4(G543), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n520), .A2(new_n522), .A3(new_n527), .A4(new_n529), .ZN(new_n531));
  INV_X1    g106(.A(G88), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n535), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n526), .B1(new_n534), .B2(new_n536), .ZN(G166));
  AND2_X1   g112(.A1(new_n527), .A2(new_n529), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  INV_X1    g116(.A(new_n531), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G89), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n541), .A2(new_n543), .A3(new_n544), .A4(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  AOI22_X1  g123(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n518), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n539), .A2(new_n551), .B1(new_n552), .B2(new_n531), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n550), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n518), .ZN(new_n557));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n539), .A2(new_n558), .B1(new_n559), .B2(new_n531), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  XOR2_X1   g139(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n565));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n520), .A2(new_n522), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  INV_X1    g145(.A(G78), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n569), .A2(new_n570), .B1(new_n571), .B2(new_n519), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI221_X1 g149(.A(KEYINPUT73), .B1(new_n571), .B2(new_n519), .C1(new_n569), .C2(new_n570), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(G651), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n538), .A2(G53), .A3(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n538), .A2(new_n579), .A3(G53), .A4(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n542), .A2(G91), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n576), .A2(new_n581), .A3(new_n582), .ZN(G299));
  XNOR2_X1  g158(.A(G166), .B(KEYINPUT74), .ZN(G303));
  OAI21_X1  g159(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI221_X1 g162(.A(new_n585), .B1(new_n586), .B2(new_n531), .C1(new_n587), .C2(new_n539), .ZN(G288));
  INV_X1    g163(.A(G73), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT75), .B1(new_n589), .B2(new_n519), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(G73), .A3(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n590), .B(new_n592), .C1(new_n569), .C2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n540), .A2(G48), .B1(new_n594), .B2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n542), .A2(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n518), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n539), .A2(new_n600), .B1(new_n601), .B2(new_n531), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n531), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT10), .B1(new_n531), .B2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n610), .A2(new_n518), .B1(new_n611), .B2(new_n539), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n605), .B1(G868), .B2(new_n613), .ZN(G284));
  OAI21_X1  g189(.A(new_n605), .B1(G868), .B2(new_n613), .ZN(G321));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(G168), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(G168), .A2(new_n617), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G299), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n620), .B2(new_n616), .ZN(G297));
  OAI21_X1  g196(.A(new_n618), .B1(new_n620), .B2(new_n616), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n613), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n613), .A2(new_n623), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT77), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n478), .A2(G135), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT78), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n483), .B(KEYINPUT66), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G123), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n478), .A2(KEYINPUT78), .A3(G135), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n632), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT15), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n652), .A2(G2435), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(G2435), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT81), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n649), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n648), .A3(new_n662), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n667), .A3(G14), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  XOR2_X1   g246(.A(G2067), .B(G2678), .Z(new_n672));
  AOI21_X1  g247(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n671), .B(KEYINPUT17), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n673), .B1(new_n675), .B2(new_n672), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT82), .ZN(new_n677));
  INV_X1    g252(.A(new_n671), .ZN(new_n678));
  INV_X1    g253(.A(new_n672), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n679), .A3(new_n670), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n675), .A2(new_n670), .A3(new_n672), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  OR3_X1    g272(.A1(new_n690), .A2(new_n693), .A3(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  INV_X1    g277(.A(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1986), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n701), .B(new_n705), .Z(G229));
  NAND2_X1  g281(.A1(G288), .A2(G16), .ZN(new_n707));
  INV_X1    g282(.A(G23), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G16), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT33), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n707), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n712), .A2(G1976), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G1976), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n713), .B1(new_n707), .B2(new_n710), .ZN(new_n717));
  AOI211_X1 g292(.A(KEYINPUT33), .B(new_n709), .C1(G288), .C2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(KEYINPUT85), .A2(G16), .ZN(new_n720));
  NOR2_X1   g295(.A1(KEYINPUT85), .A2(G16), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G22), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G166), .B2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G1971), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n715), .A2(new_n719), .A3(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n725), .A2(G1971), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n729), .A2(G6), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G305), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT32), .B(G1981), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT86), .B(KEYINPUT34), .Z(new_n735));
  NAND4_X1  g310(.A1(new_n727), .A2(new_n728), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n735), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n715), .A2(new_n719), .A3(new_n728), .A4(new_n726), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n733), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n636), .A2(G119), .B1(new_n478), .B2(G131), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n461), .A2(G107), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT84), .B(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT35), .B(G1991), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n744), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G25), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n745), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n747), .B1(new_n745), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n723), .A2(G24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n603), .B2(new_n723), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1986), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n750), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n736), .A2(new_n739), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT87), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n757), .A2(new_n758), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(G162), .A2(new_n744), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n744), .A2(G35), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n748), .B1(new_n490), .B2(new_n491), .ZN(new_n770));
  OAI21_X1  g345(.A(KEYINPUT29), .B1(new_n770), .B2(new_n767), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n769), .A2(new_n771), .A3(G2090), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(KEYINPUT91), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n769), .A2(new_n771), .A3(new_n774), .A4(G2090), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n639), .ZN(new_n777));
  INV_X1    g352(.A(G29), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT90), .B(KEYINPUT30), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G28), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n777), .A2(new_n744), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(G29), .A2(G32), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n636), .A2(G129), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n478), .A2(G141), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n783), .A2(new_n784), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n782), .B1(new_n788), .B2(new_n778), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT27), .B(G1996), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(G2090), .B1(new_n769), .B2(new_n771), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n723), .A2(G19), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n561), .B2(new_n723), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT88), .B(G1341), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(G164), .A2(new_n744), .ZN(new_n797));
  INV_X1    g372(.A(G2078), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n744), .A2(G27), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n798), .B1(new_n797), .B2(new_n799), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n792), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n776), .A2(new_n781), .A3(new_n791), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G171), .A2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G5), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n729), .A2(G4), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n613), .B2(new_n729), .ZN(new_n810));
  INV_X1    g385(.A(G1348), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT31), .B(G11), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n636), .A2(G128), .B1(new_n478), .B2(G140), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n461), .A2(G116), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n748), .A2(G26), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n818), .A2(G29), .B1(KEYINPUT28), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(KEYINPUT28), .B2(new_n819), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G2067), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n804), .A2(new_n808), .A3(new_n814), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n789), .A2(new_n790), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT24), .B(G34), .ZN(new_n825));
  AOI22_X1  g400(.A1(G160), .A2(G29), .B1(new_n748), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G2084), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n806), .B2(new_n807), .ZN(new_n828));
  AND4_X1   g403(.A1(new_n764), .A2(new_n823), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(G299), .A2(G16), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n723), .A2(KEYINPUT23), .A3(G20), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT23), .ZN(new_n832));
  INV_X1    g407(.A(G20), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n722), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT92), .B(G1956), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n478), .A2(G139), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT25), .Z(new_n840));
  AOI22_X1  g415(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(new_n840), .C1(new_n461), .C2(new_n841), .ZN(new_n842));
  MUX2_X1   g417(.A(G33), .B(new_n842), .S(G29), .Z(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(G2072), .Z(new_n844));
  NAND2_X1  g419(.A1(G168), .A2(G16), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G16), .B2(G21), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT89), .B(G1966), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n829), .A2(new_n837), .A3(new_n844), .A4(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(G311));
  INV_X1    g426(.A(KEYINPUT93), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n823), .A2(new_n824), .A3(new_n828), .ZN(new_n854));
  INV_X1    g429(.A(new_n764), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n854), .A2(new_n855), .A3(new_n848), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n856), .A2(KEYINPUT93), .A3(new_n837), .A4(new_n844), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n857), .ZN(G150));
  XNOR2_X1  g433(.A(KEYINPUT94), .B(G55), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n540), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT95), .B(G93), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n542), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(new_n518), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G860), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT37), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n863), .B2(new_n865), .ZN(new_n871));
  INV_X1    g446(.A(new_n865), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n872), .A2(KEYINPUT96), .A3(new_n862), .A4(new_n860), .ZN(new_n873));
  INV_X1    g448(.A(new_n561), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n866), .A2(KEYINPUT96), .A3(new_n561), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n613), .A2(G559), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT97), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n867), .B1(new_n880), .B2(new_n881), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n869), .B1(new_n883), .B2(new_n884), .ZN(G145));
  XNOR2_X1  g460(.A(G162), .B(G160), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n777), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n818), .B(new_n842), .Z(new_n888));
  AND2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n636), .A2(G130), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n478), .A2(G142), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n896), .B(new_n897), .C1(G118), .C2(new_n461), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n892), .A2(new_n893), .A3(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n743), .B(new_n899), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n788), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n511), .B(new_n642), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n891), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n891), .A2(new_n903), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g483(.A(G305), .B(G166), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n603), .B(G288), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT100), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n914), .B(KEYINPUT101), .C1(KEYINPUT42), .C2(new_n911), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(KEYINPUT101), .B2(new_n914), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n613), .A2(G299), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n613), .A2(G299), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(KEYINPUT99), .A3(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n918), .A2(KEYINPUT99), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n917), .A2(new_n918), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n626), .B(new_n877), .ZN(new_n927));
  MUX2_X1   g502(.A(new_n926), .B(new_n921), .S(new_n927), .Z(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n916), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n916), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(G868), .B2(new_n866), .ZN(G295));
  OAI21_X1  g508(.A(new_n932), .B1(G868), .B2(new_n866), .ZN(G331));
  XNOR2_X1  g509(.A(G301), .B(G286), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n877), .B(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(new_n921), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n877), .A2(new_n935), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n938), .A2(KEYINPUT102), .ZN(new_n939));
  XNOR2_X1  g514(.A(G168), .B(G301), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n940), .A2(KEYINPUT103), .A3(new_n876), .A4(new_n875), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n877), .B2(new_n935), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n938), .A2(KEYINPUT102), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n939), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n937), .B1(new_n925), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n913), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(KEYINPUT104), .A3(new_n913), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n946), .A2(new_n921), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n924), .A2(new_n922), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n921), .A2(new_n922), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n953), .A2(new_n954), .A3(new_n936), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n912), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n950), .A2(new_n951), .A3(new_n956), .A4(new_n906), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n950), .A2(new_n951), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n947), .A2(new_n913), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n906), .A4(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n957), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n960), .A2(KEYINPUT44), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n961), .A2(KEYINPUT43), .A3(new_n906), .A4(new_n963), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n957), .A2(new_n962), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(G397));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n972));
  NOR2_X1   g547(.A1(G166), .A2(KEYINPUT74), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT74), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n974), .B(new_n526), .C1(new_n534), .C2(new_n536), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT55), .B(G8), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(G303), .A2(KEYINPUT108), .A3(KEYINPUT55), .A4(G8), .ZN(new_n979));
  OAI21_X1  g554(.A(G8), .B1(new_n973), .B2(new_n975), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND4_X1   g557(.A1(new_n972), .A2(new_n978), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n513), .A2(new_n984), .A3(new_n516), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT107), .B(G40), .Z(new_n987));
  NOR3_X1   g562(.A1(new_n465), .A2(new_n472), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n514), .B2(new_n515), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n986), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G2090), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n985), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n988), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1971), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n992), .A2(new_n993), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n983), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G2084), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n986), .A2(new_n1002), .A3(new_n988), .A4(new_n991), .ZN(new_n1003));
  INV_X1    g578(.A(new_n988), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n511), .A2(new_n984), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(new_n994), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n984), .A4(new_n516), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1966), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1003), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(G286), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n997), .A2(new_n998), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n986), .A2(new_n993), .A3(new_n988), .A4(new_n991), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n978), .A2(new_n979), .A3(new_n982), .A4(new_n972), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(G8), .A3(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1001), .A2(new_n1013), .A3(new_n1018), .A4(KEYINPUT63), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n594), .A2(G651), .ZN(new_n1020));
  INV_X1    g595(.A(G48), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1020), .B1(new_n1021), .B2(new_n539), .ZN(new_n1022));
  NOR2_X1   g597(.A1(KEYINPUT112), .A2(G86), .ZN(new_n1023));
  AND2_X1   g598(.A1(KEYINPUT112), .A2(G86), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n531), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(G1981), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n595), .A2(new_n703), .A3(new_n596), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT49), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT49), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n511), .A2(new_n984), .A3(new_n988), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT109), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1034), .A3(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G288), .A2(new_n716), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1039), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT109), .B(new_n1000), .C1(new_n989), .C2(new_n988), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1034), .B1(new_n1031), .B2(G8), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1037), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(G288), .B2(new_n716), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1043), .B(new_n1049), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1036), .A2(KEYINPUT111), .A3(new_n1043), .A4(new_n1049), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1019), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n513), .A2(new_n984), .A3(new_n516), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n990), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n998), .A2(new_n997), .B1(new_n1061), .B2(new_n993), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1058), .B1(new_n1062), .B2(new_n1000), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1016), .A2(G8), .A3(new_n1057), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1046), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT110), .B1(new_n1046), .B2(KEYINPUT52), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT114), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1065), .B(new_n1013), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1056), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1066), .A2(new_n716), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1027), .B1(new_n1078), .B2(G288), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1036), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1055), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1064), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT117), .B1(new_n1077), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1081), .A2(new_n1036), .B1(new_n1084), .B2(new_n1083), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1071), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1048), .A2(KEYINPUT114), .A3(new_n1054), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1075), .B1(new_n1093), .B2(new_n1013), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1088), .B(new_n1089), .C1(new_n1094), .C2(new_n1056), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n578), .A2(KEYINPUT119), .A3(new_n580), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT119), .B1(new_n578), .B2(new_n580), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n576), .A2(KEYINPUT120), .A3(new_n582), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT120), .B1(new_n576), .B2(new_n582), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1098), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT121), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1106), .A3(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT118), .B(G1956), .Z(new_n1109));
  NOR2_X1   g684(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n1059), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n995), .A2(new_n988), .A3(new_n996), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1108), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1105), .A2(new_n1111), .A3(new_n1107), .A4(new_n1113), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT61), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n986), .A2(new_n988), .A3(new_n991), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n811), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1031), .A2(KEYINPUT122), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n989), .B2(new_n988), .ZN(new_n1122));
  OR3_X1    g697(.A1(new_n1120), .A2(new_n1122), .A3(G2067), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n613), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1124), .A2(KEYINPUT60), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1117), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1124), .A2(new_n613), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1125), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT60), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1114), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1111), .A2(new_n1113), .A3(KEYINPUT123), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1108), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1004), .B1(new_n985), .B2(new_n994), .ZN(new_n1136));
  INV_X1    g711(.A(G1996), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n996), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT124), .B(new_n1139), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1138), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1144), .A2(KEYINPUT59), .A3(new_n561), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT59), .B1(new_n1144), .B2(new_n561), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1127), .A2(new_n1130), .A3(new_n1135), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1134), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1116), .B1(new_n1149), .B2(new_n1129), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1011), .A2(G8), .A3(G286), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1000), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(KEYINPUT125), .A3(G286), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT51), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(G286), .A2(G8), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1012), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1012), .A2(new_n1158), .A3(KEYINPUT51), .A4(new_n1160), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1157), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AND4_X1   g739(.A1(KEYINPUT53), .A2(new_n996), .A3(G40), .A4(new_n798), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n989), .A2(KEYINPUT106), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n989), .A2(KEYINPUT106), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(new_n994), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1168), .A3(G160), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT127), .Z(new_n1170));
  XNOR2_X1  g745(.A(G301), .B(KEYINPUT54), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1136), .A2(new_n798), .A3(new_n996), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT53), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1173), .A2(new_n1174), .B1(new_n1118), .B2(new_n807), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1008), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1172), .A2(new_n1175), .B1(new_n1171), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1151), .A2(new_n1164), .A3(new_n1093), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1164), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1157), .A2(new_n1162), .A3(KEYINPUT62), .A4(new_n1163), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1183), .A2(G171), .A3(new_n1093), .A4(new_n1177), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1087), .A2(new_n1095), .A3(new_n1179), .A4(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1168), .A2(new_n1004), .ZN(new_n1186));
  INV_X1    g761(.A(G2067), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n818), .B(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n788), .B(G1996), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n743), .A2(new_n746), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n743), .A2(new_n746), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(G1986), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1196), .B1(new_n1197), .B2(new_n603), .ZN(new_n1198));
  NOR2_X1   g773(.A1(G290), .A2(G1986), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1186), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1185), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT46), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1186), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1202), .B1(new_n1203), .B2(G1996), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1186), .B1(new_n1189), .B2(new_n788), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1186), .A2(KEYINPUT46), .A3(new_n1137), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  XOR2_X1   g782(.A(new_n1207), .B(KEYINPUT47), .Z(new_n1208));
  NAND2_X1  g783(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1209));
  OR2_X1    g784(.A1(new_n818), .A2(G2067), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1203), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1186), .A2(new_n1199), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT48), .Z(new_n1213));
  AOI21_X1  g788(.A(new_n1213), .B1(new_n1186), .B2(new_n1195), .ZN(new_n1214));
  NOR3_X1   g789(.A1(new_n1208), .A2(new_n1211), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1201), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g791(.A(G229), .ZN(new_n1218));
  NAND4_X1  g792(.A1(new_n967), .A2(G319), .A3(new_n1218), .A4(new_n969), .ZN(new_n1219));
  NAND3_X1  g793(.A1(new_n907), .A2(new_n668), .A3(new_n685), .ZN(new_n1220));
  NOR2_X1   g794(.A1(new_n1219), .A2(new_n1220), .ZN(G308));
  AND2_X1   g795(.A1(new_n967), .A2(new_n969), .ZN(new_n1222));
  INV_X1    g796(.A(new_n1220), .ZN(new_n1223));
  NAND4_X1  g797(.A1(new_n1222), .A2(G319), .A3(new_n1223), .A4(new_n1218), .ZN(G225));
endmodule


