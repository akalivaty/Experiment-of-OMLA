

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  NAND2_X1 U322 ( .A1(n473), .A2(n472), .ZN(n483) );
  XOR2_X1 U323 ( .A(n446), .B(n329), .Z(n471) );
  XOR2_X1 U324 ( .A(n371), .B(n346), .Z(n290) );
  XOR2_X1 U325 ( .A(G120GAT), .B(KEYINPUT0), .Z(n291) );
  XOR2_X1 U326 ( .A(KEYINPUT25), .B(n463), .Z(n292) );
  XNOR2_X1 U327 ( .A(n372), .B(KEYINPUT79), .ZN(n373) );
  XNOR2_X1 U328 ( .A(n374), .B(n373), .ZN(n377) );
  INV_X1 U329 ( .A(KEYINPUT55), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U331 ( .A(KEYINPUT100), .B(KEYINPUT37), .ZN(n485) );
  XNOR2_X1 U332 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U333 ( .A(n486), .B(n485), .ZN(n513) );
  XNOR2_X1 U334 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n456) );
  XNOR2_X1 U335 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n296) );
  XOR2_X1 U337 ( .A(G29GAT), .B(G43GAT), .Z(n294) );
  XNOR2_X1 U338 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n403) );
  XOR2_X1 U340 ( .A(G36GAT), .B(G190GAT), .Z(n434) );
  XNOR2_X1 U341 ( .A(n403), .B(n434), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n302) );
  XOR2_X1 U343 ( .A(G162GAT), .B(KEYINPUT74), .Z(n298) );
  XNOR2_X1 U344 ( .A(G50GAT), .B(G218GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n359) );
  XOR2_X1 U346 ( .A(n359), .B(G134GAT), .Z(n300) );
  NAND2_X1 U347 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U349 ( .A(n302), .B(n301), .Z(n311) );
  XOR2_X1 U350 ( .A(KEYINPUT73), .B(G92GAT), .Z(n304) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(G85GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U353 ( .A(G106GAT), .B(n305), .Z(n399) );
  INV_X1 U354 ( .A(n399), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n307) );
  XNOR2_X1 U356 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U358 ( .A(n309), .B(n308), .Z(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n549) );
  XNOR2_X1 U360 ( .A(KEYINPUT78), .B(n549), .ZN(n534) );
  XOR2_X1 U361 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n313) );
  XNOR2_X1 U362 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(n314), .ZN(n446) );
  XOR2_X1 U365 ( .A(G176GAT), .B(G99GAT), .Z(n316) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(G190GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U368 ( .A(G183GAT), .B(KEYINPUT81), .Z(n318) );
  XNOR2_X1 U369 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n320), .B(n319), .Z(n328) );
  XOR2_X1 U372 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n322) );
  XNOR2_X1 U373 ( .A(G71GAT), .B(KEYINPUT83), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U375 ( .A(G15GAT), .B(G127GAT), .Z(n371) );
  XNOR2_X1 U376 ( .A(G113GAT), .B(G134GAT), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n291), .B(n323), .ZN(n346) );
  NAND2_X1 U378 ( .A1(G227GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n290), .B(n324), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n329) );
  NAND2_X1 U382 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XOR2_X1 U383 ( .A(G148GAT), .B(G155GAT), .Z(n331) );
  XNOR2_X1 U384 ( .A(G29GAT), .B(G127GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n333) );
  XOR2_X1 U386 ( .A(G162GAT), .B(G85GAT), .Z(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n352) );
  XOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT92), .Z(n337) );
  XNOR2_X1 U390 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n350) );
  XOR2_X1 U392 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n339) );
  XNOR2_X1 U393 ( .A(KEYINPUT1), .B(KEYINPUT95), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U395 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n341) );
  XNOR2_X1 U396 ( .A(KEYINPUT4), .B(KEYINPUT94), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U398 ( .A(n343), .B(n342), .Z(n348) );
  XOR2_X1 U399 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n345) );
  XNOR2_X1 U400 ( .A(G141GAT), .B(KEYINPUT88), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n358) );
  XNOR2_X1 U402 ( .A(n346), .B(n358), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U404 ( .A(n350), .B(n349), .Z(n351) );
  XOR2_X1 U405 ( .A(n352), .B(n351), .Z(n465) );
  XOR2_X1 U406 ( .A(G211GAT), .B(KEYINPUT22), .Z(n354) );
  XNOR2_X1 U407 ( .A(G106GAT), .B(KEYINPUT23), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n367) );
  XOR2_X1 U409 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n356) );
  NAND2_X1 U410 ( .A1(G228GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U412 ( .A(n357), .B(KEYINPUT87), .Z(n361) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n363) );
  XNOR2_X1 U415 ( .A(G78GAT), .B(G204GAT), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n362), .B(G148GAT), .ZN(n394) );
  XOR2_X1 U417 ( .A(n363), .B(n394), .Z(n365) );
  XOR2_X1 U418 ( .A(G22GAT), .B(G155GAT), .Z(n383) );
  XOR2_X1 U419 ( .A(G197GAT), .B(KEYINPUT21), .Z(n443) );
  XNOR2_X1 U420 ( .A(n383), .B(n443), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U422 ( .A(n367), .B(n366), .Z(n469) );
  NAND2_X1 U423 ( .A1(n465), .A2(n469), .ZN(n450) );
  XOR2_X1 U424 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n369) );
  XNOR2_X1 U425 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n387) );
  XNOR2_X1 U427 ( .A(G71GAT), .B(G57GAT), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n370), .B(KEYINPUT13), .ZN(n390) );
  XNOR2_X1 U429 ( .A(n390), .B(n371), .ZN(n374) );
  AND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(G8GAT), .B(G183GAT), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n375), .B(G211GAT), .ZN(n435) );
  XOR2_X1 U433 ( .A(n435), .B(KEYINPUT15), .Z(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n380) );
  INV_X1 U435 ( .A(n380), .ZN(n378) );
  NAND2_X1 U436 ( .A1(n378), .A2(G78GAT), .ZN(n382) );
  INV_X1 U437 ( .A(G78GAT), .ZN(n379) );
  NAND2_X1 U438 ( .A1(n380), .A2(n379), .ZN(n381) );
  NAND2_X1 U439 ( .A1(n382), .A2(n381), .ZN(n385) );
  XNOR2_X1 U440 ( .A(G1GAT), .B(n383), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U442 ( .A(n387), .B(n386), .Z(n577) );
  XOR2_X1 U443 ( .A(KEYINPUT112), .B(n577), .Z(n560) );
  NOR2_X1 U444 ( .A1(n549), .A2(n560), .ZN(n424) );
  XOR2_X1 U445 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n422) );
  XOR2_X1 U446 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n389) );
  XNOR2_X1 U447 ( .A(G120GAT), .B(KEYINPUT72), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n398) );
  XOR2_X1 U449 ( .A(G176GAT), .B(G64GAT), .Z(n442) );
  XOR2_X1 U450 ( .A(n442), .B(n390), .Z(n392) );
  NAND2_X1 U451 ( .A1(G230GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U453 ( .A(n393), .B(KEYINPUT71), .Z(n396) );
  XNOR2_X1 U454 ( .A(n394), .B(KEYINPUT31), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U456 ( .A(n398), .B(n397), .Z(n400) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n574) );
  XNOR2_X1 U458 ( .A(KEYINPUT41), .B(n574), .ZN(n542) );
  XOR2_X1 U459 ( .A(G36GAT), .B(G50GAT), .Z(n402) );
  NAND2_X1 U460 ( .A1(G229GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U462 ( .A(n404), .B(n403), .Z(n412) );
  XOR2_X1 U463 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n406) );
  XNOR2_X1 U464 ( .A(KEYINPUT67), .B(KEYINPUT70), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U466 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n408) );
  XNOR2_X1 U467 ( .A(KEYINPUT29), .B(KEYINPUT65), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n420) );
  XOR2_X1 U471 ( .A(G8GAT), .B(G1GAT), .Z(n414) );
  XNOR2_X1 U472 ( .A(G197GAT), .B(G141GAT), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U474 ( .A(G22GAT), .B(G15GAT), .Z(n416) );
  XNOR2_X1 U475 ( .A(G169GAT), .B(G113GAT), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U477 ( .A(n418), .B(n417), .Z(n419) );
  XOR2_X1 U478 ( .A(n420), .B(n419), .Z(n568) );
  INV_X1 U479 ( .A(n568), .ZN(n552) );
  NAND2_X1 U480 ( .A1(n542), .A2(n552), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  NAND2_X1 U482 ( .A1(n424), .A2(n423), .ZN(n425) );
  XNOR2_X1 U483 ( .A(KEYINPUT47), .B(n425), .ZN(n432) );
  INV_X1 U484 ( .A(n574), .ZN(n430) );
  XOR2_X1 U485 ( .A(KEYINPUT36), .B(n534), .Z(n581) );
  NOR2_X1 U486 ( .A1(n577), .A2(n581), .ZN(n427) );
  XNOR2_X1 U487 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  NAND2_X1 U489 ( .A1(n428), .A2(n568), .ZN(n429) );
  NOR2_X1 U490 ( .A1(n430), .A2(n429), .ZN(n431) );
  NOR2_X1 U491 ( .A1(n432), .A2(n431), .ZN(n433) );
  XNOR2_X1 U492 ( .A(KEYINPUT48), .B(n433), .ZN(n539) );
  XOR2_X1 U493 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U494 ( .A1(G226GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U496 ( .A(KEYINPUT96), .B(G92GAT), .Z(n439) );
  XNOR2_X1 U497 ( .A(G218GAT), .B(G204GAT), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U499 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n460) );
  NOR2_X1 U503 ( .A1(n539), .A2(n460), .ZN(n449) );
  INV_X1 U504 ( .A(KEYINPUT54), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(n564) );
  NOR2_X1 U506 ( .A1(n450), .A2(n564), .ZN(n454) );
  XNOR2_X1 U507 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n452) );
  NOR2_X1 U508 ( .A1(n471), .A2(n455), .ZN(n561) );
  NAND2_X1 U509 ( .A1(n534), .A2(n561), .ZN(n457) );
  INV_X1 U510 ( .A(n465), .ZN(n565) );
  NAND2_X1 U511 ( .A1(n552), .A2(n574), .ZN(n487) );
  NOR2_X1 U512 ( .A1(n577), .A2(n534), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT16), .ZN(n474) );
  INV_X1 U514 ( .A(n471), .ZN(n525) );
  NOR2_X1 U515 ( .A1(n469), .A2(n525), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(KEYINPUT26), .ZN(n566) );
  INV_X1 U517 ( .A(n460), .ZN(n515) );
  XNOR2_X1 U518 ( .A(n515), .B(KEYINPUT27), .ZN(n467) );
  NAND2_X1 U519 ( .A1(n566), .A2(n467), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n515), .A2(n525), .ZN(n461) );
  NAND2_X1 U521 ( .A1(n461), .A2(n469), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT98), .ZN(n463) );
  NAND2_X1 U523 ( .A1(n464), .A2(n292), .ZN(n466) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n473) );
  NAND2_X1 U525 ( .A1(n467), .A2(n565), .ZN(n468) );
  XOR2_X1 U526 ( .A(KEYINPUT97), .B(n468), .Z(n538) );
  XOR2_X1 U527 ( .A(n469), .B(KEYINPUT64), .Z(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT28), .B(n470), .ZN(n519) );
  NOR2_X1 U529 ( .A1(n538), .A2(n519), .ZN(n524) );
  NAND2_X1 U530 ( .A1(n524), .A2(n471), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n474), .A2(n483), .ZN(n501) );
  NOR2_X1 U532 ( .A1(n487), .A2(n501), .ZN(n481) );
  NAND2_X1 U533 ( .A1(n565), .A2(n481), .ZN(n475) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(n475), .ZN(n476) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U536 ( .A1(n515), .A2(n481), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n479) );
  NAND2_X1 U539 ( .A1(n481), .A2(n525), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U541 ( .A(G15GAT), .B(n480), .Z(G1326GAT) );
  NAND2_X1 U542 ( .A1(n519), .A2(n481), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT39), .Z(n491) );
  NAND2_X1 U545 ( .A1(n577), .A2(n483), .ZN(n484) );
  NOR2_X1 U546 ( .A1(n581), .A2(n484), .ZN(n486) );
  OR2_X1 U547 ( .A1(n513), .A2(n487), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U549 ( .A(KEYINPUT38), .B(n489), .ZN(n497) );
  NAND2_X1 U550 ( .A1(n565), .A2(n497), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n497), .A2(n515), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n497), .A2(n525), .ZN(n495) );
  XOR2_X1 U556 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  NAND2_X1 U559 ( .A1(n497), .A2(n519), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(KEYINPUT104), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n504) );
  XOR2_X1 U563 ( .A(n542), .B(KEYINPUT105), .Z(n557) );
  NAND2_X1 U564 ( .A1(n557), .A2(n568), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(KEYINPUT106), .ZN(n512) );
  NOR2_X1 U566 ( .A1(n512), .A2(n501), .ZN(n502) );
  XOR2_X1 U567 ( .A(KEYINPUT107), .B(n502), .Z(n509) );
  NAND2_X1 U568 ( .A1(n509), .A2(n565), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n505), .Z(G1332GAT) );
  NAND2_X1 U571 ( .A1(n515), .A2(n509), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT109), .Z(n508) );
  NAND2_X1 U574 ( .A1(n509), .A2(n525), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U577 ( .A1(n509), .A2(n519), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n520) );
  NAND2_X1 U580 ( .A1(n565), .A2(n520), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n515), .A2(n520), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(KEYINPUT110), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n525), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n522) );
  NAND2_X1 U588 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U592 ( .A1(n539), .A2(n526), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n552), .A2(n535), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U596 ( .A1(n535), .A2(n557), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n533) );
  XOR2_X1 U599 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n531) );
  NAND2_X1 U600 ( .A1(n535), .A2(n560), .ZN(n530) );
  XNOR2_X1 U601 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U604 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U607 ( .A1(n540), .A2(n566), .ZN(n547) );
  NOR2_X1 U608 ( .A1(n568), .A2(n547), .ZN(n541) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n541), .Z(G1344GAT) );
  XOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT117), .Z(n544) );
  INV_X1 U611 ( .A(n547), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n550), .A2(n542), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U614 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  OR2_X1 U616 ( .A1(n577), .A2(n547), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n548), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n552), .A2(n561), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n555) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(n556), .Z(n559) );
  NAND2_X1 U626 ( .A1(n557), .A2(n561), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G183GAT), .B(n563), .ZN(G1350GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n580) );
  NOR2_X1 U633 ( .A1(n568), .A2(n580), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT60), .B(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n580), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n580), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(G218GAT), .B(n584), .Z(G1355GAT) );
endmodule

