//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT80), .ZN(new_n190));
  INV_X1    g004(.A(G227), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n190), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT81), .A3(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT3), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(G104), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n210), .A2(new_n204), .A3(KEYINPUT81), .A4(G104), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n208), .A3(new_n209), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G107), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n214), .B2(new_n207), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n219), .A3(G143), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n221), .B2(G146), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n220), .A2(new_n222), .B1(G128), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n212), .B(new_n215), .C1(new_n225), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT10), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n221), .A2(G146), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(G146), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(G143), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n233), .B2(G143), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n236), .B2(new_n223), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n229), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n212), .A2(new_n215), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT84), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n223), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n217), .A2(new_n219), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n231), .B1(new_n243), .B2(new_n221), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n238), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n245), .A2(new_n240), .A3(KEYINPUT84), .A4(KEYINPUT10), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n230), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n206), .A2(new_n211), .A3(new_n208), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT82), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n206), .A2(new_n208), .A3(new_n252), .A4(new_n211), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n250), .A2(new_n251), .A3(G101), .A4(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n220), .A2(new_n222), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n255), .A2(new_n256), .B1(new_n234), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n250), .A2(G101), .A3(new_n253), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n261), .A2(KEYINPUT83), .A3(new_n262), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n260), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n203), .B1(new_n248), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT87), .ZN(new_n269));
  OR2_X1    g083(.A1(new_n225), .A2(new_n227), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT10), .B1(new_n270), .B2(new_n240), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n245), .A2(new_n240), .A3(KEYINPUT10), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n271), .B1(new_n274), .B2(new_n246), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n254), .A2(new_n259), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n261), .A2(KEYINPUT83), .A3(new_n262), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT83), .B1(new_n261), .B2(new_n262), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT87), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n203), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n269), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n275), .A2(new_n279), .A3(new_n202), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n193), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n212), .A2(new_n215), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n237), .A2(new_n238), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT85), .A3(new_n228), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n237), .A2(new_n286), .A3(new_n289), .A4(new_n238), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n288), .A2(KEYINPUT12), .A3(new_n203), .A4(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT86), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n203), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n295), .A2(KEYINPUT86), .A3(KEYINPUT12), .A4(new_n288), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT12), .ZN(new_n297));
  INV_X1    g111(.A(new_n288), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(new_n294), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n300), .A2(new_n284), .A3(new_n193), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n187), .B(new_n188), .C1(new_n285), .C2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n193), .B1(new_n300), .B2(new_n284), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n284), .A2(new_n193), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n283), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G469), .B1(new_n305), .B2(G902), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT9), .B(G234), .ZN(new_n308));
  OAI21_X1  g122(.A(G221), .B1(new_n308), .B2(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(G237), .A2(G953), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(G143), .A3(G214), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(G143), .B1(new_n311), .B2(G214), .ZN(new_n314));
  OAI21_X1  g128(.A(G131), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT17), .ZN(new_n316));
  INV_X1    g130(.A(G237), .ZN(new_n317));
  INV_X1    g131(.A(G953), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G214), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n221), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n201), .A3(new_n312), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n315), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G125), .B(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT16), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(G125), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT74), .B1(new_n329), .B2(KEYINPUT16), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n216), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n324), .A2(G146), .A3(new_n328), .A4(new_n330), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT17), .B(G131), .C1(new_n313), .C2(new_n314), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n322), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n336), .B1(new_n243), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n233), .A2(new_n323), .A3(KEYINPUT77), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(G146), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT18), .A2(G131), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n313), .B2(new_n314), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n320), .A2(new_n312), .A3(new_n345), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(G113), .B(G122), .Z(new_n351));
  XOR2_X1   g165(.A(KEYINPUT91), .B(G104), .Z(new_n352));
  XOR2_X1   g166(.A(new_n351), .B(new_n352), .Z(new_n353));
  AND3_X1   g167(.A1(new_n335), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n335), .B2(new_n350), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n188), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G475), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT20), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n323), .A2(KEYINPUT19), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n329), .A2(new_n338), .A3(KEYINPUT19), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n333), .B1(new_n361), .B2(new_n243), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n315), .A2(new_n321), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n340), .A2(new_n341), .B1(G146), .B2(new_n339), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n347), .A2(new_n348), .ZN(new_n365));
  OAI22_X1  g179(.A1(new_n362), .A2(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n353), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n335), .A2(new_n350), .A3(new_n353), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G475), .A2(G902), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n358), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n371), .ZN(new_n373));
  AOI211_X1 g187(.A(KEYINPUT20), .B(new_n373), .C1(new_n368), .C2(new_n369), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n357), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT92), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT92), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n357), .B(new_n377), .C1(new_n372), .C2(new_n374), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G478), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(KEYINPUT15), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n223), .A2(G143), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n221), .A2(KEYINPUT13), .A3(G128), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n223), .B2(G143), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n382), .B(new_n383), .C1(new_n385), .C2(KEYINPUT94), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n385), .A2(KEYINPUT94), .ZN(new_n387));
  OAI21_X1  g201(.A(G134), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n221), .A2(G128), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n382), .A3(new_n195), .ZN(new_n390));
  INV_X1    g204(.A(G116), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G122), .ZN(new_n392));
  INV_X1    g206(.A(G122), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G116), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n392), .A2(new_n394), .A3(new_n204), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n204), .B1(new_n392), .B2(new_n394), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT93), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n394), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G107), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT93), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n392), .A2(new_n394), .A3(new_n204), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n388), .A2(new_n390), .A3(new_n397), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n389), .A2(new_n382), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G134), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n390), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n391), .A2(KEYINPUT14), .A3(G122), .ZN(new_n407));
  OAI211_X1 g221(.A(G107), .B(new_n407), .C1(new_n398), .C2(KEYINPUT14), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n408), .A3(new_n401), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G217), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n308), .A2(new_n411), .A3(G953), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n403), .A2(new_n409), .A3(new_n412), .ZN(new_n415));
  AOI21_X1  g229(.A(G902), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT95), .B1(new_n416), .B2(KEYINPUT96), .ZN(new_n417));
  INV_X1    g231(.A(new_n415), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n412), .B1(new_n403), .B2(new_n409), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT95), .B(new_n188), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n381), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n414), .A2(new_n415), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT96), .A3(new_n188), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT95), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n381), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(G234), .A2(G237), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(G952), .A3(new_n318), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(G898), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(G902), .A3(G953), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n436), .B(KEYINPUT97), .Z(new_n437));
  AND3_X1   g251(.A1(new_n379), .A2(new_n430), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n337), .B(new_n238), .C1(new_n242), .C2(new_n244), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n440), .A2(KEYINPUT88), .ZN(new_n441));
  OAI211_X1 g255(.A(KEYINPUT88), .B(new_n440), .C1(new_n259), .C2(new_n337), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n318), .A2(G224), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n441), .B2(new_n442), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT7), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT8), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n452));
  XOR2_X1   g266(.A(G116), .B(G119), .Z(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT2), .B(G113), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT2), .B(G113), .Z(new_n456));
  XNOR2_X1  g270(.A(G116), .B(G119), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(KEYINPUT66), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(KEYINPUT5), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n391), .A2(KEYINPUT5), .A3(G119), .ZN(new_n460));
  INV_X1    g274(.A(G113), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n455), .A2(new_n458), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(KEYINPUT89), .A3(new_n240), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n240), .B2(new_n463), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT89), .B1(new_n463), .B2(new_n240), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n451), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n441), .A2(new_n442), .A3(new_n446), .A4(new_n443), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n449), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n240), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n277), .A2(new_n278), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n455), .A2(new_n458), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n457), .B1(new_n456), .B2(KEYINPUT65), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n454), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n254), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n471), .B(new_n450), .C1(new_n472), .C2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n470), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n450), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n479), .B1(new_n265), .B2(new_n266), .ZN(new_n483));
  INV_X1    g297(.A(new_n471), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n480), .A3(KEYINPUT6), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n487), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n444), .A2(new_n445), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n481), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n491), .B(KEYINPUT90), .Z(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n481), .B2(new_n490), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n438), .B(new_n439), .C1(new_n492), .C2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n310), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n318), .A2(G221), .A3(G234), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT79), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT22), .B(G137), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n499), .B(new_n500), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n223), .A2(G119), .ZN(new_n503));
  INV_X1    g317(.A(G119), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G128), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT72), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT72), .ZN(new_n507));
  INV_X1    g321(.A(G110), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT24), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT24), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G110), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n509), .B2(new_n511), .ZN(new_n514));
  OAI22_X1  g328(.A1(new_n506), .A2(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT75), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n503), .A2(new_n505), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT72), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n510), .A2(G110), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n508), .A2(KEYINPUT24), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT73), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(new_n528), .A3(KEYINPUT75), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n223), .A2(KEYINPUT23), .A3(G119), .ZN(new_n530));
  INV_X1    g344(.A(new_n503), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n505), .B(new_n530), .C1(new_n531), .C2(KEYINPUT23), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(G110), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n517), .A2(new_n518), .A3(new_n529), .A4(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n342), .A2(new_n333), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n521), .A2(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n533), .B1(new_n538), .B2(KEYINPUT75), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n518), .B1(new_n539), .B2(new_n517), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT78), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n529), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n538), .A2(KEYINPUT75), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT76), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT78), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n535), .A4(new_n536), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n523), .A2(new_n528), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(G110), .B2(new_n532), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n332), .A2(new_n333), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n502), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n551), .ZN(new_n553));
  AOI211_X1 g367(.A(new_n553), .B(new_n501), .C1(new_n541), .C2(new_n546), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n411), .B1(G234), .B2(new_n188), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n555), .A2(G902), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n188), .B1(new_n552), .B2(new_n554), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT25), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT25), .B(new_n188), .C1(new_n552), .C2(new_n554), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n557), .B1(new_n562), .B2(new_n556), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n564));
  NAND2_X1  g378(.A1(new_n311), .A2(G210), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT26), .B(G101), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n455), .A2(new_n458), .B1(new_n474), .B2(new_n476), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n234), .A2(new_n258), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n220), .A2(new_n256), .A3(new_n222), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(new_n202), .ZN(new_n574));
  INV_X1    g388(.A(new_n199), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n195), .A2(G137), .ZN(new_n576));
  OAI21_X1  g390(.A(G131), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n196), .A2(new_n198), .A3(new_n201), .A4(new_n199), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n237), .B2(new_n238), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT30), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n579), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n245), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n200), .A2(G131), .ZN(new_n584));
  INV_X1    g398(.A(new_n578), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n571), .B(new_n572), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT30), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n570), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n583), .A2(new_n586), .A3(new_n570), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n569), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT29), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n570), .B1(new_n583), .B2(new_n586), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT28), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n583), .A2(new_n586), .A3(new_n570), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT28), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n594), .A2(new_n597), .A3(new_n568), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n591), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT69), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT69), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n591), .A2(new_n598), .A3(new_n601), .A4(new_n592), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n597), .A2(KEYINPUT71), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT71), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n595), .A2(new_n606), .A3(new_n596), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g422(.A(KEYINPUT70), .B(KEYINPUT28), .C1(new_n590), .C2(new_n593), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n569), .A2(new_n592), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n604), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n600), .A2(new_n188), .A3(new_n602), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT32), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n583), .A2(new_n587), .A3(new_n586), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n587), .B1(new_n583), .B2(new_n586), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n478), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(new_n595), .A3(new_n568), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT31), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n617), .A2(KEYINPUT31), .A3(new_n595), .A4(new_n568), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n594), .A2(new_n597), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n620), .A2(new_n621), .B1(new_n622), .B2(new_n569), .ZN(new_n623));
  NOR2_X1   g437(.A1(G472), .A2(G902), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT68), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n614), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n620), .A2(new_n621), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n569), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n625), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(KEYINPUT32), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n613), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n563), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n497), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G101), .ZN(G3));
  AOI21_X1  g449(.A(new_n491), .B1(new_n481), .B2(new_n490), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n439), .B(new_n437), .C1(new_n492), .C2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n423), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT33), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n423), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n380), .A2(G902), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(G478), .B2(new_n416), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n376), .A3(new_n378), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n309), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n302), .B2(new_n306), .ZN(new_n649));
  INV_X1    g463(.A(new_n556), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n560), .B2(new_n561), .ZN(new_n651));
  AOI21_X1  g465(.A(G902), .B1(new_n627), .B2(new_n628), .ZN(new_n652));
  INV_X1    g466(.A(G472), .ZN(new_n653));
  OAI22_X1  g467(.A1(new_n652), .A2(new_n653), .B1(new_n623), .B2(new_n625), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n651), .A2(new_n654), .A3(new_n557), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n647), .A2(new_n649), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT99), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT34), .B(G104), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  INV_X1    g473(.A(new_n375), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n429), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n637), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n649), .A3(new_n655), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT100), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NAND2_X1  g480(.A1(new_n562), .A2(new_n556), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n547), .A2(new_n551), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n502), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n556), .A2(G902), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n654), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n497), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  AND2_X1   g490(.A1(new_n631), .A2(new_n626), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n667), .A2(new_n672), .B1(new_n677), .B2(new_n613), .ZN(new_n678));
  INV_X1    g492(.A(new_n439), .ZN(new_n679));
  INV_X1    g493(.A(new_n491), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n489), .A2(new_n447), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n480), .A3(new_n468), .A4(new_n467), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n188), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n481), .A2(new_n490), .A3(new_n491), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n679), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n661), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n435), .A2(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n432), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n678), .A2(new_n649), .A3(new_n687), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  XNOR2_X1  g508(.A(new_n690), .B(KEYINPUT39), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n649), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT40), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n492), .A2(new_n495), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n569), .B1(new_n590), .B2(new_n593), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT102), .ZN(new_n703));
  INV_X1    g517(.A(new_n618), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n188), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n677), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n667), .A2(new_n672), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n429), .A2(new_n376), .A3(new_n378), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n708), .A2(new_n679), .A3(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n697), .A2(new_n701), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT103), .B(G143), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G45));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n439), .B1(new_n492), .B2(new_n636), .ZN(new_n715));
  INV_X1    g529(.A(new_n690), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n646), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n714), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n646), .A2(new_n716), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n687), .A2(KEYINPUT104), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n678), .A2(new_n718), .A3(new_n649), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  AOI21_X1  g536(.A(new_n281), .B1(new_n280), .B2(new_n203), .ZN(new_n723));
  AOI211_X1 g537(.A(KEYINPUT87), .B(new_n202), .C1(new_n275), .C2(new_n279), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n284), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n193), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n301), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(G469), .B1(new_n727), .B2(G902), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n728), .A2(new_n302), .A3(new_n309), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n647), .A2(new_n729), .A3(new_n632), .A4(new_n563), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND4_X1  g546(.A1(new_n662), .A2(new_n729), .A3(new_n632), .A4(new_n563), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  AND3_X1   g548(.A1(new_n708), .A2(new_n632), .A3(new_n438), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n729), .B2(new_n687), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n728), .A2(new_n302), .A3(new_n309), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n738), .A2(KEYINPUT105), .A3(new_n715), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n735), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  NAND3_X1  g555(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n569), .A2(new_n742), .B1(new_n620), .B2(new_n621), .ZN(new_n743));
  OAI22_X1  g557(.A1(new_n652), .A2(new_n653), .B1(new_n743), .B2(new_n625), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n651), .A2(new_n744), .A3(new_n557), .ZN(new_n745));
  AOI211_X1 g559(.A(new_n679), .B(new_n709), .C1(new_n685), .C2(new_n686), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n729), .A2(new_n745), .A3(new_n746), .A4(new_n437), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n557), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n742), .A2(new_n569), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n625), .B1(new_n751), .B2(new_n627), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n629), .A2(new_n188), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n752), .B1(new_n753), .B2(G472), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n667), .A2(new_n750), .A3(new_n437), .A4(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(KEYINPUT106), .A3(new_n729), .A4(new_n746), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  INV_X1    g573(.A(new_n672), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n719), .B(new_n754), .C1(new_n651), .C2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n737), .B2(new_n739), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  NOR3_X1   g578(.A1(new_n492), .A2(new_n495), .A3(new_n679), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n646), .A2(new_n766), .A3(new_n716), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n649), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n631), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n629), .A2(KEYINPUT107), .A3(KEYINPUT32), .A4(new_n630), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n770), .A2(new_n613), .A3(new_n626), .A4(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n772), .A2(new_n773), .A3(new_n563), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n772), .B2(new_n563), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n768), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n649), .A2(new_n632), .A3(new_n563), .A4(new_n765), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n766), .B1(new_n777), .B2(new_n717), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  NOR2_X1   g594(.A1(new_n777), .A2(new_n691), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n195), .ZN(G36));
  NAND2_X1  g596(.A1(new_n379), .A2(new_n645), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT43), .Z(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n654), .A3(new_n708), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n305), .A2(KEYINPUT45), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n305), .A2(KEYINPUT45), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(G469), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(G469), .A2(G902), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT46), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n302), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n790), .A2(KEYINPUT46), .A3(new_n791), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n648), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n765), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n785), .B2(new_n786), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n787), .A2(new_n796), .A3(new_n695), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  AND2_X1   g614(.A1(new_n796), .A2(KEYINPUT47), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n796), .A2(KEYINPUT47), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n797), .A2(new_n563), .A3(new_n632), .A4(new_n717), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT109), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n804), .A2(KEYINPUT109), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NOR3_X1   g625(.A1(new_n701), .A2(new_n707), .A3(new_n783), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n563), .A2(new_n309), .A3(new_n439), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT110), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n728), .A2(new_n302), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT49), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n755), .A2(new_n738), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT106), .B1(new_n818), .B2(new_n746), .ZN(new_n819));
  INV_X1    g633(.A(new_n709), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n687), .A2(new_n820), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n755), .A2(new_n821), .A3(new_n738), .A4(new_n748), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n740), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n497), .B1(new_n633), .B2(new_n673), .ZN(new_n824));
  INV_X1    g638(.A(new_n437), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n698), .A2(new_n679), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n379), .A2(new_n429), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n379), .A2(KEYINPUT111), .A3(new_n429), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n646), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n826), .A2(new_n655), .A3(new_n649), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n824), .A2(new_n730), .A3(new_n733), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n823), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n708), .A2(new_n716), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n649), .A3(new_n707), .A4(new_n746), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n763), .A2(new_n693), .A3(new_n721), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n721), .A2(new_n693), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n840), .A3(new_n763), .A4(new_n836), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n649), .A2(new_n765), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n429), .A2(new_n375), .A3(new_n716), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n632), .B(new_n843), .C1(new_n651), .C2(new_n760), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n844), .B2(new_n761), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n781), .B(new_n845), .C1(new_n776), .C2(new_n778), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n834), .A2(new_n838), .A3(new_n841), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n730), .A2(new_n733), .A3(new_n832), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n758), .A3(new_n740), .A4(new_n824), .ZN(new_n851));
  INV_X1    g665(.A(new_n781), .ZN(new_n852));
  INV_X1    g666(.A(new_n845), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n779), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n841), .A4(new_n838), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n849), .A2(new_n856), .A3(KEYINPUT54), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT54), .B1(new_n849), .B2(new_n856), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n861));
  INV_X1    g675(.A(new_n563), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n729), .A2(new_n765), .ZN(new_n863));
  OR4_X1    g677(.A1(new_n862), .A2(new_n863), .A3(new_n432), .A4(new_n707), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n645), .B(new_n864), .C1(new_n376), .C2(new_n378), .ZN(new_n865));
  INV_X1    g679(.A(new_n432), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n784), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n863), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n708), .A3(new_n754), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT113), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n867), .A2(new_n862), .A3(new_n744), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n679), .A3(new_n700), .A4(new_n729), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT50), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n875), .A2(KEYINPUT112), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT112), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n815), .A2(new_n648), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n803), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n765), .A3(new_n872), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n861), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n864), .A2(new_n646), .ZN(new_n885));
  INV_X1    g699(.A(G952), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n885), .A2(new_n886), .A3(G953), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n774), .A2(new_n775), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n868), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT48), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n872), .B1(new_n739), .B2(new_n737), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n861), .B1(new_n875), .B2(new_n876), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n871), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n894), .B2(new_n882), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n860), .A2(new_n884), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(G952), .A2(G953), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n817), .B1(new_n896), .B2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n318), .A2(G952), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT114), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n486), .A2(new_n488), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n489), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n188), .B1(new_n849), .B2(new_n856), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(G210), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n905), .A2(new_n493), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n904), .A2(new_n907), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n901), .B(new_n908), .C1(new_n909), .C2(new_n910), .ZN(G51));
  XNOR2_X1  g725(.A(new_n727), .B(KEYINPUT116), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n791), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n860), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n790), .B(KEYINPUT117), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n905), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n899), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT118), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n905), .A2(new_n370), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n370), .B1(new_n905), .B2(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n899), .ZN(G60));
  NAND2_X1  g737(.A1(new_n849), .A2(new_n856), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n849), .A2(new_n856), .A3(KEYINPUT54), .ZN(new_n927));
  XNOR2_X1  g741(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n380), .A2(new_n188), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n640), .A2(new_n642), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n901), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n932), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n859), .A2(KEYINPUT120), .A3(new_n934), .A4(new_n930), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n926), .A2(new_n934), .A3(new_n927), .A4(new_n930), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n933), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n933), .A2(new_n935), .A3(new_n938), .A4(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT60), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n924), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n555), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n924), .A2(new_n670), .A3(new_n945), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n901), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n947), .A2(new_n900), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n954), .B2(new_n950), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G66));
  NAND2_X1  g770(.A1(new_n851), .A2(new_n318), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT123), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n318), .B1(new_n434), .B2(G224), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n902), .B1(G898), .B2(new_n318), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(G69));
  INV_X1    g776(.A(G900), .ZN(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n191), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT125), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n615), .A2(new_n616), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(new_n361), .ZN(new_n968));
  NAND2_X1  g782(.A1(G900), .A2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n839), .A2(new_n763), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n781), .B1(new_n776), .B2(new_n778), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n796), .A2(new_n695), .A3(new_n746), .A4(new_n888), .ZN(new_n973));
  AND4_X1   g787(.A1(new_n799), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n810), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n970), .B1(new_n976), .B2(new_n318), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n971), .A2(new_n711), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT62), .Z(new_n979));
  NAND4_X1  g793(.A1(new_n696), .A2(new_n633), .A3(new_n765), .A4(new_n831), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n799), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT124), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n810), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n968), .B1(new_n983), .B2(new_n318), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n966), .B1(new_n977), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n968), .B(new_n969), .C1(new_n975), .C2(G953), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n983), .A2(new_n318), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n986), .B(new_n965), .C1(new_n987), .C2(new_n968), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n985), .A2(new_n988), .ZN(G72));
  XNOR2_X1  g803(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n653), .A2(new_n188), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n983), .B2(new_n851), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n617), .A2(new_n595), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n993), .A2(new_n568), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n975), .B2(new_n851), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n994), .A2(new_n568), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT127), .Z(new_n998));
  AOI21_X1  g812(.A(new_n899), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n591), .A2(new_n618), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n924), .A2(new_n992), .A3(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n995), .A2(new_n999), .A3(new_n1001), .ZN(G57));
endmodule


