//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n451, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT67), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g025(.A(G2106), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n455), .A2(new_n451), .B1(new_n459), .B2(new_n456), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT69), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n463), .B1(new_n468), .B2(KEYINPUT70), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n466), .ZN(new_n475));
  NAND3_X1  g050(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  NAND2_X1  g053(.A1(G101), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n473), .A2(new_n480), .ZN(G160));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n464), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n477), .A2(new_n462), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n489));
  AND3_X1   g064(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT3), .B1(KEYINPUT71), .B2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n489), .B1(new_n492), .B2(new_n462), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n477), .A2(KEYINPUT72), .A3(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n488), .B1(G124), .B2(new_n495), .ZN(G162));
  OAI211_X1 g071(.A(KEYINPUT4), .B(G138), .C1(new_n490), .C2(new_n491), .ZN(new_n497));
  NAND2_X1  g072(.A1(G102), .A2(G2104), .ZN(new_n498));
  AOI21_X1  g073(.A(G2105), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G126), .B1(new_n490), .B2(new_n491), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(G114), .B2(G2104), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n462), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT4), .B1(new_n470), .B2(G138), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n499), .A2(new_n503), .A3(new_n504), .ZN(G164));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT73), .B(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n508), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n510), .A2(G50), .B1(G75), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n511), .A2(G62), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(new_n517), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n514), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n510), .A2(G89), .A3(new_n517), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT73), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n509), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g103(.A(G51), .B(G543), .C1(new_n528), .C2(new_n506), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n517), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n523), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND3_X1  g111(.A1(new_n510), .A2(G90), .A3(new_n517), .ZN(new_n537));
  OAI211_X1 g112(.A(G52), .B(G543), .C1(new_n528), .C2(new_n506), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n515), .B2(new_n516), .ZN(new_n540));
  AND2_X1   g115(.A1(G77), .A2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n511), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n537), .A2(new_n538), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND3_X1  g119(.A1(new_n510), .A2(G81), .A3(new_n517), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n510), .A2(G43), .A3(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n515), .B2(new_n516), .ZN(new_n548));
  AND2_X1   g123(.A1(G68), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n511), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND3_X1  g133(.A1(new_n510), .A2(G53), .A3(G543), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n524), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n510), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n510), .A2(G91), .A3(new_n517), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n561), .A2(new_n563), .A3(new_n564), .A4(new_n565), .ZN(G299));
  OAI221_X1 g141(.A(new_n518), .B1(new_n519), .B2(new_n520), .C1(new_n512), .C2(new_n513), .ZN(G303));
  NAND3_X1  g142(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n568), .B(new_n569), .C1(new_n519), .C2(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n517), .A2(G61), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n508), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT75), .B1(new_n577), .B2(new_n508), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n510), .A2(G86), .A3(new_n517), .ZN(new_n580));
  AND2_X1   g155(.A1(G48), .A2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n581), .B1(new_n528), .B2(new_n506), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(G305));
  NAND3_X1  g159(.A1(new_n510), .A2(G85), .A3(new_n517), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n510), .A2(G543), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT76), .B(G47), .Z(new_n588));
  OAI221_X1 g163(.A(new_n585), .B1(new_n508), .B2(new_n586), .C1(new_n587), .C2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  OAI211_X1 g165(.A(G54), .B(G543), .C1(new_n528), .C2(new_n506), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n515), .B2(new_n516), .ZN(new_n593));
  AND2_X1   g168(.A1(G79), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT77), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n591), .A2(new_n598), .A3(new_n595), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n510), .A2(G92), .A3(new_n517), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n510), .A2(KEYINPUT10), .A3(G92), .A4(new_n517), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n597), .A2(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n590), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n590), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n602), .A2(new_n603), .ZN(new_n613));
  INV_X1    g188(.A(new_n599), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n598), .B1(new_n591), .B2(new_n595), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT78), .B1(new_n616), .B2(G559), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n604), .A2(new_n618), .A3(new_n611), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n617), .A2(G868), .A3(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n552), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT11), .Z(G282));
  INV_X1    g199(.A(new_n623), .ZN(G323));
  NAND3_X1  g200(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G2100), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT79), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n495), .A2(G123), .ZN(new_n631));
  INV_X1    g206(.A(new_n486), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n464), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n632), .A2(G135), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  OAI211_X1 g213(.A(new_n630), .B(new_n638), .C1(G2100), .C2(new_n628), .ZN(G156));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT80), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT14), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n646), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n655), .A3(G14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n661), .B(KEYINPUT17), .Z(new_n665));
  INV_X1    g240(.A(new_n658), .ZN(new_n666));
  INV_X1    g241(.A(new_n659), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n662), .A3(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(new_n660), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n664), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT81), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(new_n684), .B(new_n683), .S(new_n676), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT82), .B(G1986), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G32), .ZN(new_n697));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT26), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n701));
  INV_X1    g276(.A(G141), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n700), .B(new_n701), .C1(new_n486), .C2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G129), .B2(new_n495), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n697), .B1(new_n704), .B2(new_n696), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT91), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT27), .B(G1996), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G21), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G168), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n706), .A2(new_n708), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n706), .A2(new_n708), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n709), .A2(G5), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G301), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G1961), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT95), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n715), .A2(new_n716), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n723));
  INV_X1    g298(.A(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G160), .B2(new_n696), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(G2084), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(KEYINPUT96), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n696), .A2(G26), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G128), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n493), .B2(new_n494), .ZN(new_n734));
  INV_X1    g309(.A(G140), .ZN(new_n735));
  NOR2_X1   g310(.A1(G104), .A2(G2105), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n486), .A2(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n696), .ZN(new_n740));
  INV_X1    g315(.A(G2067), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n728), .A2(KEYINPUT96), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n729), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n709), .A2(G19), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n552), .B2(new_n709), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(G1341), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n719), .B2(new_n718), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT25), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n470), .A2(G127), .ZN(new_n751));
  NAND2_X1  g326(.A1(G115), .A2(G2104), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n750), .B1(new_n753), .B2(G2105), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n632), .A2(G139), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n696), .A2(G33), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G11), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT94), .B(G28), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(new_n696), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n762), .B1(new_n764), .B2(new_n766), .C1(new_n637), .C2(new_n696), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n758), .B1(new_n757), .B2(new_n759), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n760), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n696), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n696), .ZN(new_n771));
  INV_X1    g346(.A(G2078), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n746), .A2(G1341), .B1(new_n727), .B2(G2084), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n748), .A2(new_n769), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n722), .A2(new_n744), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n709), .A2(G20), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n608), .B2(new_n709), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n696), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n696), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT29), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n780), .B1(G2090), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n709), .A2(G4), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n604), .B2(new_n709), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT88), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT89), .B(G1348), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n713), .A2(new_n714), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n783), .A2(G2090), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND3_X1   g367(.A1(new_n784), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n787), .A2(new_n788), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n776), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G23), .B(G288), .S(G16), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT33), .B(G1976), .Z(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G16), .A2(G22), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G166), .B2(G16), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n798), .B1(G1971), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n579), .A2(G16), .A3(new_n583), .ZN(new_n802));
  OR2_X1    g377(.A1(G6), .A2(G16), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT32), .B(G1981), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n800), .ZN(new_n807));
  INV_X1    g382(.A(G1971), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n807), .A2(new_n808), .B1(new_n796), .B2(new_n797), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n801), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT86), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n801), .A2(new_n806), .A3(new_n809), .A4(KEYINPUT86), .ZN(new_n813));
  AOI21_X1  g388(.A(KEYINPUT34), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(KEYINPUT34), .A3(new_n813), .ZN(new_n816));
  MUX2_X1   g391(.A(G24), .B(G290), .S(G16), .Z(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G1986), .Z(new_n818));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(KEYINPUT87), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n696), .A2(G25), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT83), .Z(new_n822));
  OR2_X1    g397(.A1(G95), .A2(G2105), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n823), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT85), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n632), .A2(G131), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT84), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n495), .B2(G119), .ZN(new_n828));
  INV_X1    g403(.A(G119), .ZN(new_n829));
  AOI211_X1 g404(.A(KEYINPUT84), .B(new_n829), .C1(new_n493), .C2(new_n494), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n825), .B(new_n826), .C1(new_n828), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n822), .B1(new_n831), .B2(G29), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT35), .B(G1991), .Z(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n820), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n815), .A2(new_n816), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n819), .A2(KEYINPUT87), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n795), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n815), .A2(new_n838), .A3(new_n816), .A4(new_n836), .ZN(new_n841));
  AOI21_X1  g416(.A(KEYINPUT97), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n836), .A2(new_n816), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n839), .B1(new_n843), .B2(new_n814), .ZN(new_n844));
  INV_X1    g419(.A(new_n795), .ZN(new_n845));
  AND4_X1   g420(.A1(KEYINPUT97), .A2(new_n844), .A3(new_n841), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n842), .A2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n840), .A2(new_n841), .ZN(G150));
  NAND3_X1  g423(.A1(new_n510), .A2(G93), .A3(new_n517), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n510), .A2(G55), .A3(G543), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n515), .B2(new_n516), .ZN(new_n852));
  AND2_X1   g427(.A1(G80), .A2(G543), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n511), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n551), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n551), .A2(new_n855), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT38), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n604), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n862), .A2(new_n863), .A3(G860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n855), .A2(G860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT37), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  OAI21_X1  g442(.A(G162), .B1(new_n480), .B2(new_n473), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n495), .A2(G124), .ZN(new_n869));
  INV_X1    g444(.A(new_n488), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G160), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n868), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n873), .B1(new_n868), .B2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n637), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n868), .A2(new_n872), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT98), .ZN(new_n878));
  INV_X1    g453(.A(new_n637), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n868), .A2(new_n872), .A3(new_n873), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G142), .ZN(new_n883));
  NOR2_X1   g458(.A1(G106), .A2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n486), .A2(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(G130), .B2(new_n495), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n627), .ZN(new_n888));
  INV_X1    g463(.A(G126), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n475), .B2(new_n476), .ZN(new_n890));
  INV_X1    g465(.A(new_n502), .ZN(new_n891));
  OAI21_X1  g466(.A(G2105), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(KEYINPUT4), .A2(G138), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n475), .B2(new_n476), .ZN(new_n894));
  INV_X1    g469(.A(new_n498), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n462), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n504), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n739), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(G164), .B1(new_n734), .B2(new_n738), .ZN(new_n900));
  INV_X1    g475(.A(new_n756), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n888), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n756), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n907));
  INV_X1    g482(.A(new_n627), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n887), .B(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n704), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n831), .B(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n904), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n904), .B2(new_n910), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n882), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n912), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n902), .A2(new_n888), .A3(new_n903), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n909), .B1(new_n906), .B2(new_n907), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n876), .A2(new_n881), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n904), .A2(new_n910), .A3(new_n912), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n915), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT99), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n915), .A2(new_n922), .A3(new_n926), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  XNOR2_X1  g505(.A(G305), .B(G290), .ZN(new_n931));
  XNOR2_X1  g506(.A(G303), .B(G288), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT42), .ZN(new_n934));
  XNOR2_X1  g509(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n616), .B2(new_n608), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n604), .A2(KEYINPUT100), .A3(G299), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT100), .B1(new_n604), .B2(G299), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n616), .A2(new_n608), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n604), .A2(G299), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT41), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n858), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n617), .B2(new_n619), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n617), .A3(new_n619), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n941), .B1(new_n938), .B2(new_n939), .ZN(new_n951));
  INV_X1    g526(.A(new_n949), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n947), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT102), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n953), .A3(KEYINPUT102), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n934), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n931), .A2(new_n932), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n931), .A2(new_n932), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT42), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(new_n954), .ZN(new_n962));
  OAI21_X1  g537(.A(G868), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n855), .A2(new_n621), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n930), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n950), .A2(new_n953), .A3(KEYINPUT102), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n961), .B1(new_n966), .B2(new_n954), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n955), .A2(new_n934), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n621), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n964), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n969), .A2(KEYINPUT103), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n965), .A2(new_n971), .ZN(G295));
  NAND2_X1  g547(.A1(new_n963), .A2(new_n964), .ZN(G331));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g549(.A1(G168), .A2(G171), .ZN(new_n975));
  NAND2_X1  g550(.A1(G286), .A2(G301), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n856), .A2(new_n975), .A3(new_n857), .A4(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n551), .A2(new_n855), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n551), .A2(new_n855), .ZN(new_n979));
  AND2_X1   g554(.A1(G286), .A2(G301), .ZN(new_n980));
  NOR2_X1   g555(.A1(G286), .A2(G301), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n978), .A2(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT104), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n975), .A2(new_n976), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT104), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n858), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n951), .A2(new_n977), .A3(new_n983), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n977), .ZN(new_n988));
  INV_X1    g563(.A(new_n935), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n604), .B2(G299), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT100), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n616), .B2(new_n608), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n992), .B2(new_n937), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n988), .B1(new_n993), .B2(new_n943), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n923), .B1(new_n995), .B2(new_n960), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n987), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n933), .B1(new_n995), .B2(KEYINPUT105), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n974), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n941), .A2(new_n942), .A3(KEYINPUT41), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n604), .A2(G299), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n992), .B2(new_n937), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1005), .B2(new_n989), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n983), .A2(new_n977), .A3(new_n986), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n977), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n992), .A2(new_n937), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(new_n941), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n982), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n933), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n983), .A2(new_n986), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n945), .A2(new_n988), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(G37), .B1(new_n1016), .B2(new_n933), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1017), .A3(KEYINPUT107), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n996), .B2(new_n1013), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1020), .A3(KEYINPUT43), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1002), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1014), .A2(new_n1017), .A3(new_n1001), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1025), .B2(new_n974), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n983), .A2(new_n986), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1027), .A2(new_n1005), .A3(new_n1009), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n982), .A2(new_n977), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n940), .B2(new_n944), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT105), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(new_n960), .A3(new_n998), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1001), .B1(new_n1032), .B2(new_n1017), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n996), .A2(new_n1013), .A3(KEYINPUT43), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1023), .B(new_n974), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1022), .B1(new_n1026), .B2(new_n1036), .ZN(G397));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT45), .B1(new_n898), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G40), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n473), .A2(new_n1040), .A3(new_n480), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G290), .A2(G1986), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(KEYINPUT108), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G290), .A2(G1986), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1048));
  INV_X1    g623(.A(new_n833), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n831), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n739), .B(new_n741), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n704), .B(G1996), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n831), .A2(new_n1049), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1048), .B1(new_n1043), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n898), .A2(new_n1038), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT50), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT50), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n898), .A2(new_n1059), .A3(new_n1038), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1058), .A2(new_n1041), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n719), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT45), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n898), .A2(KEYINPUT45), .A3(new_n1038), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(new_n772), .A3(new_n1041), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1066), .A2(new_n1067), .A3(KEYINPUT53), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT53), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1062), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1066), .A2(new_n1067), .A3(KEYINPUT53), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1061), .A2(KEYINPUT124), .A3(new_n719), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT124), .B1(new_n1061), .B2(new_n719), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1079), .A3(G301), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1071), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n1082));
  INV_X1    g657(.A(G8), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1041), .A2(new_n1065), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n714), .B1(new_n1084), .B2(new_n1039), .ZN(new_n1085));
  INV_X1    g660(.A(G2084), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1058), .A2(new_n1086), .A3(new_n1041), .A4(new_n1060), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1083), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT110), .B(G8), .Z(new_n1089));
  NOR2_X1   g664(.A1(G168), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT51), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(KEYINPUT51), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1060), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1059), .B1(new_n898), .B2(new_n1038), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n478), .A2(new_n479), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n462), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n469), .A2(new_n472), .ZN(new_n1097));
  OAI211_X1 g672(.A(G40), .B(new_n1096), .C1(new_n1097), .C2(new_n462), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1093), .A2(new_n1094), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1064), .A2(new_n1041), .A3(new_n1065), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1099), .A2(new_n1086), .B1(new_n1100), .B2(new_n714), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1092), .B1(new_n1101), .B2(new_n1089), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1091), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(new_n1090), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1081), .A2(new_n1082), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1062), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1061), .A2(KEYINPUT124), .A3(new_n719), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(G171), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT125), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(G171), .C1(new_n1108), .C2(new_n1112), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1074), .A2(new_n1075), .B1(new_n719), .B2(new_n1061), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1082), .B1(new_n1117), .B2(G301), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT55), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(G303), .B2(G8), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1120), .B(G8), .C1(new_n514), .C2(new_n521), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n808), .B1(new_n1084), .B2(new_n1039), .ZN(new_n1125));
  INV_X1    g700(.A(G2090), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1058), .A2(new_n1126), .A3(new_n1041), .A4(new_n1060), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1089), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT109), .ZN(new_n1132));
  AND4_X1   g707(.A1(new_n1132), .A2(new_n1128), .A3(G8), .A4(new_n1124), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1083), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1134), .B2(new_n1124), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1131), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT112), .B(G1981), .Z(new_n1137));
  NAND3_X1  g712(.A1(new_n579), .A2(new_n583), .A3(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT113), .B(G86), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n517), .B(new_n1139), .C1(new_n528), .C2(new_n506), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1140), .A2(KEYINPUT114), .A3(new_n582), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT114), .B1(new_n1140), .B2(new_n582), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1141), .A2(new_n1142), .A3(new_n574), .ZN(new_n1143));
  INV_X1    g718(.A(G1981), .ZN(new_n1144));
  OAI211_X1 g719(.A(KEYINPUT49), .B(new_n1138), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT115), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1140), .A2(new_n582), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT114), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n574), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1140), .A2(KEYINPUT114), .A3(new_n582), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G1981), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1153), .A2(KEYINPUT115), .A3(KEYINPUT49), .A4(new_n1138), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT49), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1138), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1144), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n898), .A2(new_n1038), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1089), .B1(new_n1159), .B2(new_n1041), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1147), .A2(new_n1154), .A3(new_n1158), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT52), .ZN(new_n1162));
  INV_X1    g737(.A(G1976), .ZN(new_n1163));
  OR2_X1    g738(.A1(G288), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1162), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1166));
  XNOR2_X1  g741(.A(KEYINPUT111), .B(G1976), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT52), .B1(G288), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1165), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT117), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1161), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1161), .B2(new_n1169), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1136), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1107), .A2(new_n1119), .A3(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1099), .A2(G1956), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1084), .A2(new_n1039), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT56), .B(G2072), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(KEYINPUT119), .A3(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1064), .A2(new_n1177), .A3(new_n1041), .A4(new_n1065), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT119), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1175), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n563), .A2(KEYINPUT118), .A3(new_n565), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(G299), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1186), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1175), .A2(new_n1188), .A3(new_n1178), .A4(new_n1181), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n1191));
  OAI21_X1  g766(.A(KEYINPUT122), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT59), .ZN(new_n1193));
  INV_X1    g768(.A(G1996), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1176), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT120), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n1098), .B2(new_n1057), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1159), .A2(KEYINPUT120), .A3(new_n1041), .ZN(new_n1198));
  XNOR2_X1  g773(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(G1341), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1195), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1193), .B1(new_n1202), .B2(new_n552), .ZN(new_n1203));
  AOI211_X1 g778(.A(KEYINPUT59), .B(new_n551), .C1(new_n1195), .C2(new_n1201), .ZN(new_n1204));
  AOI21_X1  g779(.A(G2067), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1061), .A2(new_n788), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT60), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n604), .A2(new_n1209), .ZN(new_n1210));
  OAI22_X1  g785(.A1(new_n1203), .A2(new_n1204), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1208), .A2(new_n604), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1206), .A2(new_n616), .A3(new_n1207), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1209), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT122), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1187), .A2(new_n1189), .A3(new_n1216), .A4(KEYINPUT61), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1192), .A2(new_n1215), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1189), .A2(new_n604), .A3(new_n1208), .ZN(new_n1220));
  AND2_X1   g795(.A1(new_n1220), .A2(new_n1187), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1174), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1128), .A2(G8), .A3(new_n1124), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1223), .A2(KEYINPUT109), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1134), .A2(new_n1132), .A3(new_n1124), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1161), .A2(new_n1169), .ZN(new_n1227));
  XOR2_X1   g802(.A(new_n1138), .B(KEYINPUT116), .Z(new_n1228));
  NOR2_X1   g803(.A1(G288), .A2(G1976), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1228), .B1(new_n1161), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(new_n1160), .ZN(new_n1231));
  OAI22_X1  g806(.A1(new_n1226), .A2(new_n1227), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1233), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1234));
  AOI211_X1 g809(.A(KEYINPUT62), .B(new_n1105), .C1(new_n1091), .C2(new_n1102), .ZN(new_n1235));
  NOR2_X1   g810(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1130), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1227), .A2(KEYINPUT117), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1161), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1239));
  AOI21_X1  g814(.A(G301), .B1(new_n1076), .B2(new_n1062), .ZN(new_n1240));
  AND4_X1   g815(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1232), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  NOR3_X1   g817(.A1(new_n1101), .A2(G286), .A3(new_n1089), .ZN(new_n1243));
  NAND4_X1  g818(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1243), .ZN(new_n1244));
  INV_X1    g819(.A(KEYINPUT63), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1243), .A2(KEYINPUT63), .ZN(new_n1247));
  NOR2_X1   g822(.A1(new_n1134), .A2(new_n1124), .ZN(new_n1248));
  NOR3_X1   g823(.A1(new_n1247), .A2(new_n1227), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1249), .A2(new_n1226), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1242), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g827(.A(new_n1056), .B1(new_n1222), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g828(.A(new_n1043), .B1(new_n1051), .B2(new_n911), .ZN(new_n1254));
  NAND3_X1  g829(.A1(new_n1043), .A2(KEYINPUT46), .A3(new_n1194), .ZN(new_n1255));
  INV_X1    g830(.A(KEYINPUT46), .ZN(new_n1256));
  OAI21_X1  g831(.A(new_n1256), .B1(new_n1042), .B2(G1996), .ZN(new_n1257));
  NAND3_X1  g832(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  XOR2_X1   g833(.A(new_n1258), .B(KEYINPUT47), .Z(new_n1259));
  NAND2_X1  g834(.A1(new_n1055), .A2(new_n1043), .ZN(new_n1260));
  NAND2_X1  g835(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1261));
  XNOR2_X1  g836(.A(new_n1261), .B(KEYINPUT48), .ZN(new_n1262));
  AOI21_X1  g837(.A(new_n1259), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g838(.A1(new_n739), .A2(new_n741), .ZN(new_n1264));
  AOI21_X1  g839(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1265));
  OAI21_X1  g840(.A(new_n1264), .B1(new_n1265), .B2(new_n1050), .ZN(new_n1266));
  INV_X1    g841(.A(KEYINPUT126), .ZN(new_n1267));
  AOI21_X1  g842(.A(new_n1042), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g843(.A(new_n1268), .B1(new_n1267), .B2(new_n1266), .ZN(new_n1269));
  AND2_X1   g844(.A1(new_n1263), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g845(.A1(new_n1253), .A2(new_n1270), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g846(.A1(G227), .A2(new_n460), .ZN(new_n1273));
  NAND3_X1  g847(.A1(new_n694), .A2(new_n656), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g848(.A(new_n1274), .B1(new_n925), .B2(new_n927), .ZN(new_n1275));
  INV_X1    g849(.A(KEYINPUT127), .ZN(new_n1276));
  OAI211_X1 g850(.A(new_n1275), .B(new_n1276), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1277));
  INV_X1    g851(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g852(.A(new_n1276), .B1(new_n1025), .B2(new_n1275), .ZN(new_n1279));
  NOR2_X1   g853(.A1(new_n1278), .A2(new_n1279), .ZN(G308));
  NAND2_X1  g854(.A1(new_n1025), .A2(new_n1275), .ZN(new_n1281));
  NAND2_X1  g855(.A1(new_n1281), .A2(KEYINPUT127), .ZN(new_n1282));
  NAND2_X1  g856(.A1(new_n1282), .A2(new_n1277), .ZN(G225));
endmodule


