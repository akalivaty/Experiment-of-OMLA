//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n211), .B(new_n213), .C1(G50), .C2(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G116), .ZN(new_n217));
  INV_X1    g0017(.A(G270), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n206), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(G1), .ZN(new_n230));
  INV_X1    g0030(.A(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n229), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n224), .A2(new_n227), .A3(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT66), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n232), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n254), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G223), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G1698), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G222), .B2(G1698), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n256), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G77), .B2(new_n260), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n230), .B1(G41), .B2(G45), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n256), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G226), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n265), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G190), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G200), .ZN(new_n276));
  INV_X1    g0076(.A(new_n272), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n203), .A2(G20), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT8), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G58), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT67), .B(G58), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n254), .A2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n278), .B1(new_n279), .B2(new_n281), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n206), .A2(new_n254), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(new_n232), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n230), .A2(G13), .A3(G20), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n291), .A2(new_n294), .B1(new_n202), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n293), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n230), .A2(G20), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT70), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(G50), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n307), .A2(KEYINPUT9), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(KEYINPUT9), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n275), .B1(new_n276), .B2(new_n277), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(KEYINPUT72), .A3(KEYINPUT10), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n307), .B1(G169), .B2(new_n277), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT71), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n317), .C1(G179), .C2(new_n272), .ZN(new_n318));
  NAND2_X1  g0118(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n310), .A2(new_n319), .A3(new_n311), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n302), .A2(G77), .A3(new_n305), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G20), .A2(G77), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n322), .B1(new_n323), .B2(new_n281), .C1(new_n324), .C2(new_n290), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(new_n294), .B1(new_n299), .B2(new_n207), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n256), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G232), .A2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G238), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n260), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n328), .B(new_n332), .C1(G107), .C2(new_n260), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n256), .A2(new_n266), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n271), .C1(new_n208), .C2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n327), .B1(G200), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n273), .B2(new_n335), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n313), .A2(new_n318), .A3(new_n320), .A4(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT78), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(KEYINPUT3), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n257), .A2(KEYINPUT78), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n254), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n343), .A2(KEYINPUT7), .A3(new_n234), .A4(new_n259), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n260), .B2(G20), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n220), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n280), .A2(G159), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n201), .B1(new_n286), .B2(G68), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n234), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n339), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n257), .A2(KEYINPUT78), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n340), .A2(KEYINPUT3), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(G33), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(new_n234), .A3(new_n258), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT7), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n354), .A2(new_n345), .A3(new_n234), .A4(new_n258), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(G68), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n286), .A2(G68), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n228), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n351), .A2(new_n294), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n270), .B1(new_n267), .B2(G232), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n354), .A2(new_n258), .B1(new_n261), .B2(new_n330), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n330), .A2(G226), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n365), .A2(new_n366), .B1(G33), .B2(G87), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n364), .B(G190), .C1(new_n367), .C2(new_n256), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n288), .A2(new_n304), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n302), .B1(new_n299), .B2(new_n288), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n354), .A2(new_n258), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n261), .A2(new_n330), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n372), .A3(new_n366), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G87), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n256), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n271), .B1(new_n334), .B2(new_n216), .ZN(new_n376));
  OAI21_X1  g0176(.A(G200), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n363), .A2(new_n368), .A3(new_n370), .A4(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT17), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n285), .A2(new_n287), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n305), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n382), .A2(new_n301), .B1(new_n298), .B2(new_n381), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n220), .B1(new_n355), .B2(KEYINPUT7), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n350), .B1(new_n384), .B2(new_n357), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n293), .B1(new_n385), .B2(KEYINPUT16), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n351), .ZN(new_n387));
  OAI21_X1  g0187(.A(G169), .B1(new_n375), .B2(new_n376), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n364), .B(G179), .C1(new_n367), .C2(new_n256), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n380), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n362), .A2(new_n294), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n344), .A2(new_n346), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G68), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT16), .B1(new_n395), .B2(new_n361), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n370), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(KEYINPUT18), .A3(new_n390), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n379), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT79), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n335), .A2(G179), .ZN(new_n402));
  INV_X1    g0202(.A(G169), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n335), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n327), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n260), .B1(G232), .B2(new_n330), .ZN(new_n407));
  NOR2_X1   g0207(.A1(G226), .A2(G1698), .ZN(new_n408));
  INV_X1    g0208(.A(G97), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n407), .A2(new_n408), .B1(new_n254), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n270), .B1(new_n410), .B2(new_n328), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n221), .B2(new_n334), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n412), .A2(KEYINPUT13), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(KEYINPUT13), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OR3_X1    g0215(.A1(new_n415), .A2(KEYINPUT14), .A3(new_n403), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(G179), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT14), .B1(new_n415), .B2(new_n403), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n298), .B2(G68), .ZN(new_n421));
  XOR2_X1   g0221(.A(new_n421), .B(KEYINPUT76), .Z(new_n422));
  NAND2_X1  g0222(.A1(new_n299), .A2(new_n220), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(KEYINPUT12), .B2(new_n423), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n290), .A2(new_n207), .B1(new_n234), .B2(G68), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n281), .A2(new_n202), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n294), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT11), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n301), .A2(new_n220), .A3(new_n304), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT74), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT77), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n419), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT73), .B1(new_n415), .B2(new_n276), .ZN(new_n435));
  INV_X1    g0235(.A(new_n431), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n415), .A2(G190), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT73), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(G200), .C1(new_n413), .C2(new_n414), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n338), .A2(new_n406), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G87), .ZN(new_n443));
  AOI211_X1 g0243(.A(G20), .B(new_n443), .C1(new_n354), .C2(new_n258), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT22), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT86), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n443), .A2(KEYINPUT22), .A3(G20), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n260), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT87), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n371), .A2(new_n234), .A3(G87), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT86), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT22), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n446), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT23), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n234), .B2(G107), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n209), .A2(KEYINPUT23), .A3(G20), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n455), .A2(new_n456), .B1(new_n289), .B2(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT88), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT88), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n453), .A2(new_n460), .A3(new_n457), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(KEYINPUT24), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(KEYINPUT88), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n294), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n298), .A2(G107), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n230), .A2(G33), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n302), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n468), .A2(new_n469), .B1(new_n472), .B2(G107), .ZN(new_n473));
  OR2_X1    g0273(.A1(G250), .A2(G1698), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n330), .A2(G257), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n371), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G294), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n254), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT90), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n371), .A2(new_n474), .A3(new_n475), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT90), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n481), .C1(new_n254), .C2(new_n477), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n328), .A3(new_n482), .ZN(new_n483));
  XOR2_X1   g0283(.A(KEYINPUT5), .B(G41), .Z(new_n484));
  NAND3_X1  g0284(.A1(new_n230), .A2(G45), .A3(G274), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XOR2_X1   g0286(.A(new_n486), .B(KEYINPUT82), .Z(new_n487));
  NAND2_X1  g0287(.A1(new_n230), .A2(G45), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n256), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G264), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n483), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n276), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(G190), .B2(new_n492), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n465), .A2(new_n473), .A3(new_n494), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n486), .B(KEYINPUT82), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(G257), .B2(new_n490), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT80), .ZN(new_n500));
  XNOR2_X1  g0300(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n371), .A2(new_n503), .A3(G244), .A4(new_n330), .ZN(new_n504));
  AOI21_X1  g0304(.A(G1698), .B1(new_n258), .B2(new_n259), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G244), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n502), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT81), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n508), .A2(new_n509), .A3(new_n256), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n498), .A2(new_n501), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n503), .A2(G244), .ZN(new_n512));
  AOI211_X1 g0312(.A(G1698), .B(new_n512), .C1(new_n354), .C2(new_n258), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n503), .B1(new_n505), .B2(G244), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT81), .B1(new_n515), .B2(new_n328), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n497), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT83), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n497), .B(KEYINPUT83), .C1(new_n510), .C2(new_n516), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(G200), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n298), .A2(G97), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n471), .A2(new_n409), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n394), .A2(G107), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT6), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n409), .A2(new_n209), .ZN(new_n526));
  NOR2_X1   g0326(.A1(G97), .A2(G107), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI221_X1 g0330(.A(new_n524), .B1(new_n234), .B2(new_n530), .C1(new_n207), .C2(new_n281), .ZN(new_n531));
  AOI211_X1 g0331(.A(new_n522), .B(new_n523), .C1(new_n531), .C2(new_n294), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n515), .A2(new_n328), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n497), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G190), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n521), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n489), .A2(new_n218), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n210), .A2(G1698), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n371), .B(new_n540), .C1(G257), .C2(G1698), .ZN(new_n541));
  INV_X1    g0341(.A(new_n260), .ZN(new_n542));
  XOR2_X1   g0342(.A(KEYINPUT85), .B(G303), .Z(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n487), .B(new_n539), .C1(new_n545), .C2(new_n256), .ZN(new_n546));
  INV_X1    g0346(.A(G179), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n298), .A2(new_n293), .A3(G116), .A4(new_n470), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n299), .A2(new_n217), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n234), .A2(G116), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n293), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(G20), .B1(new_n254), .B2(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n501), .A2(new_n553), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n552), .A2(new_n554), .A3(KEYINPUT20), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT20), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n549), .B(new_n550), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n256), .B1(new_n541), .B2(new_n544), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(new_n496), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(G190), .A3(new_n539), .ZN(new_n561));
  INV_X1    g0361(.A(new_n557), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n559), .A2(new_n496), .A3(new_n538), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n562), .C1(new_n276), .C2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n546), .A2(KEYINPUT21), .A3(G169), .A4(new_n557), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n557), .A2(G169), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n563), .ZN(new_n568));
  AND4_X1   g0368(.A1(new_n558), .A2(new_n564), .A3(new_n565), .A4(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n522), .B1(new_n531), .B2(new_n294), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n409), .B2(new_n471), .ZN(new_n571));
  INV_X1    g0371(.A(new_n517), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n547), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n534), .A2(new_n403), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n495), .A2(new_n537), .A3(new_n569), .A4(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n492), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(G169), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n492), .A2(G179), .ZN(new_n579));
  AOI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n465), .C2(new_n473), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT84), .ZN(new_n581));
  INV_X1    g0381(.A(new_n258), .ZN(new_n582));
  XNOR2_X1  g0382(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(G33), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n208), .A2(new_n330), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n581), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G116), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n371), .A2(G238), .A3(new_n330), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n371), .A2(KEYINPUT84), .A3(new_n585), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n328), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n256), .A2(G250), .A3(new_n488), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n485), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n299), .A2(new_n324), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n371), .A2(new_n234), .A3(G68), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT19), .B1(new_n289), .B2(G97), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n527), .A2(new_n443), .ZN(new_n599));
  NAND3_X1  g0399(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n234), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n293), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  AOI211_X1 g0403(.A(new_n596), .B(new_n603), .C1(new_n472), .C2(G87), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n595), .B(new_n604), .C1(new_n273), .C2(new_n594), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n594), .A2(new_n403), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n596), .A2(new_n603), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n324), .B2(new_n471), .ZN(new_n608));
  INV_X1    g0408(.A(new_n485), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n591), .B2(new_n328), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n547), .A3(new_n593), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n576), .A2(new_n580), .A3(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n442), .A2(new_n614), .ZN(G372));
  INV_X1    g0415(.A(KEYINPUT92), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT91), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n606), .B2(new_n611), .ZN(new_n618));
  AOI21_X1  g0418(.A(G169), .B1(new_n610), .B2(new_n593), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(KEYINPUT91), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n616), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n610), .A2(new_n547), .A3(new_n593), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT91), .B1(new_n622), .B2(new_n619), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n606), .A2(new_n617), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(KEYINPUT92), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n621), .A2(new_n625), .A3(new_n608), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n495), .A2(new_n537), .A3(new_n605), .A4(new_n575), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n465), .A2(new_n473), .ZN(new_n630));
  INV_X1    g0430(.A(new_n578), .ZN(new_n631));
  INV_X1    g0431(.A(new_n579), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n568), .A2(new_n565), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n558), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n627), .B1(new_n629), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  INV_X1    g0439(.A(new_n575), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n626), .A2(new_n639), .A3(new_n605), .A4(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT26), .B1(new_n575), .B2(new_n613), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n442), .A2(new_n643), .ZN(new_n644));
  AOI221_X4 g0444(.A(new_n380), .B1(new_n388), .B2(new_n389), .C1(new_n363), .C2(new_n370), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT18), .B1(new_n397), .B2(new_n390), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n440), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n434), .B1(new_n648), .B2(new_n405), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n649), .B2(new_n379), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n313), .A2(new_n320), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n318), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n644), .A2(new_n652), .ZN(G369));
  AND2_X1   g0453(.A1(new_n633), .A2(new_n495), .ZN(new_n654));
  XOR2_X1   g0454(.A(KEYINPUT93), .B(KEYINPUT27), .Z(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n231), .A2(G20), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(G1), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n655), .A2(new_n230), .A3(new_n657), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n630), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n663), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n633), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n557), .A2(new_n663), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n569), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n636), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n580), .A2(new_n666), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n636), .A2(new_n663), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n654), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n225), .ZN(new_n678));
  OR3_X1    g0478(.A1(new_n678), .A2(KEYINPUT94), .A3(G41), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT94), .B1(new_n678), .B2(G41), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n527), .A2(new_n443), .A3(new_n217), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n682), .A2(new_n230), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n229), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT28), .Z(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  INV_X1    g0488(.A(new_n594), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n483), .A2(new_n491), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n535), .A2(new_n548), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT30), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n572), .A2(new_n689), .A3(new_n563), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n547), .A3(new_n492), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n666), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n495), .A2(new_n575), .A3(new_n537), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n578), .B1(new_n465), .B2(new_n473), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n613), .B1(new_n697), .B2(new_n632), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n696), .A2(new_n698), .A3(new_n569), .A4(new_n666), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n695), .B1(new_n699), .B2(KEYINPUT31), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n695), .A2(KEYINPUT95), .A3(KEYINPUT31), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n695), .A2(KEYINPUT31), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT95), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n688), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n643), .A2(new_n708), .A3(new_n666), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n575), .A2(new_n613), .A3(KEYINPUT26), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n626), .A2(new_n605), .A3(new_n640), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(KEYINPUT26), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n663), .B1(new_n638), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n709), .B1(new_n708), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n707), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n687), .B1(new_n715), .B2(G1), .ZN(G364));
  AOI21_X1  g0516(.A(new_n230), .B1(new_n657), .B2(G45), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n682), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n672), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G330), .B2(new_n670), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n371), .A2(new_n678), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n248), .B2(G45), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(G45), .B2(new_n229), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n260), .A2(G355), .A3(new_n225), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n725), .B(new_n726), .C1(G116), .C2(new_n225), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n233), .B1(G20), .B2(new_n403), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n234), .A2(new_n273), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G179), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n276), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n234), .A2(G190), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(G179), .A3(new_n276), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n736), .A2(G326), .B1(new_n739), .B2(G311), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G179), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G329), .ZN(new_n744));
  INV_X1    g0544(.A(G303), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n276), .A2(G179), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n734), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n740), .B(new_n744), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n737), .A2(G179), .A3(G200), .ZN(new_n749));
  OR2_X1    g0549(.A1(KEYINPUT33), .A2(G317), .ZN(new_n750));
  NAND2_X1  g0550(.A1(KEYINPUT33), .A2(G317), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n737), .A2(new_n746), .ZN(new_n753));
  INV_X1    g0553(.A(G283), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n748), .A2(new_n260), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n735), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G322), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n234), .B1(new_n741), .B2(G190), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n756), .B(new_n758), .C1(new_n477), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT97), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n749), .A2(new_n220), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n753), .A2(new_n209), .ZN(new_n763));
  INV_X1    g0563(.A(new_n736), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n743), .A2(G159), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n202), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n763), .B(new_n767), .C1(new_n765), .C2(new_n766), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n542), .B1(new_n739), .B2(G77), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n759), .A2(new_n409), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n747), .A2(new_n443), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n770), .B(new_n771), .C1(new_n286), .C2(new_n757), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n768), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n761), .B1(new_n762), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n733), .B1(new_n774), .B2(new_n728), .ZN(new_n775));
  INV_X1    g0575(.A(new_n731), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n775), .B(new_n719), .C1(new_n670), .C2(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n721), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  NOR2_X1   g0579(.A1(new_n405), .A2(new_n663), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n327), .A2(new_n663), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n337), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(new_n782), .B2(new_n405), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT98), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n729), .ZN(new_n786));
  INV_X1    g0586(.A(new_n749), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n757), .A2(G143), .B1(new_n787), .B2(G150), .ZN(new_n788));
  INV_X1    g0588(.A(G137), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n788), .B1(new_n789), .B2(new_n764), .C1(new_n790), .C2(new_n738), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT34), .ZN(new_n792));
  INV_X1    g0592(.A(new_n759), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n286), .ZN(new_n794));
  INV_X1    g0594(.A(new_n747), .ZN(new_n795));
  INV_X1    g0595(.A(new_n753), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G50), .A2(new_n795), .B1(new_n796), .B2(G68), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n584), .B1(G132), .B2(new_n743), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n792), .A2(new_n794), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n749), .A2(new_n754), .ZN(new_n800));
  INV_X1    g0600(.A(new_n757), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n477), .B1(new_n742), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G303), .B2(new_n736), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n260), .B1(new_n796), .B2(G87), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n739), .A2(G116), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n770), .B1(G107), .B2(new_n795), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n799), .B1(new_n800), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n728), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n728), .A2(new_n729), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n207), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n786), .A2(new_n719), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n785), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n643), .B2(new_n666), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n641), .A2(new_n642), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n635), .B1(new_n697), .B2(new_n632), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n626), .B1(new_n817), .B2(new_n628), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n814), .B(new_n666), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(new_n707), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n813), .B1(new_n822), .B2(new_n719), .ZN(G384));
  INV_X1    g0623(.A(new_n695), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n576), .A2(new_n580), .A3(new_n613), .A4(new_n663), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT31), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n704), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n442), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT102), .ZN(new_n830));
  INV_X1    g0630(.A(new_n661), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n358), .A2(new_n361), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n339), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n383), .B1(new_n386), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n387), .A2(KEYINPUT17), .A3(new_n368), .A4(new_n377), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT17), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n378), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n831), .B(new_n835), .C1(new_n647), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n390), .A2(new_n831), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n378), .B1(new_n841), .B2(new_n834), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT37), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n351), .A2(new_n294), .A3(new_n362), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n844), .A2(new_n383), .B1(new_n390), .B2(new_n831), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(new_n846), .A3(new_n378), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n840), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n433), .A2(new_n663), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n434), .A2(new_n440), .A3(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n433), .B(new_n663), .C1(new_n648), .C2(new_n419), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n785), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n704), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n853), .B(new_n857), .C1(new_n700), .C2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT40), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n397), .A2(new_n831), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n379), .B2(new_n399), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n845), .A2(new_n846), .A3(new_n378), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n846), .B1(new_n845), .B2(new_n378), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n850), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n867), .A2(new_n852), .A3(KEYINPUT101), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT101), .B1(new_n867), .B2(new_n852), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n868), .A2(new_n869), .A3(new_n860), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n828), .A2(new_n870), .A3(new_n857), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n861), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n830), .B(new_n872), .Z(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(G330), .ZN(new_n874));
  INV_X1    g0674(.A(new_n853), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n855), .A2(new_n856), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n780), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n875), .B(new_n877), .C1(new_n819), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n434), .A2(new_n663), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT99), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n867), .A2(new_n852), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT100), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n875), .B2(new_n882), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n840), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n840), .B2(new_n848), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT100), .B(KEYINPUT39), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n881), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n399), .A2(new_n831), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n879), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n652), .B1(new_n714), .B2(new_n442), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n891), .B(new_n892), .Z(new_n893));
  XNOR2_X1  g0693(.A(new_n874), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n230), .B2(new_n657), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT35), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n234), .B(new_n233), .C1(new_n530), .C2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(G116), .C1(new_n896), .C2(new_n530), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n685), .A2(new_n359), .A3(G77), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(G50), .B2(new_n220), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(G1), .A3(new_n231), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n895), .A2(new_n899), .A3(new_n902), .ZN(G367));
  OAI221_X1 g0703(.A(new_n732), .B1(new_n225), .B2(new_n324), .C1(new_n723), .C2(new_n244), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT105), .ZN(new_n905));
  INV_X1    g0705(.A(G317), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n738), .A2(new_n754), .B1(new_n742), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n757), .A2(new_n543), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n747), .A2(new_n217), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n908), .B1(KEYINPUT46), .B2(new_n909), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n907), .B(new_n910), .C1(KEYINPUT46), .C2(new_n909), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n753), .A2(new_n409), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n749), .A2(new_n477), .B1(new_n759), .B2(new_n209), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(G311), .B2(new_n736), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n911), .A2(new_n584), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n757), .A2(G150), .B1(new_n787), .B2(G159), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n207), .B2(new_n753), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n542), .B(new_n918), .C1(G137), .C2(new_n743), .ZN(new_n919));
  AOI22_X1  g0719(.A1(G50), .A2(new_n739), .B1(new_n795), .B2(new_n286), .ZN(new_n920));
  INV_X1    g0720(.A(G143), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n919), .B(new_n920), .C1(new_n921), .C2(new_n764), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n759), .A2(new_n220), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT47), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n905), .B1(new_n925), .B2(new_n728), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n604), .A2(new_n666), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n626), .A2(new_n605), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n626), .B2(new_n927), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n926), .B(new_n719), .C1(new_n929), .C2(new_n776), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n676), .A2(new_n674), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n537), .A2(new_n575), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n571), .B2(new_n663), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n640), .B2(new_n663), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT44), .Z(new_n936));
  NOR2_X1   g0736(.A1(new_n931), .A2(new_n934), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n673), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(KEYINPUT104), .B(new_n676), .C1(new_n667), .C2(new_n675), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(KEYINPUT104), .B2(new_n676), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(new_n671), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n715), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n715), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n681), .B(KEYINPUT41), .Z(new_n948));
  AOI21_X1  g0748(.A(new_n718), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n934), .A2(new_n676), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT42), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n580), .A2(new_n537), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n663), .B1(new_n953), .B2(new_n575), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n950), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT103), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n673), .A2(new_n934), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n955), .B(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n930), .B1(new_n949), .B2(new_n960), .ZN(G387));
  OR2_X1    g0761(.A1(new_n944), .A2(new_n715), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(new_n682), .A3(new_n945), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n944), .A2(new_n718), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n667), .A2(new_n776), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n801), .A2(new_n202), .B1(new_n742), .B2(new_n279), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n912), .B(new_n966), .C1(G68), .C2(new_n739), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n759), .A2(new_n324), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n747), .A2(new_n207), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(G159), .C2(new_n736), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n381), .A2(new_n787), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n967), .A2(new_n371), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n736), .A2(G322), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n802), .B2(new_n749), .C1(new_n801), .C2(new_n906), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n543), .B2(new_n739), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT48), .Z(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n754), .B2(new_n759), .C1(new_n477), .C2(new_n747), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT49), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n743), .A2(G326), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n979), .B(new_n584), .C1(new_n217), .C2(new_n753), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n972), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n728), .ZN(new_n982));
  INV_X1    g0782(.A(G45), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n722), .B1(new_n241), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n260), .A2(new_n683), .A3(new_n225), .ZN(new_n985));
  AOI211_X1 g0785(.A(G45), .B(new_n683), .C1(G68), .C2(G77), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n323), .A2(G50), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT50), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n225), .A2(G107), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n732), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n965), .A2(new_n719), .A3(new_n982), .A4(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n963), .A2(new_n964), .A3(new_n992), .ZN(G393));
  NAND2_X1  g0793(.A1(new_n934), .A2(new_n731), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT106), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n260), .B(new_n763), .C1(G322), .C2(new_n743), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n754), .B2(new_n747), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT107), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n787), .A2(new_n543), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n739), .A2(G294), .B1(new_n793), .B2(G116), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n757), .A2(G311), .B1(new_n736), .B2(G317), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT52), .Z(new_n1002));
  NAND4_X1  g0802(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n749), .A2(new_n202), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n757), .A2(G159), .B1(new_n736), .B2(G150), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT51), .Z(new_n1006));
  OAI22_X1  g0806(.A1(new_n747), .A2(new_n220), .B1(new_n753), .B2(new_n443), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n921), .A2(new_n742), .B1(new_n759), .B2(new_n207), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n738), .A2(new_n323), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n371), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1003), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n728), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n252), .A2(new_n722), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n732), .C1(new_n409), .C2(new_n225), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n995), .A2(new_n719), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n941), .A2(new_n945), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT108), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n946), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n682), .B1(new_n1017), .B2(KEYINPUT108), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1016), .B1(new_n717), .B2(new_n941), .C1(new_n1019), .C2(new_n1020), .ZN(G390));
  NOR2_X1   g0821(.A1(new_n868), .A2(new_n869), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n780), .B1(new_n713), .B2(new_n814), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1022), .B(new_n881), .C1(new_n1023), .C2(new_n877), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n853), .A2(KEYINPUT39), .B1(new_n883), .B2(KEYINPUT100), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n888), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n877), .B1(new_n819), .B2(new_n878), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n881), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n826), .B1(new_n614), .B2(new_n666), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n706), .B(new_n701), .C1(new_n1031), .C2(new_n695), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1032), .A2(G330), .A3(new_n814), .A4(new_n876), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1024), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT109), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1024), .A2(new_n1030), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n876), .A2(new_n814), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n827), .B2(new_n704), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(G330), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT109), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1024), .A2(new_n1030), .A3(new_n1042), .A4(new_n1033), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1035), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n828), .A2(new_n442), .A3(G330), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT110), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n892), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(G330), .B1(new_n700), .B2(new_n858), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT111), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g0852(.A(KEYINPUT111), .B(G330), .C1(new_n700), .C2(new_n858), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n814), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n877), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n1023), .A3(new_n1033), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n876), .B1(new_n707), .B2(new_n814), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1057), .A2(new_n1040), .B1(new_n780), .B2(new_n820), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1049), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT112), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1044), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1035), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n820), .A2(new_n780), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1032), .A2(G330), .A3(new_n814), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n877), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1063), .B1(new_n1065), .B2(new_n1039), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1033), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n877), .B2(new_n1054), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1066), .B1(new_n1068), .B2(new_n1023), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1062), .B(KEYINPUT112), .C1(new_n1069), .C2(new_n1049), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1061), .A2(new_n682), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n743), .A2(G125), .ZN(new_n1072));
  INV_X1    g0872(.A(G132), .ZN(new_n1073));
  INV_X1    g0873(.A(G128), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1072), .B1(new_n801), .B2(new_n1073), .C1(new_n1074), .C2(new_n764), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT54), .B(G143), .Z(new_n1076));
  AOI21_X1  g0876(.A(new_n1075), .B1(new_n739), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n787), .A2(G137), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n795), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n747), .B2(new_n279), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1079), .A2(new_n1081), .B1(G159), .B2(new_n793), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n260), .B1(new_n753), .B2(new_n202), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT113), .Z(new_n1084));
  NAND4_X1  g0884(.A1(new_n1077), .A2(new_n1078), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n542), .B1(new_n477), .B2(new_n742), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n801), .A2(new_n217), .B1(new_n764), .B2(new_n754), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n409), .A2(new_n738), .B1(new_n749), .B2(new_n209), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(KEYINPUT114), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n771), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G68), .A2(new_n796), .B1(new_n793), .B2(G77), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1085), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1094), .A2(new_n728), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n811), .A2(new_n288), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n1027), .C2(new_n729), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1044), .A2(new_n718), .B1(new_n719), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1071), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT115), .ZN(G378));
  INV_X1    g0900(.A(new_n307), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(new_n661), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n318), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1102), .B1(new_n651), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1102), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n313), .A2(new_n318), .A3(new_n320), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1104), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n729), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1073), .A2(new_n749), .B1(new_n738), .B2(new_n789), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G125), .B2(new_n736), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n757), .A2(G128), .B1(G150), .B2(new_n793), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1076), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1115), .B(new_n1116), .C1(new_n747), .C2(new_n1117), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT59), .Z(new_n1119));
  OAI21_X1  g0919(.A(new_n254), .B1(new_n753), .B2(new_n790), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G124), .B2(new_n743), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n255), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n354), .A2(new_n255), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(G50), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n324), .B2(new_n738), .ZN(new_n1126));
  NOR4_X1   g0926(.A1(new_n1126), .A2(new_n582), .A3(new_n923), .A4(new_n969), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n796), .A2(new_n286), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n757), .A2(G107), .B1(new_n787), .B2(G97), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n736), .A2(G116), .B1(G283), .B2(new_n743), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT58), .Z(new_n1132));
  OAI21_X1  g0932(.A(new_n728), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n811), .A2(new_n202), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1113), .A2(new_n719), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT116), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n861), .A2(new_n871), .A3(G330), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1112), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1139), .A2(new_n861), .A3(G330), .A4(new_n871), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1138), .A2(new_n891), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n891), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1136), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n891), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT116), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1135), .B1(new_n1148), .B2(new_n717), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT117), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1049), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1138), .A2(new_n891), .A3(new_n1140), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1146), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1150), .B1(new_n1156), .B2(new_n682), .ZN(new_n1157));
  AOI211_X1 g0957(.A(KEYINPUT117), .B(new_n681), .C1(new_n1152), .C2(new_n1155), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1049), .B1(new_n1044), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1153), .B1(new_n1148), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1149), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(G375));
  NAND2_X1  g0964(.A1(new_n877), .A2(new_n729), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n542), .B1(new_n764), .B2(new_n477), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n747), .A2(new_n409), .B1(new_n742), .B2(new_n745), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n787), .A2(G116), .B1(new_n739), .B2(G107), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n968), .B(new_n1167), .C1(new_n1168), .C2(KEYINPUT118), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(KEYINPUT118), .B2(new_n1168), .C1(new_n754), .C2(new_n801), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1166), .B(new_n1170), .C1(G77), .C2(new_n796), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n757), .A2(G137), .B1(new_n739), .B2(G150), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1172), .B(new_n1128), .C1(new_n1074), .C2(new_n742), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n759), .A2(new_n202), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n764), .A2(new_n1073), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n371), .B1(new_n790), .B2(new_n747), .C1(new_n1117), .C2(new_n749), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n728), .B1(new_n1171), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n811), .A2(new_n220), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1165), .A2(new_n719), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n1069), .B2(new_n717), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT119), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1069), .A2(new_n1049), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1059), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n1185), .A3(new_n948), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(G381));
  INV_X1    g0988(.A(KEYINPUT121), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1071), .A2(new_n1189), .A3(new_n1098), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1189), .B1(new_n1071), .B2(new_n1098), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(G375), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  OR2_X1    g0995(.A1(G390), .A2(G387), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT120), .ZN(new_n1198));
  OR4_X1    g0998(.A1(G381), .A2(new_n1195), .A3(new_n1196), .A4(new_n1198), .ZN(G407));
  OAI211_X1 g0999(.A(G407), .B(G213), .C1(G343), .C2(new_n1195), .ZN(G409));
  NAND2_X1  g1000(.A1(G390), .A2(G387), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1196), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(G393), .B(new_n778), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT125), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1203), .B(new_n1204), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(new_n1196), .A3(new_n1201), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G213), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(G343), .ZN(new_n1211));
  OAI21_X1  g1011(.A(KEYINPUT57), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n682), .B1(new_n1161), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT117), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1156), .A2(new_n1150), .A3(new_n682), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1162), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1149), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1216), .B(new_n1217), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1044), .A2(new_n1160), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1221), .A2(new_n1151), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1222), .A2(new_n948), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n718), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1135), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1191), .A2(new_n1192), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1211), .B1(new_n1220), .B2(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(G384), .B(KEYINPUT123), .Z(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1059), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1160), .A2(new_n1151), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT122), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT122), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1184), .B(new_n1234), .C1(new_n1230), .C2(new_n1059), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n681), .B1(new_n1232), .B2(KEYINPUT60), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1229), .B1(new_n1237), .B2(new_n1183), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(G384), .A2(KEYINPUT123), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(new_n1183), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT62), .B1(new_n1227), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT126), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1225), .B1(new_n1222), .B2(new_n948), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1099), .A2(KEYINPUT121), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n1190), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1163), .B2(G378), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1244), .B1(new_n1248), .B2(new_n1211), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1220), .A2(new_n1226), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1211), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(KEYINPUT126), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1242), .A2(KEYINPUT62), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1243), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1239), .A2(G2897), .A3(new_n1211), .A4(new_n1241), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1211), .A2(G2897), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1241), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n1238), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1249), .A2(new_n1252), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1209), .B1(new_n1255), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1242), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1260), .A2(new_n1266), .A3(KEYINPUT124), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT124), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n1227), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT61), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1227), .A2(new_n1242), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1265), .A2(new_n1271), .A3(new_n1272), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1264), .A2(new_n1276), .ZN(G405));
  OAI21_X1  g1077(.A(new_n1220), .B1(new_n1163), .B2(new_n1193), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT127), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1278), .B(new_n1279), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1209), .B(new_n1280), .ZN(G402));
endmodule


