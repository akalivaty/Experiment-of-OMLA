//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT74), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G143), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(new_n190), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n193), .A2(KEYINPUT65), .A3(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT65), .B1(new_n193), .B2(new_n194), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n190), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n192), .B2(new_n190), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n199), .B(G146), .C1(new_n203), .C2(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n201), .A2(KEYINPUT0), .A3(new_n206), .A4(G128), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n197), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT11), .A2(G134), .ZN(new_n211));
  OR2_X1    g025(.A1(KEYINPUT68), .A2(G137), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT68), .A2(G137), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(G137), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n221));
  INV_X1    g035(.A(new_n211), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT68), .A2(G137), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT68), .A2(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n218), .A4(new_n217), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n220), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(KEYINPUT69), .B(G131), .C1(new_n214), .C2(new_n219), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT70), .B1(new_n210), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G128), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n193), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n201), .A2(new_n236), .A3(new_n206), .A4(G128), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n216), .A2(G137), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n223), .A2(new_n224), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n216), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n242));
  OR3_X1    g056(.A1(new_n241), .A2(new_n242), .A3(new_n226), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n241), .B2(new_n226), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n238), .A2(new_n243), .A3(new_n227), .A4(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n207), .B(KEYINPUT67), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n230), .A4(new_n197), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n232), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT30), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n230), .B(new_n197), .C1(new_n208), .C2(new_n209), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n245), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(new_n250), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G119), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G116), .ZN(new_n257));
  INV_X1    g071(.A(G116), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G119), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT2), .B(G113), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n251), .A2(new_n255), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n262), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n252), .A2(new_n245), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G237), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G210), .ZN(new_n268));
  INV_X1    g082(.A(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n270), .B(new_n271), .Z(new_n272));
  NAND3_X1  g086(.A1(new_n263), .A2(new_n265), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT31), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n263), .A2(new_n275), .A3(new_n265), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n272), .B(KEYINPUT72), .Z(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AND4_X1   g093(.A1(new_n227), .A2(new_n238), .A3(new_n243), .A4(new_n244), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n252), .B2(KEYINPUT70), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n264), .B1(new_n281), .B2(new_n248), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n265), .B1(new_n282), .B2(KEYINPUT73), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n249), .A2(KEYINPUT73), .A3(new_n262), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT28), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n265), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n279), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(KEYINPUT32), .B(new_n189), .C1(new_n277), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n288), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n249), .A2(new_n262), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n265), .A3(new_n284), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n296), .B2(KEYINPUT28), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n274), .B(new_n276), .C1(new_n297), .C2(new_n279), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT32), .B1(new_n298), .B2(new_n189), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n286), .A2(new_n288), .A3(new_n279), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n263), .A2(new_n265), .ZN(new_n302));
  INV_X1    g116(.A(new_n272), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT29), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n252), .A2(new_n245), .A3(new_n264), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n264), .B1(new_n252), .B2(new_n245), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT28), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n310), .B2(new_n288), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n288), .A2(new_n307), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n272), .A2(KEYINPUT29), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n306), .B1(new_n315), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  INV_X1    g131(.A(new_n309), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n265), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n292), .B1(new_n319), .B2(KEYINPUT28), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n312), .B1(new_n320), .B2(new_n307), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT76), .B(new_n317), .C1(new_n321), .C2(new_n314), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n305), .A2(new_n316), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n323), .A2(new_n324), .A3(G472), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n324), .B1(new_n323), .B2(G472), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n300), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XOR2_X1   g141(.A(KEYINPUT78), .B(G217), .Z(new_n328));
  INV_X1    g142(.A(G234), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(G902), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT16), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n333), .A2(KEYINPUT16), .A3(G140), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(G146), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n334), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT80), .B1(new_n341), .B2(new_n190), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n340), .A2(new_n343), .A3(G146), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n256), .A2(KEYINPUT23), .A3(G128), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT23), .B1(new_n256), .B2(G128), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n345), .A2(new_n346), .B1(new_n256), .B2(G128), .ZN(new_n347));
  INV_X1    g161(.A(G110), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g163(.A(G119), .B(G128), .Z(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT24), .B(G110), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI221_X1 g166(.A(new_n339), .B1(new_n342), .B2(new_n344), .C1(new_n349), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n335), .A2(new_n336), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n190), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n337), .ZN(new_n356));
  OAI221_X1 g170(.A(new_n356), .B1(new_n348), .B2(new_n347), .C1(new_n350), .C2(new_n351), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT22), .B(G137), .ZN(new_n359));
  INV_X1    g173(.A(G221), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n360), .A2(new_n329), .A3(G953), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n359), .B(new_n361), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n357), .A3(new_n362), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n317), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n367), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n330), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n372));
  AOI21_X1  g186(.A(G902), .B1(new_n328), .B2(new_n329), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n364), .A2(new_n365), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n374), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT81), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(G469), .A2(G902), .ZN(new_n379));
  INV_X1    g193(.A(G469), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT82), .B(G107), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n382), .A2(KEYINPUT3), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT3), .B1(new_n382), .B2(G107), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(G104), .B2(new_n386), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n384), .A2(new_n387), .A3(G101), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n382), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(G104), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n269), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n238), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n201), .A2(new_n206), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n236), .B1(new_n192), .B2(new_n190), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n394), .B1(new_n233), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n237), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n392), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n231), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT12), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n269), .A2(KEYINPUT83), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n384), .B2(new_n387), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n386), .A2(G104), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(KEYINPUT3), .B2(new_n390), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n412), .B(new_n269), .C1(new_n381), .C2(new_n383), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n407), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n381), .B2(new_n383), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT4), .B1(new_n415), .B2(new_n409), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n406), .B1(new_n210), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n413), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT4), .ZN(new_n420));
  INV_X1    g234(.A(new_n416), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n422), .A2(new_n246), .A3(KEYINPUT84), .A4(new_n197), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT10), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n398), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n238), .A2(new_n392), .A3(KEYINPUT10), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n428), .A3(new_n231), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G140), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n267), .A2(G227), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n430), .B(new_n431), .Z(new_n432));
  AND3_X1   g246(.A1(new_n405), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n428), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n230), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n432), .B1(new_n435), .B2(new_n429), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n380), .B(new_n317), .C1(new_n433), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n405), .A2(new_n429), .ZN(new_n438));
  INV_X1    g252(.A(new_n432), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n426), .A2(new_n427), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n418), .B2(new_n423), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n439), .B1(new_n442), .B2(new_n231), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n435), .B1(new_n443), .B2(KEYINPUT86), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n445), .B(new_n439), .C1(new_n442), .C2(new_n231), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n440), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n379), .B(new_n437), .C1(new_n447), .C2(new_n380), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT9), .B(G234), .Z(new_n449));
  AOI21_X1  g263(.A(new_n360), .B1(new_n449), .B2(new_n317), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n356), .ZN(new_n453));
  INV_X1    g267(.A(G214), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n454), .A2(G237), .A3(G953), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G143), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n192), .B2(new_n455), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT17), .A3(G131), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(G131), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n456), .B(new_n226), .C1(new_n192), .C2(new_n455), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n453), .B(new_n458), .C1(new_n461), .C2(KEYINPUT17), .ZN(new_n462));
  OAI22_X1  g276(.A1(new_n342), .A2(new_n344), .B1(new_n190), .B2(new_n341), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n457), .A2(KEYINPUT18), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n457), .A2(KEYINPUT18), .A3(G131), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .A4(new_n460), .ZN(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n382), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT93), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n462), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n462), .A2(new_n466), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n317), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n474), .A2(G475), .ZN(new_n475));
  NOR2_X1   g289(.A1(G475), .A2(G902), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n337), .A2(new_n338), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n337), .A2(new_n338), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT91), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT19), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n478), .A2(new_n479), .B1(new_n482), .B2(new_n190), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n461), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n190), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n339), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n466), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n468), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n477), .B(new_n470), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT94), .B1(new_n491), .B2(new_n471), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n476), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT20), .ZN(new_n494));
  INV_X1    g308(.A(new_n476), .ZN(new_n495));
  AOI211_X1 g309(.A(KEYINPUT20), .B(new_n495), .C1(new_n491), .C2(new_n471), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n475), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT100), .ZN(new_n499));
  INV_X1    g313(.A(G952), .ZN(new_n500));
  AOI211_X1 g314(.A(G953), .B(new_n500), .C1(G234), .C2(G237), .ZN(new_n501));
  XOR2_X1   g315(.A(KEYINPUT21), .B(G898), .Z(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n317), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n204), .A2(G128), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n216), .B(new_n508), .C1(new_n192), .C2(new_n233), .ZN(new_n509));
  INV_X1    g323(.A(G122), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G116), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n258), .A2(G122), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n513), .A2(new_n381), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n381), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n202), .A2(G143), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n233), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT95), .B1(new_n519), .B2(KEYINPUT13), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n507), .B1(new_n519), .B2(KEYINPUT13), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n523), .C1(new_n192), .C2(new_n233), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n516), .B1(new_n525), .B2(G134), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n510), .A2(G116), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT14), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n511), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT96), .B(new_n511), .C1(new_n528), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n529), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G107), .ZN(new_n536));
  OAI21_X1  g350(.A(G134), .B1(new_n519), .B2(new_n507), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n515), .B1(new_n537), .B2(new_n509), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n328), .A2(new_n449), .A3(new_n267), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n527), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n536), .A2(new_n538), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n540), .B1(new_n543), .B2(new_n526), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT97), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n527), .A2(new_n546), .A3(new_n539), .A4(new_n541), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n317), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G478), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT98), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(KEYINPUT98), .A3(new_n550), .ZN(new_n554));
  INV_X1    g368(.A(new_n550), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n545), .A2(new_n317), .A3(new_n547), .A4(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n556), .A2(KEYINPUT99), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(KEYINPUT99), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n553), .A2(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n498), .A2(new_n499), .A3(new_n506), .A4(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n475), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT20), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n339), .A2(new_n486), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT92), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n483), .A2(new_n484), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n461), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n468), .B1(new_n566), .B2(new_n466), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n477), .B1(new_n567), .B2(new_n470), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n491), .A2(KEYINPUT94), .A3(new_n471), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n562), .B1(new_n570), .B2(new_n476), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n561), .B1(new_n571), .B2(new_n496), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n553), .A2(new_n554), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n557), .A2(new_n558), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n506), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT100), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n560), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G210), .B1(G237), .B2(G902), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT90), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n260), .A2(new_n261), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n581), .A2(G113), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT5), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n392), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT88), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT88), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n392), .A2(new_n587), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT87), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n422), .B2(new_n262), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n590), .B(new_n262), .C1(new_n414), .C2(new_n416), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n589), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(G110), .B(G122), .Z(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n595), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n597), .B(new_n589), .C1(new_n591), .C2(new_n593), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(KEYINPUT6), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n210), .A2(G125), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n235), .A2(new_n333), .A3(new_n237), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G224), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G953), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n602), .B(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT6), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n594), .A2(new_n606), .A3(new_n595), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n599), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n584), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n609), .B(KEYINPUT89), .C1(new_n388), .C2(new_n391), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT89), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n611), .B1(new_n392), .B2(new_n584), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n585), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n595), .B(KEYINPUT8), .Z(new_n614));
  AOI22_X1  g428(.A1(new_n602), .A2(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n604), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n600), .A2(KEYINPUT7), .A3(new_n616), .A4(new_n601), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT7), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n602), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n615), .A2(new_n598), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n317), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n579), .B1(new_n608), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n620), .A2(new_n317), .ZN(new_n623));
  INV_X1    g437(.A(new_n579), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n599), .A2(new_n605), .A3(new_n607), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G214), .B1(G237), .B2(G902), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n452), .A2(new_n577), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n327), .A2(new_n378), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  NAND2_X1  g447(.A1(new_n548), .A2(new_n549), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT33), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n545), .A2(new_n547), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n635), .B1(new_n636), .B2(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n317), .A2(G478), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n572), .A2(new_n506), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n578), .B1(new_n608), .B2(new_n621), .ZN(new_n641));
  INV_X1    g455(.A(new_n578), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n623), .A2(new_n642), .A3(new_n625), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n641), .A2(new_n628), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  OR3_X1    g459(.A1(new_n640), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n645), .B1(new_n640), .B2(new_n644), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n378), .A2(new_n448), .A3(new_n451), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n298), .A2(new_n189), .ZN(new_n650));
  INV_X1    g464(.A(G472), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n298), .B2(new_n317), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  INV_X1    g470(.A(new_n559), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n657), .A2(new_n641), .A3(new_n628), .A4(new_n643), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n570), .A2(new_n562), .A3(new_n476), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n494), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n561), .A3(new_n506), .ZN(new_n662));
  OR3_X1    g476(.A1(new_n658), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n659), .B1(new_n658), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n653), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NOR2_X1   g482(.A1(new_n363), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n358), .B(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n373), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n370), .A2(new_n671), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n452), .A2(new_n577), .A3(new_n630), .A4(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n650), .A2(new_n652), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n501), .B1(new_n504), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AOI211_X1 g494(.A(KEYINPUT20), .B(new_n495), .C1(new_n568), .C2(new_n569), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n561), .B(new_n680), .C1(new_n571), .C2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n559), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n448), .A2(new_n451), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n644), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n327), .A2(new_n672), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  INV_X1    g501(.A(new_n302), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n688), .A2(new_n272), .B1(new_n278), .B2(new_n319), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n689), .B2(G902), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n300), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n679), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n452), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n627), .B(KEYINPUT38), .ZN(new_n697));
  OR4_X1    g511(.A1(new_n629), .A2(new_n498), .A3(new_n672), .A4(new_n559), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n691), .A2(new_n695), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(new_n192), .Z(G45));
  NAND2_X1  g515(.A1(new_n572), .A2(new_n639), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n679), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n327), .A2(new_n672), .A3(new_n685), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  INV_X1    g519(.A(new_n436), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n443), .A2(new_n405), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n380), .B1(new_n708), .B2(new_n317), .ZN(new_n709));
  INV_X1    g523(.A(new_n437), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n451), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n327), .A2(new_n378), .A3(new_n648), .A4(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT41), .B(G113), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT104), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n714), .B(new_n716), .ZN(G15));
  NAND4_X1  g531(.A1(new_n327), .A2(new_n378), .A3(new_n665), .A4(new_n713), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  INV_X1    g533(.A(new_n644), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n451), .A2(new_n577), .A3(new_n720), .A4(new_n711), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n327), .A2(new_n721), .A3(new_n672), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  INV_X1    g537(.A(new_n658), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n572), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n712), .A3(new_n505), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n370), .A2(new_n376), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n321), .A2(new_n278), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n274), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n728), .A2(KEYINPUT106), .A3(new_n274), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n732), .A3(new_n276), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n188), .B(KEYINPUT105), .Z(new_n734));
  AOI21_X1  g548(.A(new_n652), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n726), .A2(new_n727), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NOR2_X1   g551(.A1(new_n712), .A2(new_n644), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n735), .A3(new_n672), .A4(new_n703), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  NAND3_X1  g554(.A1(new_n622), .A2(new_n628), .A3(new_n626), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n684), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n327), .A2(new_n378), .A3(new_n703), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n742), .A2(KEYINPUT42), .A3(new_n703), .ZN(new_n746));
  INV_X1    g560(.A(new_n299), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(KEYINPUT107), .A3(new_n290), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n325), .B2(new_n326), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n300), .A2(KEYINPUT107), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n727), .B(new_n746), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  NAND4_X1  g567(.A1(new_n327), .A2(new_n378), .A3(new_n683), .A4(new_n742), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NAND2_X1  g569(.A1(new_n498), .A2(new_n639), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n758), .B(new_n672), .C1(new_n650), .C2(new_n652), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n380), .B1(new_n447), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n764), .B2(new_n447), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n379), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n437), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT46), .B1(new_n766), .B2(new_n379), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n451), .B(new_n693), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n741), .B(KEYINPUT108), .Z(new_n771));
  NOR4_X1   g585(.A1(new_n761), .A2(new_n763), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(G137), .Z(G39));
  OAI21_X1  g587(.A(new_n451), .B1(new_n768), .B2(new_n769), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT47), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n774), .A2(KEYINPUT47), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n327), .ZN(new_n779));
  INV_X1    g593(.A(new_n378), .ZN(new_n780));
  INV_X1    g594(.A(new_n741), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n703), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  NAND4_X1  g600(.A1(new_n735), .A2(new_n672), .A3(new_n703), .A4(new_n742), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n682), .A2(new_n657), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n781), .A2(KEYINPUT112), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n661), .A2(new_n561), .A3(new_n559), .A4(new_n680), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n790), .B1(new_n791), .B2(new_n741), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n789), .A2(new_n452), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n327), .A2(new_n793), .A3(new_n672), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n754), .A2(new_n787), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n702), .B1(new_n572), .B2(new_n559), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n630), .A2(new_n796), .A3(new_n506), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n673), .A2(new_n674), .B1(new_n653), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n632), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n714), .A2(new_n718), .A3(new_n722), .A4(new_n736), .ZN(new_n801));
  AND4_X1   g615(.A1(KEYINPUT53), .A2(new_n800), .A3(new_n752), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n725), .A2(new_n684), .A3(new_n672), .A4(new_n679), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n691), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n686), .A2(new_n704), .A3(new_n805), .A4(new_n739), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n802), .A2(new_n803), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n806), .B(KEYINPUT52), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT53), .A4(new_n752), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  INV_X1    g628(.A(new_n799), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n754), .A2(new_n787), .A3(new_n794), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n801), .A2(new_n752), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT113), .A4(new_n752), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n810), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n813), .B(new_n814), .C1(KEYINPUT53), .C2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n819), .A2(new_n820), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n824), .B2(new_n808), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n822), .B1(new_n826), .B2(new_n814), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n735), .A2(new_n727), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n758), .A2(new_n501), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n628), .B1(KEYINPUT116), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(new_n697), .A3(new_n713), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n834), .B(new_n835), .Z(new_n836));
  NAND2_X1  g650(.A1(new_n713), .A2(new_n781), .ZN(new_n837));
  INV_X1    g651(.A(new_n501), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n837), .A2(new_n691), .A3(new_n780), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n572), .A2(new_n639), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n829), .A2(new_n713), .A3(new_n781), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n735), .A2(new_n672), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n839), .A2(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n836), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n778), .B1(new_n450), .B2(new_n711), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n830), .A2(new_n771), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n846), .B2(KEYINPUT117), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n845), .B(KEYINPUT51), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n727), .B1(new_n749), .B2(new_n750), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n851), .A2(new_n841), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT48), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  INV_X1    g669(.A(new_n839), .ZN(new_n856));
  OAI211_X1 g670(.A(G952), .B(new_n267), .C1(new_n856), .C2(new_n702), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n738), .B2(new_n831), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n850), .A2(new_n854), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n778), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(KEYINPUT115), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  INV_X1    g676(.A(new_n711), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n778), .A2(new_n862), .B1(new_n451), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n848), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT51), .B1(new_n845), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n827), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(G952), .A2(G953), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n697), .B1(KEYINPUT49), .B2(new_n863), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n727), .A2(new_n451), .A3(new_n628), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n756), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT49), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n871), .B1(new_n872), .B2(new_n711), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n869), .B1(KEYINPUT111), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(KEYINPUT111), .B2(new_n873), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n867), .A2(new_n868), .B1(new_n691), .B2(new_n875), .ZN(G75));
  NOR2_X1   g690(.A1(new_n267), .A2(G952), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n599), .A2(new_n607), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n605), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT55), .Z(new_n880));
  OAI21_X1  g694(.A(new_n813), .B1(KEYINPUT53), .B2(new_n821), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(G210), .A3(G902), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n880), .B1(new_n884), .B2(KEYINPUT118), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n882), .A2(new_n887), .A3(new_n883), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n877), .B(new_n885), .C1(new_n889), .C2(new_n880), .ZN(G51));
  AOI21_X1  g704(.A(new_n803), .B1(new_n802), .B2(new_n808), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT114), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n893), .B2(new_n825), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(KEYINPUT119), .A3(new_n822), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n893), .A2(new_n825), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n897), .A3(new_n814), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n379), .B(KEYINPUT57), .Z(new_n899));
  NAND3_X1  g713(.A1(new_n895), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n895), .A2(new_n898), .A3(new_n902), .A4(new_n899), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n708), .A3(new_n903), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n896), .A2(new_n317), .A3(new_n766), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n877), .B1(new_n904), .B2(new_n905), .ZN(G54));
  NAND4_X1  g720(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n907));
  INV_X1    g721(.A(new_n570), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n877), .ZN(G60));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT59), .Z(new_n913));
  NOR2_X1   g727(.A1(new_n637), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n895), .A2(new_n898), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n827), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n877), .B1(new_n919), .B2(new_n637), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n915), .A2(new_n916), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(G63));
  XOR2_X1   g736(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n923));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n881), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n364), .A2(new_n365), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n877), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n881), .A2(new_n925), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n670), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n929), .B2(new_n670), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(KEYINPUT61), .B(new_n928), .C1(new_n931), .C2(new_n932), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(G66));
  NAND2_X1  g751(.A1(new_n801), .A2(new_n815), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n267), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n503), .B2(new_n603), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n878), .B1(G898), .B2(new_n267), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT124), .Z(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n796), .A2(new_n781), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n779), .A2(new_n780), .A3(new_n694), .A4(new_n946), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n947), .B(new_n772), .C1(new_n778), .C2(new_n784), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n686), .A2(new_n704), .A3(new_n739), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n700), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n948), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n948), .B2(new_n954), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n267), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n251), .A2(new_n255), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n482), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n772), .B1(new_n778), .B2(new_n784), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n965), .A2(new_n752), .A3(new_n754), .A4(new_n950), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n851), .A2(new_n725), .A3(new_n770), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT126), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n964), .B1(new_n969), .B2(new_n267), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n945), .B1(new_n962), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n962), .A2(new_n945), .A3(new_n971), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n974), .ZN(new_n977));
  AOI211_X1 g791(.A(KEYINPUT127), .B(new_n970), .C1(new_n959), .C2(new_n961), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n972), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(G72));
  NAND2_X1  g794(.A1(G472), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT63), .Z(new_n982));
  OR2_X1    g796(.A1(new_n957), .A2(new_n958), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n938), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n688), .A2(new_n303), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n982), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n302), .A2(new_n272), .ZN(new_n988));
  NOR4_X1   g802(.A1(new_n826), .A2(new_n987), .A3(new_n985), .A4(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n969), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n982), .B1(new_n990), .B2(new_n938), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n991), .A2(new_n988), .ZN(new_n992));
  NOR4_X1   g806(.A1(new_n986), .A2(new_n877), .A3(new_n989), .A4(new_n992), .ZN(G57));
endmodule


