//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT84), .ZN(new_n188));
  XNOR2_X1  g002(.A(G113), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT18), .A2(G131), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G237), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G953), .ZN(new_n197));
  INV_X1    g011(.A(G953), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT67), .ZN(new_n199));
  OAI211_X1 g013(.A(G214), .B(new_n195), .C1(new_n197), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(KEYINPUT67), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(G953), .ZN(new_n204));
  AOI21_X1  g018(.A(G237), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(G143), .B1(new_n205), .B2(G214), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT82), .B1(new_n202), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n200), .A2(new_n201), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(G143), .A3(G214), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n194), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n211), .A2(new_n194), .ZN(new_n213));
  XNOR2_X1  g027(.A(G125), .B(G140), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n212), .A2(new_n213), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(KEYINPUT16), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT16), .ZN(new_n221));
  INV_X1    g035(.A(G140), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G125), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT71), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT71), .A4(G125), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n220), .A2(G146), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n214), .A2(KEYINPUT83), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT19), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n214), .A2(KEYINPUT83), .A3(KEYINPUT19), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n227), .B1(new_n232), .B2(G146), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT64), .A2(G131), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT64), .A2(G131), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n202), .B2(new_n206), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n234), .A2(new_n235), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n208), .A2(new_n238), .A3(new_n210), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n233), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n188), .B(new_n192), .C1(new_n219), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT17), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n237), .A2(new_n242), .A3(new_n239), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT85), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n220), .A2(new_n225), .A3(new_n226), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n215), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n227), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n238), .B1(new_n208), .B2(new_n210), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(KEYINPUT17), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n237), .A2(KEYINPUT85), .A3(new_n242), .A4(new_n239), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n207), .A2(new_n211), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n193), .ZN(new_n254));
  INV_X1    g068(.A(new_n213), .ZN(new_n255));
  INV_X1    g069(.A(new_n218), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n257), .A3(new_n191), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n241), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n237), .A2(new_n239), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n260), .B(new_n227), .C1(G146), .C2(new_n232), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n188), .B1(new_n262), .B2(new_n192), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n187), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT20), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT86), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT86), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n267), .A3(KEYINPUT20), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n219), .A2(new_n240), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT84), .B1(new_n269), .B2(new_n191), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n258), .A3(new_n241), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT20), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n187), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n266), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n201), .A2(G128), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT89), .ZN(new_n276));
  INV_X1    g090(.A(G128), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(G143), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(G134), .ZN(new_n279));
  INV_X1    g093(.A(G107), .ZN(new_n280));
  INV_X1    g094(.A(G116), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G122), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n280), .B1(new_n283), .B2(KEYINPUT14), .ZN(new_n284));
  XNOR2_X1  g098(.A(G116), .B(G122), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT14), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n284), .A2(new_n287), .B1(new_n280), .B2(new_n285), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT9), .B(G234), .Z(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G217), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n291), .A2(new_n292), .A3(G953), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n285), .B(new_n280), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(KEYINPUT88), .ZN(new_n295));
  INV_X1    g109(.A(G134), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT13), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n276), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n298), .A2(new_n278), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n278), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n289), .A2(new_n293), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n293), .B1(new_n289), .B2(new_n301), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  INV_X1    g119(.A(G478), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n306), .A2(KEYINPUT15), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n304), .B2(new_n305), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(G234), .A2(G237), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n312), .A2(G952), .A3(new_n198), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n203), .A2(new_n204), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n315), .A2(G902), .A3(new_n312), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT21), .B(G898), .Z(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n313), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n252), .A2(new_n257), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n192), .A2(KEYINPUT87), .ZN(new_n322));
  AOI21_X1  g136(.A(G902), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n321), .B2(new_n322), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G475), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n274), .A2(new_n311), .A3(new_n320), .A4(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n277), .A2(KEYINPUT1), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n215), .A2(G143), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n201), .A2(G146), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n277), .A2(new_n215), .A3(G143), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n201), .B(G146), .C1(new_n277), .C2(KEYINPUT1), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  XNOR2_X1  g150(.A(G143), .B(G146), .ZN(new_n337));
  NAND2_X1  g151(.A1(KEYINPUT0), .A2(G128), .ZN(new_n338));
  OR2_X1    g152(.A1(KEYINPUT0), .A2(G128), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n337), .A2(new_n338), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n336), .B1(G125), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT78), .ZN(new_n344));
  INV_X1    g158(.A(G224), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G953), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n344), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT6), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n280), .A3(G104), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT73), .B1(new_n280), .B2(G104), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n190), .A3(G107), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n349), .A2(new_n353), .A3(new_n351), .A4(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(G101), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n363));
  INV_X1    g177(.A(new_n359), .ZN(new_n364));
  INV_X1    g178(.A(G101), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n361), .A2(new_n366), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n358), .A2(new_n360), .A3(new_n363), .A4(G101), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT75), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT2), .A2(G113), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT66), .ZN(new_n373));
  OR2_X1    g187(.A1(KEYINPUT2), .A2(G113), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G116), .B(G119), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n380));
  INV_X1    g194(.A(G119), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G116), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n380), .B(G113), .C1(KEYINPUT5), .C2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n190), .A2(G107), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n280), .A2(G104), .ZN(new_n387));
  OAI21_X1  g201(.A(G101), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n359), .B2(G101), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT76), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(new_n388), .C1(new_n359), .C2(G101), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n385), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(G110), .B(G122), .Z(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n379), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n395), .B(KEYINPUT77), .Z(new_n398));
  NAND2_X1  g212(.A1(new_n361), .A2(new_n366), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT75), .A3(new_n369), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n377), .B1(new_n400), .B2(new_n367), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n398), .B1(new_n401), .B2(new_n393), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n348), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n379), .A2(new_n394), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT6), .B1(new_n404), .B2(new_n398), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n347), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n395), .B(KEYINPUT8), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n385), .A2(new_n389), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n394), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n401), .A2(new_n393), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(new_n396), .ZN(new_n411));
  INV_X1    g225(.A(new_n346), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n343), .B1(KEYINPUT7), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n342), .ZN(new_n414));
  INV_X1    g228(.A(G125), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT79), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT7), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n346), .B2(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n413), .A2(new_n416), .B1(new_n343), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n411), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n406), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n328), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n406), .A2(new_n423), .A3(new_n421), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n406), .A2(new_n423), .A3(new_n421), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT81), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n423), .B1(new_n406), .B2(new_n421), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT80), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n424), .A2(new_n427), .A3(new_n429), .A4(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G469), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n342), .B1(new_n400), .B2(new_n367), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n390), .A2(new_n392), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT10), .A3(new_n335), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n389), .A2(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n438), .A2(KEYINPUT10), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT11), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n296), .B2(G137), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n296), .A2(G137), .ZN(new_n443));
  INV_X1    g257(.A(G137), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT11), .A3(G134), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G131), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT65), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n238), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n446), .A2(KEYINPUT65), .A3(new_n236), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n434), .A2(new_n440), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n390), .A2(new_n437), .A3(new_n392), .ZN(new_n454));
  INV_X1    g268(.A(new_n438), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT12), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT12), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n444), .A2(KEYINPUT11), .A3(G134), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT11), .B1(new_n444), .B2(G134), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n461), .A2(new_n448), .A3(new_n238), .A4(new_n443), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT65), .B1(new_n446), .B2(new_n236), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n462), .A2(new_n463), .B1(G131), .B2(new_n446), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n458), .B(new_n464), .C1(new_n454), .C2(new_n455), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n314), .A2(G227), .ZN(new_n467));
  XNOR2_X1  g281(.A(G110), .B(G140), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n453), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n371), .A2(new_n414), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n436), .A2(new_n439), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n464), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n452), .B1(new_n434), .B2(new_n440), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n433), .B(new_n305), .C1(new_n471), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(G469), .A2(G902), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n470), .B1(new_n453), .B2(new_n466), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n475), .A3(new_n469), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(G469), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G221), .B1(new_n291), .B2(G902), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G214), .B1(G237), .B2(G902), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n327), .A2(new_n432), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G472), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n452), .A2(new_n414), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n444), .A2(G134), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n443), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n491), .A2(G131), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n335), .B(new_n493), .C1(new_n450), .C2(new_n451), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n377), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(KEYINPUT28), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n492), .B(new_n437), .C1(new_n462), .C2(new_n463), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n462), .A2(new_n463), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n342), .B1(new_n499), .B2(new_n447), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n378), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n495), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n497), .B1(new_n502), .B2(KEYINPUT28), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n365), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n205), .A2(G210), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT29), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT30), .B1(new_n498), .B2(new_n500), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n494), .B(new_n511), .C1(new_n464), .C2(new_n342), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n496), .B1(new_n513), .B2(new_n378), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n507), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n503), .A2(KEYINPUT29), .A3(new_n508), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n488), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT68), .B1(new_n514), .B2(new_n508), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n377), .B1(new_n510), .B2(new_n512), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n523));
  NOR4_X1   g337(.A1(new_n522), .A2(new_n523), .A3(new_n496), .A4(new_n507), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT31), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n502), .A2(KEYINPUT28), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n507), .B1(new_n526), .B2(new_n497), .ZN(new_n527));
  INV_X1    g341(.A(new_n512), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n511), .B1(new_n489), .B2(new_n494), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n378), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n495), .A4(new_n508), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT69), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n514), .A2(new_n534), .A3(new_n531), .A4(new_n508), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n525), .A2(new_n527), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT32), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n520), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n314), .A2(G221), .A3(G234), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT22), .Z(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(new_n444), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n277), .A2(G119), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n381), .A2(G128), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT24), .B(G110), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G110), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n546), .A2(KEYINPUT23), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(KEYINPUT70), .A3(new_n545), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT70), .ZN(new_n553));
  OAI211_X1 g367(.A(G119), .B(new_n277), .C1(new_n553), .C2(KEYINPUT23), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n248), .B(new_n549), .C1(new_n550), .C2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT72), .B(G110), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n547), .A2(new_n548), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n227), .B(new_n217), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n544), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n556), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n543), .B(G137), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n564), .A3(new_n305), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n292), .B1(G234), .B2(new_n305), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT25), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n565), .B(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n569), .B2(new_n566), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n541), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n487), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(new_n365), .ZN(G3));
  NAND2_X1  g387(.A1(new_n536), .A2(new_n538), .ZN(new_n574));
  INV_X1    g388(.A(new_n527), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n530), .A2(new_n495), .A3(new_n508), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n523), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n514), .A2(KEYINPUT68), .A3(new_n508), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n579), .B2(KEYINPUT31), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n533), .A2(new_n535), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n574), .B1(new_n583), .B2(new_n488), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n482), .A2(new_n570), .A3(new_n483), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT90), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n585), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n531), .B1(new_n577), .B2(new_n578), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n588), .A2(new_n581), .A3(new_n575), .ZN(new_n589));
  OAI21_X1  g403(.A(G472), .B1(new_n589), .B2(G902), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT90), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n587), .A2(new_n590), .A3(new_n591), .A4(new_n574), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n486), .B1(new_n425), .B2(new_n430), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT91), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n304), .A2(new_n305), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n306), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT92), .B1(new_n302), .B2(new_n303), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(KEYINPUT92), .B(KEYINPUT33), .C1(new_n302), .C2(new_n303), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G478), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n274), .A2(new_n325), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT91), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n605), .B(new_n486), .C1(new_n425), .C2(new_n430), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n595), .A2(new_n604), .A3(new_n320), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n593), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT34), .B(G104), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  INV_X1    g424(.A(new_n325), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n264), .A2(new_n267), .A3(KEYINPUT20), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n267), .B1(new_n264), .B2(KEYINPUT20), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n273), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n271), .A2(KEYINPUT93), .A3(new_n272), .A4(new_n187), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n311), .B(new_n611), .C1(new_n614), .C2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n619), .A2(new_n320), .A3(new_n606), .A4(new_n595), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n593), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT35), .B(G107), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  INV_X1    g437(.A(new_n486), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n430), .B(new_n328), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n428), .B(new_n426), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n569), .A2(new_n566), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(new_n562), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n630), .B(new_n305), .C1(new_n292), .C2(G234), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n590), .A2(new_n574), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n627), .A2(new_n485), .A3(new_n633), .A4(new_n327), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT37), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n550), .ZN(G12));
  NAND3_X1  g450(.A1(new_n595), .A2(new_n606), .A3(new_n632), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n538), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT32), .B1(new_n589), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n519), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n484), .ZN(new_n643));
  INV_X1    g457(.A(new_n311), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n614), .A2(new_n618), .ZN(new_n645));
  INV_X1    g459(.A(new_n316), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT94), .B(G900), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n648), .A2(KEYINPUT95), .ZN(new_n649));
  INV_X1    g463(.A(new_n313), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(KEYINPUT95), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n644), .A2(new_n645), .A3(new_n325), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n638), .A2(new_n643), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  XNOR2_X1  g469(.A(new_n432), .B(KEYINPUT38), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n652), .B(KEYINPUT39), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n485), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n656), .A2(new_n486), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n640), .A2(new_n641), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n577), .A2(new_n578), .B1(new_n502), .B2(new_n507), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n662), .B2(G902), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n632), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n311), .B1(new_n274), .B2(new_n325), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n660), .A2(new_n664), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G143), .ZN(G45));
  NAND2_X1  g482(.A1(new_n274), .A2(new_n325), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n603), .A2(new_n597), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n652), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n638), .A2(new_n643), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT96), .B(G146), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G48));
  NAND2_X1  g490(.A1(new_n474), .A2(new_n475), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n470), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n474), .B(new_n469), .C1(new_n465), .C2(new_n457), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n305), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G469), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n483), .A3(new_n477), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n541), .A2(new_n570), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n607), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT97), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT41), .B(G113), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NOR2_X1   g503(.A1(new_n620), .A2(new_n685), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n281), .ZN(G18));
  NAND3_X1  g505(.A1(new_n541), .A2(new_n327), .A3(new_n684), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n637), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n381), .ZN(G21));
  NAND4_X1  g508(.A1(new_n595), .A2(new_n666), .A3(new_n684), .A4(new_n606), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n538), .B(KEYINPUT98), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n536), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n590), .A2(new_n570), .A3(new_n320), .A4(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(G122), .Z(G24));
  NAND3_X1  g514(.A1(new_n590), .A2(new_n632), .A3(new_n697), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n671), .A3(new_n672), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n595), .A2(new_n606), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n683), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT99), .B(G125), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G27));
  NAND2_X1  g521(.A1(new_n482), .A2(KEYINPUT100), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT100), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n477), .A2(new_n709), .A3(new_n478), .A4(new_n481), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n483), .A3(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n432), .A2(new_n711), .A3(new_n624), .ZN(new_n712));
  INV_X1    g526(.A(new_n570), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n642), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n714), .A3(new_n673), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n712), .A2(new_n714), .A3(KEYINPUT42), .A4(new_n673), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  NAND3_X1  g534(.A1(new_n712), .A2(new_n714), .A3(new_n653), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT101), .B(G134), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G36));
  NAND3_X1  g537(.A1(new_n274), .A2(new_n670), .A3(new_n325), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT43), .Z(new_n725));
  OAI211_X1 g539(.A(new_n584), .B(new_n632), .C1(new_n725), .C2(KEYINPUT103), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n725), .A2(KEYINPUT103), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n432), .A2(new_n624), .ZN(new_n731));
  INV_X1    g545(.A(new_n483), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n479), .A2(new_n480), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT45), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(G469), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT46), .B1(new_n735), .B2(new_n478), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT102), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(KEYINPUT46), .A3(new_n478), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n738), .A2(new_n477), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n732), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(new_n657), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n728), .A2(new_n729), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n730), .A2(new_n731), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G137), .ZN(G39));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n740), .B1(KEYINPUT104), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n747));
  AND2_X1   g561(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n673), .A3(new_n731), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n750), .A2(new_n541), .A3(new_n570), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n222), .ZN(G42));
  NOR2_X1   g566(.A1(G952), .A2(G953), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT114), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n320), .A2(new_n586), .A3(new_n627), .A4(new_n592), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n572), .B1(new_n755), .B2(new_n604), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n669), .A2(new_n311), .A3(new_n319), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n586), .A2(new_n627), .A3(new_n592), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n634), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(new_n634), .A3(KEYINPUT105), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n756), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AND4_X1   g577(.A1(new_n320), .A2(new_n619), .A3(new_n606), .A4(new_n595), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n642), .A2(new_n713), .A3(new_n683), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n642), .A2(new_n326), .A3(new_n683), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n638), .ZN(new_n767));
  OAI22_X1  g581(.A1(new_n685), .A2(new_n607), .B1(new_n695), .B2(new_n698), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI22_X1  g585(.A1(new_n620), .A2(new_n685), .B1(new_n692), .B2(new_n637), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT110), .B1(new_n772), .B2(new_n768), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n719), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(KEYINPUT111), .A3(new_n719), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n763), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n595), .A2(new_n606), .A3(new_n666), .ZN(new_n780));
  INV_X1    g594(.A(new_n711), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n664), .A3(new_n652), .A4(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n705), .A2(new_n782), .A3(new_n654), .A4(new_n674), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n637), .A2(new_n642), .A3(new_n484), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n786), .A2(new_n653), .B1(new_n704), .B2(new_n702), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT52), .A3(new_n674), .A4(new_n782), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n785), .A2(new_n788), .A3(KEYINPUT107), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n702), .A2(new_n712), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(new_n721), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n731), .A2(new_n632), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n642), .A2(new_n484), .A3(new_n611), .A4(new_n672), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n311), .A3(new_n798), .A4(new_n645), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n779), .A2(new_n794), .A3(KEYINPUT53), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n772), .A2(new_n768), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n756), .A2(new_n803), .A3(new_n761), .A4(new_n762), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n719), .A2(new_n796), .A3(new_n799), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n789), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT109), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n810), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n802), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n756), .A2(new_n803), .A3(new_n761), .A4(new_n762), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n719), .A2(new_n796), .A3(new_n799), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT106), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT53), .B1(new_n820), .B2(new_n794), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT108), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n807), .B2(new_n806), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n815), .B1(new_n823), .B2(KEYINPUT54), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n570), .A2(new_n590), .A3(new_n313), .A4(new_n697), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n725), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n684), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n703), .ZN(new_n828));
  INV_X1    g642(.A(G952), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n828), .A2(new_n829), .A3(G953), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n432), .A2(new_n650), .A3(new_n624), .A4(new_n683), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n725), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n571), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT48), .Z(new_n834));
  AND3_X1   g648(.A1(new_n661), .A2(new_n570), .A3(new_n663), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n830), .B(new_n834), .C1(new_n671), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT113), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n827), .A2(new_n486), .A3(new_n656), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT50), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n836), .A2(new_n669), .A3(new_n670), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n840), .B(new_n841), .C1(new_n701), .C2(new_n832), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n826), .A2(new_n731), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n749), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n682), .A2(new_n477), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n732), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n842), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n824), .B(new_n838), .C1(KEYINPUT51), .C2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  INV_X1    g666(.A(new_n849), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(KEYINPUT112), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n843), .B1(new_n853), .B2(KEYINPUT112), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n852), .B(new_n842), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n754), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n835), .A2(new_n486), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n656), .A2(new_n732), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n846), .A2(KEYINPUT49), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT49), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n724), .B1(new_n861), .B2(new_n847), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n857), .B1(new_n858), .B2(new_n863), .ZN(G75));
  NOR2_X1   g678(.A1(new_n314), .A2(G952), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n403), .A2(new_n405), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(new_n347), .Z(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT115), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT55), .Z(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(KEYINPUT117), .B2(KEYINPUT56), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n802), .A2(new_n812), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(G902), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n874), .A2(G210), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n871), .B(new_n875), .C1(KEYINPUT117), .C2(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n869), .B1(new_n875), .B2(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT116), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n877), .A2(KEYINPUT116), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n865), .B(new_n876), .C1(new_n878), .C2(new_n879), .ZN(G51));
  INV_X1    g694(.A(new_n763), .ZN(new_n881));
  AOI221_X4 g695(.A(new_n776), .B1(new_n717), .B2(new_n718), .C1(new_n771), .C2(new_n773), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT111), .B1(new_n774), .B2(new_n719), .ZN(new_n883));
  OAI211_X1 g697(.A(KEYINPUT53), .B(new_n881), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n884), .A2(new_n800), .A3(new_n793), .ZN(new_n885));
  AOI211_X1 g699(.A(KEYINPUT109), .B(KEYINPUT53), .C1(new_n818), .C2(new_n789), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n810), .B1(new_n806), .B2(new_n807), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT54), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n814), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n872), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n478), .B(KEYINPUT57), .Z(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT119), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n891), .A2(new_n896), .A3(new_n892), .A4(new_n893), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT120), .B1(new_n898), .B2(new_n680), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  INV_X1    g714(.A(new_n680), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n900), .B(new_n901), .C1(new_n895), .C2(new_n897), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n873), .A2(new_n735), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n865), .B1(new_n903), .B2(new_n904), .ZN(G54));
  NAND3_X1  g719(.A1(new_n874), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(new_n271), .Z(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n865), .ZN(G60));
  NAND2_X1  g722(.A1(new_n600), .A2(new_n601), .ZN(new_n909));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n891), .A2(new_n909), .A3(new_n892), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n824), .A2(new_n911), .ZN(new_n914));
  OAI221_X1 g728(.A(new_n913), .B1(G952), .B2(new_n314), .C1(new_n914), .C2(new_n909), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(G63));
  XNOR2_X1  g730(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n292), .A2(new_n305), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n872), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n865), .B1(new_n921), .B2(new_n630), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n561), .A2(new_n564), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n922), .B(new_n924), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g739(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G66));
  OAI21_X1  g741(.A(G953), .B1(new_n318), .B2(new_n345), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n804), .B2(new_n315), .ZN(new_n929));
  INV_X1    g743(.A(G898), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n866), .B1(new_n930), .B2(new_n315), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n929), .B(new_n931), .Z(G69));
  XNOR2_X1  g746(.A(new_n232), .B(KEYINPUT123), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n513), .B(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n315), .A2(G900), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n741), .A2(new_n714), .A3(new_n780), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT127), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n743), .A2(new_n719), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n787), .A2(new_n674), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT124), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n941), .B(new_n721), .C1(new_n937), .C2(KEYINPUT127), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n939), .A2(new_n751), .A3(new_n942), .ZN(new_n943));
  OAI221_X1 g757(.A(new_n935), .B1(G227), .B2(new_n936), .C1(new_n943), .C2(new_n315), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n671), .B1(new_n311), .B2(new_n669), .ZN(new_n945));
  INV_X1    g759(.A(new_n658), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n714), .A2(new_n945), .A3(new_n731), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n743), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT126), .Z(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n751), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n941), .A2(new_n667), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n951), .A2(new_n953), .ZN(new_n956));
  AND4_X1   g770(.A1(new_n314), .A2(new_n950), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(G227), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n934), .B1(new_n958), .B2(new_n936), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n944), .B1(new_n957), .B2(new_n959), .ZN(G72));
  NAND4_X1  g774(.A1(new_n950), .A2(new_n804), .A3(new_n955), .A4(new_n956), .ZN(new_n961));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT63), .Z(new_n963));
  AOI211_X1 g777(.A(new_n507), .B(new_n514), .C1(new_n961), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n579), .A2(new_n516), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n823), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n943), .A2(new_n804), .ZN(new_n967));
  AOI211_X1 g781(.A(new_n508), .B(new_n515), .C1(new_n967), .C2(new_n963), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n964), .A2(new_n966), .A3(new_n865), .A4(new_n968), .ZN(G57));
endmodule


