//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n204), .ZN(new_n228));
  NOR2_X1   g0028(.A1(G58), .A2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT64), .Z(new_n232));
  AOI211_X1 g0032(.A(new_n209), .B(new_n226), .C1(new_n228), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n223), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n214), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G222), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G223), .A2(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  OAI211_X1 g0059(.A(G1), .B(G13), .C1(new_n251), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n258), .B(new_n261), .C1(G77), .C2(new_n254), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n263), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n262), .B(new_n266), .C1(new_n218), .C2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G179), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n270));
  OAI21_X1  g0070(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n271));
  INV_X1    g0071(.A(G150), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n204), .A2(G33), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n271), .B1(new_n272), .B2(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n227), .ZN(new_n279));
  INV_X1    g0079(.A(G13), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n280), .A2(new_n204), .A3(G1), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n277), .A2(new_n279), .B1(new_n217), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(new_n203), .B2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n268), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n270), .A2(new_n285), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT70), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n268), .A2(G200), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(new_n291), .B2(new_n285), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n294), .B2(KEYINPUT71), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n268), .A2(new_n300), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n297), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n299), .B1(new_n297), .B2(new_n301), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n290), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT16), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n252), .A2(new_n204), .A3(new_n253), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT7), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n253), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n211), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n222), .A2(new_n211), .ZN(new_n311));
  OAI21_X1  g0111(.A(G20), .B1(new_n311), .B2(new_n229), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n273), .A2(G159), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n305), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT74), .ZN(new_n316));
  INV_X1    g0116(.A(new_n279), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n308), .A2(new_n309), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n314), .B1(new_n318), .B2(G68), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n317), .B1(new_n319), .B2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT74), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n321), .B(new_n305), .C1(new_n310), .C2(new_n314), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n316), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n283), .A2(new_n275), .ZN(new_n324));
  INV_X1    g0124(.A(new_n281), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n275), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n218), .A2(G1698), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n329), .B1(G223), .B2(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G87), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n265), .B1(new_n334), .B2(new_n261), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n260), .A2(G232), .A3(new_n263), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G169), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(new_n338), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n328), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT18), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n328), .A2(KEYINPUT18), .A3(new_n341), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n283), .A2(G77), .ZN(new_n348));
  XOR2_X1   g0148(.A(new_n348), .B(KEYINPUT68), .Z(new_n349));
  INV_X1    g0149(.A(new_n275), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n273), .B1(G20), .B2(G77), .ZN(new_n351));
  XOR2_X1   g0151(.A(KEYINPUT15), .B(G87), .Z(new_n352));
  NOR2_X1   g0152(.A1(new_n251), .A2(G20), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n355), .A2(new_n317), .B1(G77), .B2(new_n325), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  INV_X1    g0158(.A(new_n254), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(G238), .B2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n223), .B2(G1698), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n261), .C1(G107), .C2(new_n254), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n266), .B1(new_n267), .B2(new_n220), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT67), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n358), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT69), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n349), .A2(new_n356), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT69), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n362), .A2(new_n364), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(new_n358), .ZN(new_n370));
  INV_X1    g0170(.A(new_n369), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n366), .B(new_n370), .C1(new_n300), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n286), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n340), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n357), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n358), .B1(new_n335), .B2(new_n337), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n260), .B1(new_n332), .B2(new_n333), .ZN(new_n378));
  NOR4_X1   g0178(.A1(new_n378), .A2(new_n300), .A3(new_n336), .A4(new_n265), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n323), .A2(new_n327), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g0183(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n384));
  NAND4_X1  g0184(.A1(new_n323), .A2(new_n327), .A3(new_n380), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n347), .A2(new_n376), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n260), .A2(G238), .A3(new_n263), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n218), .A2(new_n255), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n254), .B(new_n389), .C1(G232), .C2(new_n255), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT72), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(G33), .A3(G97), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n266), .B(new_n388), .C1(new_n396), .C2(new_n260), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT13), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n397), .A2(KEYINPUT13), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G190), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n280), .A2(G1), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n211), .A2(G20), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT12), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(G68), .B2(new_n283), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n405), .B1(new_n276), .B2(new_n219), .C1(new_n274), .C2(new_n217), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n279), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT11), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(G200), .B1(new_n399), .B2(new_n400), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n402), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT14), .B1(new_n401), .B2(new_n286), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n401), .A2(KEYINPUT73), .A3(G179), .ZN(new_n416));
  INV_X1    g0216(.A(new_n400), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(G179), .A3(new_n398), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT73), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT14), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(G169), .C1(new_n399), .C2(new_n400), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n415), .A2(new_n416), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n412), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n414), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n304), .A2(new_n387), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n325), .A2(new_n352), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n325), .B(new_n317), .C1(G1), .C2(new_n251), .ZN(new_n429));
  INV_X1    g0229(.A(new_n352), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n254), .A2(new_n204), .A3(G68), .ZN(new_n433));
  OR2_X1    g0233(.A1(KEYINPUT76), .A2(G97), .ZN(new_n434));
  NAND2_X1  g0234(.A1(KEYINPUT76), .A2(G97), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n353), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT80), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT19), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n436), .B2(new_n438), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n433), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT19), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n204), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT79), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n434), .A2(new_n435), .ZN(new_n445));
  INV_X1    g0245(.A(G87), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n213), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n444), .B1(new_n443), .B2(new_n447), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n441), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n428), .B(new_n432), .C1(new_n450), .C2(new_n317), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n220), .A2(G1698), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n254), .B(new_n453), .C1(G238), .C2(G1698), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G116), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n260), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G250), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n457), .A2(G1), .A3(G274), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n261), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n340), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT78), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT78), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n465), .A3(new_n340), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n456), .A2(new_n461), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n464), .A2(new_n466), .B1(new_n286), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n433), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT76), .A2(G97), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT76), .A2(G97), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n276), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT80), .B1(new_n472), .B2(KEYINPUT19), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n443), .A2(new_n447), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT79), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n427), .B1(new_n479), .B2(new_n279), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n432), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n452), .A2(new_n468), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n279), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n467), .A2(G200), .ZN(new_n485));
  INV_X1    g0285(.A(new_n429), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G87), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n428), .A4(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n467), .A2(new_n300), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n255), .A2(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n254), .A2(G244), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n220), .B1(new_n252), .B2(new_n253), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n493), .B(new_n494), .C1(new_n495), .C2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n254), .A2(G250), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n255), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n261), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT77), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n458), .B(new_n500), .C1(KEYINPUT5), .C2(new_n259), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n203), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT77), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G257), .A3(new_n260), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n501), .A2(new_n503), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(G274), .A3(new_n260), .A4(new_n504), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n499), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G200), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n213), .B1(new_n308), .B2(new_n309), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n434), .A2(KEYINPUT6), .A3(new_n213), .A4(new_n435), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT6), .ZN(new_n514));
  AND2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  NOR2_X1   g0315(.A1(G97), .A2(G107), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n204), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n274), .A2(new_n219), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n317), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n429), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n325), .A2(G97), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n499), .A2(new_n506), .A3(new_n508), .A4(G190), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n510), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n509), .A2(new_n286), .ZN(new_n528));
  INV_X1    g0328(.A(new_n523), .ZN(new_n529));
  INV_X1    g0329(.A(new_n524), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n511), .A2(new_n518), .A3(new_n519), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n317), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n499), .A2(new_n506), .A3(new_n508), .A4(new_n340), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n204), .B(G87), .C1(new_n330), .C2(new_n331), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT22), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n254), .A2(new_n537), .A3(new_n204), .A4(G87), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n213), .A2(G20), .ZN(new_n540));
  XOR2_X1   g0340(.A(new_n540), .B(KEYINPUT23), .Z(new_n541));
  NAND3_X1  g0341(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n539), .A2(KEYINPUT24), .A3(new_n541), .A4(new_n542), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n279), .A3(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(G250), .B(new_n255), .C1(new_n330), .C2(new_n331), .ZN(new_n548));
  OAI211_X1 g0348(.A(G257), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G294), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT85), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT85), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n548), .A2(new_n549), .A3(new_n553), .A4(new_n550), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n261), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n505), .A2(G264), .A3(new_n260), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(G190), .A3(new_n508), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n486), .A2(G107), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n404), .A2(new_n540), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n559), .B(KEYINPUT25), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n547), .A2(new_n557), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n555), .A2(new_n508), .A3(new_n556), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(new_n358), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n527), .B(new_n534), .C1(new_n561), .C2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n491), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n486), .A2(G116), .ZN(new_n566));
  INV_X1    g0366(.A(G116), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n281), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g0368(.A(new_n568), .B(KEYINPUT83), .Z(new_n569));
  AOI21_X1  g0369(.A(G20), .B1(G33), .B2(G283), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n445), .B2(G33), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n278), .A2(new_n227), .B1(G20), .B2(new_n567), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT20), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(KEYINPUT20), .A3(new_n572), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n573), .B1(KEYINPUT84), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT84), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n576), .B(KEYINPUT20), .C1(new_n571), .C2(new_n572), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n566), .B(new_n569), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n505), .A2(G270), .A3(new_n260), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n254), .A2(G257), .A3(new_n255), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n254), .A2(G264), .A3(G1698), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT82), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n359), .A2(G303), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT82), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n254), .A2(new_n584), .A3(G264), .A4(G1698), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n508), .B(new_n579), .C1(new_n586), .C2(new_n260), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n578), .A2(G169), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n547), .A2(new_n558), .A3(new_n560), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n562), .A2(new_n340), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n555), .A2(new_n508), .A3(new_n556), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n286), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n587), .A2(new_n340), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n578), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n578), .A2(KEYINPUT21), .A3(new_n587), .A4(G169), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n590), .A2(new_n595), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n587), .A2(G200), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n587), .A2(new_n300), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n600), .A2(new_n601), .A3(new_n578), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n426), .A2(new_n565), .A3(new_n603), .ZN(G372));
  NOR2_X1   g0404(.A1(new_n414), .A2(new_n375), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n424), .B2(new_n423), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n346), .B1(new_n606), .B2(new_n386), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n302), .A2(new_n303), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n290), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n426), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n488), .A2(new_n489), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n448), .A2(new_n449), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n317), .B1(new_n612), .B2(new_n475), .ZN(new_n613));
  NOR4_X1   g0413(.A1(new_n613), .A2(KEYINPUT81), .A3(new_n427), .A4(new_n431), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n481), .B1(new_n480), .B2(new_n432), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n611), .B1(new_n616), .B2(new_n468), .ZN(new_n617));
  INV_X1    g0417(.A(new_n534), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n617), .A2(KEYINPUT87), .A3(KEYINPUT26), .A4(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT86), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n488), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n489), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n480), .A2(KEYINPUT86), .A3(new_n485), .A4(new_n487), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n451), .B(new_n463), .C1(G169), .C2(new_n462), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n618), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n483), .A2(new_n490), .A3(KEYINPUT26), .A4(new_n618), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT87), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n619), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n564), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(new_n599), .A3(new_n625), .A4(new_n624), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n625), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n609), .B1(new_n610), .B2(new_n637), .ZN(G369));
  NAND3_X1  g0438(.A1(new_n590), .A2(new_n597), .A3(new_n598), .ZN(new_n639));
  OR3_X1    g0439(.A1(new_n404), .A2(KEYINPUT27), .A3(G20), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT27), .B1(new_n404), .B2(G20), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n578), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n639), .A2(new_n645), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n646), .A2(new_n647), .A3(new_n602), .ZN(new_n648));
  INV_X1    g0448(.A(G330), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n561), .A2(new_n563), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n591), .B2(new_n644), .ZN(new_n653));
  INV_X1    g0453(.A(new_n595), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n595), .A2(new_n644), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n644), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(new_n639), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n595), .B2(new_n644), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n659), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n207), .ZN(new_n664));
  OR3_X1    g0464(.A1(new_n664), .A2(KEYINPUT88), .A3(G41), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT88), .B1(new_n664), .B2(G41), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n447), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(G1), .A3(new_n567), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n232), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n667), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT89), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n636), .A2(new_n660), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(KEYINPUT29), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n483), .A2(new_n490), .A3(new_n627), .A4(new_n618), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n644), .B1(new_n678), .B2(new_n635), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n565), .A2(new_n603), .A3(new_n660), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n462), .A2(new_n555), .A3(new_n556), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n499), .A2(new_n506), .A3(new_n508), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n596), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n685), .A2(G179), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n467), .A3(new_n593), .A4(new_n587), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n644), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n695), .A3(new_n644), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n649), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n682), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n673), .B1(new_n701), .B2(G1), .ZN(G364));
  INV_X1    g0502(.A(new_n667), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n280), .A2(G20), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n203), .B1(new_n704), .B2(G45), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n204), .A2(new_n340), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n709), .A2(G190), .A3(G200), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G311), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n359), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n204), .A2(G179), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n300), .A3(new_n358), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n300), .A2(new_n358), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n714), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n716), .A2(G329), .B1(new_n719), .B2(G303), .ZN(new_n720));
  INV_X1    g0520(.A(G294), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n300), .A2(G179), .A3(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n204), .ZN(new_n723));
  INV_X1    g0523(.A(G322), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n709), .A2(new_n300), .A3(G200), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n720), .B1(new_n721), .B2(new_n723), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n709), .A2(new_n358), .A3(G190), .ZN(new_n728));
  XNOR2_X1  g0528(.A(KEYINPUT33), .B(G317), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n713), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G283), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n714), .A2(new_n300), .A3(G200), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT93), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G326), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n708), .A2(new_n717), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n730), .B1(new_n731), .B2(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G159), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT32), .B1(new_n715), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n217), .B2(new_n738), .ZN(new_n742));
  INV_X1    g0542(.A(new_n728), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n743), .A2(new_n211), .B1(new_n522), .B2(new_n723), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n742), .B(new_n744), .C1(G77), .C2(new_n710), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n725), .A2(G58), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n715), .A2(KEYINPUT32), .A3(new_n740), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n718), .A2(new_n446), .ZN(new_n748));
  INV_X1    g0548(.A(new_n736), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n359), .B(new_n748), .C1(new_n749), .C2(G107), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n750), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n739), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(G1), .B(G13), .C1(new_n204), .C2(G169), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT92), .Z(new_n754));
  OAI21_X1  g0554(.A(new_n707), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT90), .Z(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n204), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT91), .Z(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n754), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n664), .A2(new_n359), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G355), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n245), .A2(new_n457), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n664), .A2(new_n254), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n670), .B2(G45), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n764), .B1(G116), .B2(new_n207), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n755), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT94), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n648), .B2(new_n760), .ZN(new_n772));
  INV_X1    g0572(.A(new_n707), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n651), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n649), .B2(new_n648), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(G396));
  NAND2_X1  g0577(.A1(new_n357), .A2(new_n644), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n372), .A2(new_n375), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(KEYINPUT96), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT96), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n372), .A2(new_n781), .A3(new_n375), .A4(new_n778), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n636), .A2(new_n660), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n674), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n782), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n375), .B2(new_n660), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n784), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(new_n699), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n699), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n789), .A2(new_n773), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n723), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G58), .ZN(new_n793));
  INV_X1    g0593(.A(G132), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G143), .A2(new_n725), .B1(new_n710), .B2(G159), .ZN(new_n795));
  INV_X1    g0595(.A(new_n738), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G137), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n795), .B(new_n797), .C1(new_n272), .C2(new_n743), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT34), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n793), .B1(new_n794), .B2(new_n715), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n799), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n749), .A2(G68), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n359), .B1(new_n719), .B2(G50), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n801), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n736), .A2(new_n446), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n711), .A2(new_n567), .B1(new_n712), .B2(new_n715), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n359), .B1(new_n726), .B2(new_n721), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n723), .A2(new_n522), .B1(new_n718), .B2(new_n213), .ZN(new_n809));
  NOR4_X1   g0609(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G303), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n731), .B2(new_n743), .C1(new_n811), .C2(new_n738), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n754), .B1(new_n805), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n754), .B1(G13), .B2(G33), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT95), .Z(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n773), .B(new_n813), .C1(new_n219), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n757), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n787), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n791), .A2(new_n819), .ZN(G384));
  INV_X1    g0620(.A(KEYINPUT40), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n412), .A2(new_n660), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n423), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT98), .ZN(new_n826));
  INV_X1    g0626(.A(new_n822), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n425), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n825), .B1(new_n828), .B2(new_n824), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT103), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n694), .A2(new_n830), .A3(new_n696), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(new_n694), .B2(new_n696), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n787), .B(new_n829), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n320), .A2(new_n315), .B1(new_n324), .B2(new_n326), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT99), .ZN(new_n836));
  INV_X1    g0636(.A(new_n642), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT99), .B1(new_n834), .B2(new_n642), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n347), .B2(new_n386), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n835), .A2(new_n341), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n381), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT37), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT100), .B1(new_n328), .B2(new_n837), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT100), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n846), .B(new_n642), .C1(new_n323), .C2(new_n327), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n342), .B(new_n381), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n844), .B1(new_n848), .B2(KEYINPUT37), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n841), .A2(new_n849), .A3(KEYINPUT38), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n841), .B2(new_n849), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n821), .B1(new_n833), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n697), .A2(KEYINPUT103), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n694), .A2(new_n696), .A3(new_n830), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n848), .B(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n845), .A2(new_n847), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT101), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n383), .A2(new_n862), .A3(new_n385), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n383), .B2(new_n385), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n861), .B1(new_n865), .B2(new_n346), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n858), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n821), .B1(new_n867), .B2(new_n850), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n857), .A2(new_n787), .A3(new_n829), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n854), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n426), .A2(new_n857), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n870), .B(new_n871), .Z(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(G330), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n861), .A2(new_n859), .A3(new_n342), .A4(new_n381), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n848), .A2(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n386), .A2(KEYINPUT101), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n383), .A2(new_n862), .A3(new_n385), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n346), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n861), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n875), .A2(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n874), .B(new_n850), .C1(new_n881), .C2(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT102), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT39), .B1(new_n851), .B2(new_n852), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT102), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n867), .A2(new_n885), .A3(new_n874), .A4(new_n850), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n423), .A2(new_n424), .A3(new_n660), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n347), .A2(new_n642), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n375), .A2(new_n644), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n784), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n893), .B(new_n829), .C1(new_n851), .C2(new_n852), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n889), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n426), .B1(new_n675), .B2(new_n681), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n609), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n895), .B(new_n897), .Z(new_n898));
  XNOR2_X1  g0698(.A(new_n873), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n203), .B2(new_n704), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n670), .A2(new_n219), .A3(new_n311), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n211), .A2(G50), .ZN(new_n902));
  OAI211_X1 g0702(.A(G1), .B(new_n280), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n513), .A2(new_n517), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n567), .B1(new_n904), .B2(KEYINPUT35), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(new_n228), .C1(KEYINPUT35), .C2(new_n904), .ZN(new_n906));
  XOR2_X1   g0706(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n907));
  XNOR2_X1  g0707(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n900), .A2(new_n903), .A3(new_n908), .ZN(G367));
  NOR2_X1   g0709(.A1(new_n743), .A2(new_n740), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n749), .A2(G77), .ZN(new_n911));
  AOI22_X1  g0711(.A1(G50), .A2(new_n710), .B1(new_n725), .B2(G150), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n792), .A2(G68), .B1(new_n796), .B2(G143), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n911), .A2(new_n254), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(KEYINPUT106), .B(G137), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n910), .B(new_n914), .C1(new_n716), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n719), .A2(G58), .ZN(new_n917));
  AOI22_X1  g0717(.A1(G294), .A2(new_n728), .B1(new_n725), .B2(G303), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(new_n359), .C1(new_n731), .C2(new_n711), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n736), .A2(new_n445), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n792), .A2(G107), .B1(new_n796), .B2(G311), .ZN(new_n921));
  INV_X1    g0721(.A(G317), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n715), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n919), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT105), .B1(new_n719), .B2(G116), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT46), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n916), .A2(new_n917), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT47), .Z(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n761), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n480), .A2(new_n487), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n644), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n624), .A2(new_n625), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n625), .B2(new_n931), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(new_n759), .ZN(new_n934));
  INV_X1    g0734(.A(new_n766), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n762), .B1(new_n207), .B2(new_n430), .C1(new_n240), .C2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n929), .A2(new_n707), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n527), .B(new_n534), .C1(new_n525), .C2(new_n660), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n534), .B2(new_n660), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT104), .Z(new_n941));
  NOR2_X1   g0741(.A1(new_n661), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT42), .Z(new_n943));
  INV_X1    g0743(.A(new_n941), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n654), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n644), .B1(new_n945), .B2(new_n534), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n938), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n659), .A2(new_n944), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n947), .A2(new_n949), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n953), .B1(new_n951), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n662), .A2(new_n941), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT44), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n662), .A2(new_n941), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n659), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n639), .A2(new_n660), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n658), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n661), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(new_n650), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n700), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n959), .B(new_n961), .C1(new_n651), .C2(new_n658), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n963), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n701), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n667), .B(KEYINPUT41), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n706), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n937), .B1(new_n957), .B2(new_n975), .ZN(G387));
  NAND2_X1  g0776(.A1(new_n967), .A2(new_n706), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT107), .Z(new_n978));
  NOR2_X1   g0778(.A1(new_n430), .A2(new_n723), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G50), .B2(new_n725), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT108), .Z(new_n981));
  AOI22_X1  g0781(.A1(new_n728), .A2(new_n350), .B1(new_n796), .B2(G159), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n272), .B2(new_n715), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n711), .A2(new_n211), .B1(new_n718), .B2(new_n219), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n983), .A2(new_n359), .A3(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n981), .B(new_n985), .C1(new_n522), .C2(new_n736), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G303), .A2(new_n710), .B1(new_n728), .B2(G311), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n922), .B2(new_n726), .C1(new_n724), .C2(new_n738), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT48), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n731), .B2(new_n723), .C1(new_n721), .C2(new_n718), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT49), .Z(new_n991));
  OAI221_X1 g0791(.A(new_n359), .B1(new_n737), .B2(new_n715), .C1(new_n736), .C2(new_n567), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n986), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n761), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n935), .B1(new_n237), .B2(G45), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n668), .A2(new_n567), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(new_n763), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n350), .A2(new_n217), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT50), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n211), .A2(new_n219), .ZN(new_n1000));
  NOR4_X1   g0800(.A1(new_n999), .A2(G45), .A3(new_n996), .A4(new_n1000), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n997), .A2(new_n1001), .B1(G107), .B2(new_n207), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n773), .B1(new_n1002), .B2(new_n762), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n994), .B(new_n1003), .C1(new_n657), .C2(new_n759), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT109), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n703), .B1(new_n701), .B2(new_n967), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n978), .B(new_n1005), .C1(new_n969), .C2(new_n1006), .ZN(G393));
  INV_X1    g0807(.A(KEYINPUT110), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n963), .A2(new_n1008), .A3(new_n970), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n962), .A2(KEYINPUT110), .A3(new_n659), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT111), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT111), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1009), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n706), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n773), .B1(new_n941), .B2(new_n760), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n762), .B1(new_n207), .B2(new_n445), .C1(new_n248), .C2(new_n935), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n792), .A2(G77), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n743), .B2(new_n217), .C1(new_n275), .C2(new_n711), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT113), .Z(new_n1020));
  AOI22_X1  g0820(.A1(new_n725), .A2(G159), .B1(new_n796), .B2(G150), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT112), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n359), .B1(new_n1022), .B2(KEYINPUT51), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n806), .B1(G68), .B2(new_n719), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(KEYINPUT51), .C2(new_n1022), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1020), .B(new_n1025), .C1(G143), .C2(new_n716), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n725), .A2(G311), .B1(new_n796), .B2(G317), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT52), .Z(new_n1028));
  AOI22_X1  g0828(.A1(new_n749), .A2(G107), .B1(G303), .B2(new_n728), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n731), .C2(new_n718), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n723), .A2(new_n567), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n711), .A2(new_n721), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n359), .B1(new_n715), .B2(new_n724), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n761), .B1(new_n1026), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1016), .A2(new_n1017), .A3(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n971), .B(new_n703), .C1(new_n1011), .C2(new_n969), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1015), .A2(new_n1036), .A3(new_n1037), .ZN(G390));
  NAND2_X1  g0838(.A1(new_n867), .A2(new_n850), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n888), .B(KEYINPUT114), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n891), .B1(new_n679), .B2(new_n783), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n829), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1039), .B(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n698), .A2(new_n787), .A3(new_n829), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n888), .B1(new_n893), .B2(new_n829), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1043), .B(new_n1044), .C1(new_n1045), .C2(new_n887), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n887), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n857), .A2(G330), .A3(new_n787), .A4(new_n829), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1046), .A2(KEYINPUT115), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1047), .A2(KEYINPUT115), .A3(new_n1049), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n706), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n254), .B(new_n748), .C1(G283), .C2(new_n796), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n803), .A2(new_n1018), .A3(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n711), .A2(new_n445), .B1(new_n721), .B2(new_n715), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n213), .B2(new_n743), .C1(new_n567), .C2(new_n726), .ZN(new_n1058));
  INV_X1    g0858(.A(G125), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n715), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(G128), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n254), .B1(new_n1061), .B2(new_n738), .C1(new_n726), .C2(new_n794), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(G159), .C2(new_n792), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT54), .B(G143), .Z(new_n1064));
  AOI22_X1  g0864(.A1(new_n749), .A2(G50), .B1(new_n710), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n915), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1063), .B(new_n1065), .C1(new_n743), .C2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n719), .A2(G150), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT53), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1058), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n773), .B1(new_n1070), .B2(new_n761), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n350), .B2(new_n815), .C1(new_n887), .C2(new_n818), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1053), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n426), .A2(new_n857), .A3(G330), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n896), .A2(new_n1074), .A3(new_n609), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(G330), .B(new_n787), .C1(new_n831), .C2(new_n832), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n1042), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1078), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n787), .A2(G330), .A3(new_n694), .A4(new_n696), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1042), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1048), .A2(new_n1081), .B1(new_n784), .B2(new_n892), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1076), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT117), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1083), .B(new_n1086), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1046), .A2(KEYINPUT115), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1047), .A2(KEYINPUT115), .A3(new_n1049), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1081), .B1(new_n1077), .B2(new_n1042), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n893), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1078), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1075), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(new_n1092), .A3(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1097), .A2(KEYINPUT116), .A3(new_n703), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT116), .B1(new_n1097), .B2(new_n703), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1088), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT118), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1088), .B(KEYINPUT118), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1073), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G378));
  INV_X1    g0905(.A(KEYINPUT57), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1075), .B1(new_n1052), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n854), .A2(G330), .A3(new_n869), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n285), .A2(new_n837), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n304), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n304), .A2(new_n1115), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1111), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1118), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(new_n1110), .A3(new_n1116), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1109), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1124), .A2(new_n854), .A3(G330), .A4(new_n869), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n895), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n895), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1123), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1106), .B1(new_n1108), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1129), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1128), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1097), .A2(new_n1076), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1135), .A3(KEYINPUT57), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n703), .A3(new_n1136), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1132), .A2(new_n1133), .A3(new_n705), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1124), .A2(new_n757), .ZN(new_n1139));
  INV_X1    g0939(.A(G124), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n251), .B1(new_n715), .B2(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n723), .A2(new_n272), .B1(new_n738), .B2(new_n1059), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1064), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n726), .A2(new_n1061), .B1(new_n718), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(G137), .C2(new_n710), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n794), .B2(new_n743), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G41), .B(new_n1141), .C1(new_n1146), .C2(KEYINPUT59), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(KEYINPUT59), .B2(new_n1146), .C1(new_n740), .C2(new_n736), .ZN(new_n1148));
  AOI21_X1  g0948(.A(G41), .B1(new_n710), .B2(new_n352), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n731), .B2(new_n715), .C1(new_n522), .C2(new_n743), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G107), .B2(new_n725), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n254), .B1(new_n749), .B2(G58), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n792), .A2(G68), .B1(new_n719), .B2(G77), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n796), .A2(G116), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT58), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G50), .B1(new_n253), .B2(new_n259), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT119), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1148), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n761), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n773), .B1(new_n816), .B2(new_n217), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1139), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1138), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1137), .A2(new_n1164), .ZN(G375));
  NAND3_X1  g0965(.A1(new_n1094), .A2(new_n1075), .A3(new_n1095), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1083), .A2(new_n974), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n715), .A2(new_n811), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n911), .A2(new_n359), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT122), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n711), .A2(new_n213), .B1(new_n718), .B2(new_n522), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n979), .B(new_n1171), .C1(G116), .C2(new_n728), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n721), .C2(new_n738), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1168), .B(new_n1173), .C1(G283), .C2(new_n725), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n749), .A2(G58), .B1(G150), .B2(new_n710), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n794), .B2(new_n738), .C1(new_n740), .C2(new_n718), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n726), .A2(new_n1066), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n743), .A2(new_n1143), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n254), .B1(new_n715), .B2(new_n1061), .C1(new_n723), .C2(new_n217), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n761), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n707), .C1(G68), .C2(new_n815), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1042), .B2(new_n756), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1107), .B2(new_n706), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1167), .A2(new_n1184), .ZN(G381));
  INV_X1    g0985(.A(G375), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1073), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1100), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1189), .A2(G384), .A3(G381), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(G390), .A2(G387), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(G393), .A2(G396), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(G407));
  OAI211_X1 g0993(.A(G407), .B(G213), .C1(G343), .C2(new_n1189), .ZN(G409));
  OR2_X1    g0994(.A1(G390), .A2(G387), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(G393), .B(new_n776), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(G390), .A2(G387), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AND2_X1   g0999(.A1(G390), .A2(G387), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1196), .B1(new_n1200), .B2(new_n1191), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n643), .A2(G213), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT60), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n667), .B1(new_n1166), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1094), .A2(new_n1095), .A3(new_n1075), .A4(KEYINPUT60), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1083), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G384), .B1(new_n1207), .B2(new_n1184), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT125), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1207), .A2(G384), .A3(new_n1184), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT124), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G375), .B1(new_n1214), .B2(new_n1187), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT123), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1138), .B2(new_n1163), .ZN(new_n1217));
  OAI211_X1 g1017(.A(KEYINPUT123), .B(new_n1162), .C1(new_n1130), .C2(new_n705), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1134), .A2(new_n1135), .A3(new_n974), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1188), .A2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1203), .B(new_n1213), .C1(new_n1215), .C2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT126), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1188), .A2(new_n1220), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1104), .B2(G375), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1226), .A2(KEYINPUT126), .A3(new_n1203), .A4(new_n1213), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT62), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1203), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n643), .A2(G213), .A3(G2897), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1210), .A2(new_n1212), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT61), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1222), .A2(KEYINPUT62), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1202), .B1(new_n1228), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT63), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1224), .A2(new_n1238), .A3(new_n1227), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1222), .A2(new_n1238), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1234), .A4(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1237), .A2(new_n1242), .ZN(G405));
  INV_X1    g1043(.A(new_n1215), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G375), .A2(new_n1188), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1202), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1213), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1249), .B(new_n1250), .ZN(G402));
endmodule


