//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(KEYINPUT64), .B(G68), .Z(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G58), .A2(G232), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n206), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n206), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NOR4_X1   g0026(.A1(new_n218), .A2(new_n219), .A3(new_n223), .A4(new_n226), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT66), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n222), .ZN(new_n246));
  INV_X1    g0046(.A(G107), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT7), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G20), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT74), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT74), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  AOI21_X1  g0053(.A(G33), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n250), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n249), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n259), .A2(new_n255), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n248), .B1(new_n260), .B2(G20), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n247), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT6), .ZN(new_n263));
  INV_X1    g0063(.A(G97), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n263), .A2(new_n264), .A3(G107), .ZN(new_n265));
  XNOR2_X1  g0065(.A(G97), .B(G107), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G77), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n267), .A2(new_n221), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n246), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(KEYINPUT68), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT68), .A2(G1), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n273), .A2(G13), .A3(G20), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n264), .ZN(new_n277));
  INV_X1    g0077(.A(new_n246), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n273), .A2(G33), .A3(new_n274), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n280), .B2(new_n264), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n272), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT68), .A2(G1), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT68), .A2(G1), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  OAI211_X1 g0088(.A(G1), .B(G13), .C1(new_n258), .C2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT5), .B(G41), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n287), .A2(G274), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n273), .A2(G45), .A3(new_n274), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT5), .A2(G41), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT5), .A2(G41), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(G257), .B(new_n289), .C1(new_n292), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(KEYINPUT70), .A2(G179), .ZN(new_n299));
  NOR2_X1   g0099(.A1(KEYINPUT70), .A2(G179), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(KEYINPUT4), .A2(G244), .ZN(new_n302));
  INV_X1    g0102(.A(G1698), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n259), .A2(new_n255), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n259), .A2(new_n255), .A3(G250), .A4(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G283), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n259), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(G33), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(G244), .A3(new_n303), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT4), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n307), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n298), .B(new_n301), .C1(new_n313), .C2(new_n289), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n251), .A2(new_n253), .A3(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n259), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n303), .A2(G244), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n289), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n315), .B1(new_n321), .B2(new_n297), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n283), .A2(new_n314), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n264), .A2(new_n247), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G97), .A2(G107), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n263), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n265), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(G20), .B1(G77), .B2(new_n269), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n259), .A2(new_n255), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT7), .B1(new_n330), .B2(new_n221), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n255), .B1(new_n309), .B2(G33), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n249), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n329), .B1(new_n333), .B2(new_n247), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n281), .B1(new_n334), .B2(new_n246), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n336), .B(G200), .C1(new_n321), .C2(new_n297), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n298), .B(G190), .C1(new_n313), .C2(new_n289), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n298), .B1(new_n313), .B2(new_n289), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n336), .B1(new_n340), .B2(G200), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n323), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT21), .ZN(new_n344));
  MUX2_X1   g0144(.A(G257), .B(G264), .S(G1698), .Z(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(new_n316), .A3(new_n259), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT80), .B(G303), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n330), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n289), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(G270), .B(new_n289), .C1(new_n292), .C2(new_n295), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n291), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(G169), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n275), .A2(new_n278), .A3(new_n279), .A4(G116), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G116), .B2(new_n275), .ZN(new_n354));
  INV_X1    g0154(.A(G116), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n245), .A2(new_n222), .B1(G20), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n306), .B(new_n221), .C1(G33), .C2(new_n264), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n356), .A2(KEYINPUT20), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT20), .B1(new_n356), .B2(new_n357), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n344), .B1(new_n352), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n349), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n291), .A2(new_n350), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n353), .B1(G116), .B2(new_n275), .C1(new_n358), .C2(new_n359), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n365), .A2(KEYINPUT21), .A3(G169), .A4(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(G179), .A3(new_n363), .A4(new_n364), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n362), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n363), .B2(new_n364), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(new_n366), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT81), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT81), .B1(new_n373), .B2(new_n366), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n369), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n258), .A2(G20), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT19), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(G97), .ZN(new_n381));
  INV_X1    g0181(.A(G87), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n325), .A2(new_n382), .B1(new_n383), .B2(new_n221), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n384), .B2(new_n380), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n316), .A2(new_n221), .A3(G68), .A4(new_n259), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT77), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n278), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT77), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT76), .ZN(new_n392));
  INV_X1    g0192(.A(G250), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n292), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n284), .A2(new_n285), .ZN(new_n395));
  AOI21_X1  g0195(.A(G274), .B1(new_n392), .B2(G250), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(G45), .A3(new_n396), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n394), .A2(new_n289), .A3(new_n397), .ZN(new_n398));
  MUX2_X1   g0198(.A(G238), .B(G244), .S(G1698), .Z(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(new_n316), .A3(new_n259), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G116), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n289), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(G200), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n280), .A2(new_n382), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT15), .B(G87), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n276), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n391), .A2(new_n403), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n394), .A2(new_n289), .A3(new_n397), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n310), .A2(new_n399), .B1(G33), .B2(G116), .ZN(new_n410));
  OAI211_X1 g0210(.A(G190), .B(new_n409), .C1(new_n410), .C2(new_n289), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n400), .A2(new_n401), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT79), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(G190), .A4(new_n409), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g0218(.A(new_n405), .B(KEYINPUT78), .Z(new_n419));
  OR2_X1    g0219(.A1(new_n419), .A2(new_n280), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n391), .A2(new_n406), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n315), .B1(new_n398), .B2(new_n402), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n415), .A2(new_n301), .A3(new_n409), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n408), .A2(new_n418), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n343), .A2(new_n378), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(KEYINPUT8), .A2(G58), .ZN(new_n427));
  INV_X1    g0227(.A(G58), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT69), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT69), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G58), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n427), .B1(new_n432), .B2(KEYINPUT8), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n379), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n269), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n278), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n246), .B1(new_n395), .B2(G20), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G50), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(G50), .B2(new_n275), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n260), .A2(G222), .A3(new_n303), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n260), .A2(G1698), .ZN(new_n442));
  INV_X1    g0242(.A(G223), .ZN(new_n443));
  OAI221_X1 g0243(.A(new_n441), .B1(new_n268), .B2(new_n260), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n414), .ZN(new_n445));
  NOR2_X1   g0245(.A1(G41), .A2(G45), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n289), .A2(new_n447), .A3(G274), .ZN(new_n448));
  INV_X1    g0248(.A(new_n446), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n414), .B1(new_n395), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n450), .B2(G226), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n440), .B1(new_n452), .B2(new_n315), .ZN(new_n453));
  INV_X1    g0253(.A(new_n301), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(new_n452), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n452), .A2(G200), .B1(new_n440), .B2(KEYINPUT9), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n445), .A2(G190), .A3(new_n451), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n457), .B(new_n458), .C1(KEYINPUT9), .C2(new_n440), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(KEYINPUT10), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(KEYINPUT10), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT69), .B(G58), .ZN(new_n463));
  OAI22_X1  g0263(.A1(new_n207), .A2(new_n463), .B1(G58), .B2(G68), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(G20), .B1(G159), .B2(new_n269), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n317), .A2(new_n248), .A3(new_n221), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G68), .ZN(new_n467));
  AOI21_X1  g0267(.A(G20), .B1(new_n316), .B2(new_n259), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n248), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n465), .B(KEYINPUT16), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT16), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n207), .B1(new_n257), .B2(new_n261), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT64), .B(G68), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n201), .B1(new_n432), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G159), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n474), .A2(new_n221), .B1(new_n475), .B2(new_n270), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n471), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n477), .A3(new_n246), .ZN(new_n478));
  INV_X1    g0278(.A(new_n433), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n479), .A2(new_n437), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n275), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  MUX2_X1   g0283(.A(G223), .B(G226), .S(G1698), .Z(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n316), .A3(new_n259), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G87), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n289), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n289), .A2(new_n447), .A3(G274), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n273), .A2(new_n274), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n289), .B1(new_n489), .B2(new_n446), .ZN(new_n490));
  INV_X1    g0290(.A(G232), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n487), .A2(new_n492), .A3(new_n301), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n487), .A2(new_n492), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(G169), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n483), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT18), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n372), .B1(new_n487), .B2(new_n492), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n494), .B2(G190), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n478), .A2(new_n500), .A3(new_n482), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT17), .ZN(new_n502));
  OR2_X1    g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT18), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n483), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(new_n502), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n498), .A2(new_n503), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n473), .A2(new_n221), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n221), .A2(G33), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n270), .A2(new_n202), .B1(new_n510), .B2(new_n268), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n246), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n512), .B(KEYINPUT11), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT12), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n275), .B2(G68), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n437), .A2(G68), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n276), .A2(KEYINPUT12), .A3(new_n207), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n513), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n259), .A2(new_n255), .A3(G232), .A4(G1698), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n259), .A2(new_n255), .A3(G226), .A4(new_n303), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n383), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n522), .A2(new_n414), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n488), .B1(new_n490), .B2(new_n208), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT13), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n448), .B1(new_n450), .B2(G238), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT13), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n414), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n519), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT14), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n525), .A2(G179), .A3(new_n529), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n518), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n525), .A2(new_n529), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n518), .B1(new_n537), .B2(G190), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(G200), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n442), .A2(new_n208), .B1(new_n247), .B2(new_n260), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n330), .A2(new_n491), .A3(G1698), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n414), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n448), .B1(new_n450), .B2(G244), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n405), .A2(new_n510), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(G20), .B2(G77), .ZN(new_n548));
  XOR2_X1   g0348(.A(KEYINPUT8), .B(G58), .Z(new_n549));
  OR2_X1    g0349(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n278), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT72), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n437), .A2(G77), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G77), .B2(new_n275), .ZN(new_n556));
  OR3_X1    g0356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n543), .A2(G190), .A3(new_n544), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n554), .B1(new_n553), .B2(new_n556), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n546), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n545), .A2(new_n315), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n553), .A2(new_n556), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n543), .A2(new_n301), .A3(new_n544), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n540), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n462), .A2(new_n508), .A3(new_n535), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT85), .ZN(new_n567));
  MUX2_X1   g0367(.A(G250), .B(G257), .S(G1698), .Z(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n316), .A3(new_n259), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G294), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n289), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G264), .B(new_n289), .C1(new_n292), .C2(new_n295), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n315), .B1(new_n574), .B2(new_n291), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n289), .A2(G274), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n576), .A2(new_n292), .A3(new_n295), .ZN(new_n577));
  INV_X1    g0377(.A(G179), .ZN(new_n578));
  NOR4_X1   g0378(.A1(new_n571), .A2(new_n573), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n567), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n571), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n581), .A2(G179), .A3(new_n291), .A4(new_n572), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n571), .A2(new_n573), .A3(new_n577), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(KEYINPUT85), .C1(new_n583), .C2(new_n315), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n316), .A2(new_n221), .A3(G87), .A4(new_n259), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n585), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT82), .B1(new_n585), .B2(KEYINPUT22), .ZN(new_n587));
  NOR4_X1   g0387(.A1(new_n330), .A2(KEYINPUT22), .A3(G20), .A4(new_n382), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT23), .B1(new_n221), .B2(G107), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n594));
  OR3_X1    g0394(.A1(new_n221), .A2(KEYINPUT23), .A3(G107), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT24), .B1(new_n589), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n585), .A2(KEYINPUT22), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT82), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n588), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n585), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  INV_X1    g0403(.A(new_n596), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n278), .B1(new_n597), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n280), .A2(new_n247), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n276), .A2(new_n247), .ZN(new_n608));
  XOR2_X1   g0408(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n609));
  OR2_X1    g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n580), .B(new_n584), .C1(new_n606), .C2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT86), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n603), .B1(new_n602), .B2(new_n604), .ZN(new_n616));
  AOI211_X1 g0416(.A(KEYINPUT24), .B(new_n596), .C1(new_n600), .C2(new_n601), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n246), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n569), .A2(new_n570), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n291), .B(new_n572), .C1(new_n619), .C2(new_n289), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n372), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n583), .A2(new_n370), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n618), .A2(new_n612), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n614), .A2(new_n615), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n580), .A2(new_n584), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n618), .B2(new_n612), .ZN(new_n627));
  INV_X1    g0427(.A(new_n623), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n606), .A2(new_n613), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT86), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n426), .B(new_n566), .C1(new_n625), .C2(new_n630), .ZN(G372));
  INV_X1    g0431(.A(new_n566), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n421), .A2(new_n424), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n421), .A2(new_n424), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n407), .A2(KEYINPUT87), .B1(new_n417), .B2(new_n412), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n389), .A2(new_n390), .B1(new_n276), .B2(new_n405), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n403), .A4(new_n404), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n634), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(new_n343), .A3(new_n624), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n618), .A2(new_n612), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n582), .B1(new_n583), .B2(new_n315), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n369), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n633), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n418), .A2(new_n403), .A3(new_n404), .A4(new_n636), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n283), .A2(new_n314), .A3(new_n322), .ZN(new_n646));
  AND4_X1   g0446(.A1(KEYINPUT26), .A2(new_n645), .A3(new_n633), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n635), .A2(new_n638), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n633), .A3(new_n646), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n632), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n505), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n504), .B1(new_n483), .B2(new_n496), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n535), .ZN(new_n657));
  INV_X1    g0457(.A(new_n564), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n540), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n501), .B(KEYINPUT17), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n656), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n459), .B(KEYINPUT10), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n456), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n653), .A2(new_n664), .ZN(G369));
  AND2_X1   g0465(.A1(new_n221), .A2(G13), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OR3_X1    g0467(.A1(new_n667), .A2(new_n489), .A3(KEYINPUT27), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT27), .B1(new_n489), .B2(new_n667), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n614), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n630), .A2(new_n625), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n641), .A2(new_n672), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n672), .A2(new_n366), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n378), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n369), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  XOR2_X1   g0481(.A(KEYINPUT88), .B(G330), .Z(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n369), .A2(new_n673), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n630), .B2(new_n625), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n641), .A2(new_n642), .A3(new_n673), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n686), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n224), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n325), .A2(new_n382), .A3(new_n355), .ZN(new_n695));
  INV_X1    g0495(.A(G1), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n220), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n694), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  INV_X1    g0500(.A(KEYINPUT89), .ZN(new_n701));
  INV_X1    g0501(.A(new_n626), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n369), .B1(new_n641), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n640), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n614), .A2(new_n680), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n597), .A2(new_n605), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n613), .B1(new_n706), .B2(new_n246), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n342), .B1(new_n707), .B2(new_n623), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n705), .A2(new_n708), .A3(KEYINPUT89), .A4(new_n639), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n645), .A2(new_n646), .A3(new_n650), .A4(new_n633), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n633), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(KEYINPUT26), .B2(new_n649), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n704), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n673), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n715));
  AND4_X1   g0515(.A1(new_n425), .A2(new_n343), .A3(new_n378), .A4(new_n673), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n614), .A2(new_n615), .A3(new_n624), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n615), .B1(new_n614), .B2(new_n624), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n321), .A2(new_n297), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n398), .A2(new_n402), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n574), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n363), .A2(new_n364), .A3(G179), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n722), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n454), .B1(new_n363), .B2(new_n364), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n340), .A2(new_n726), .A3(new_n727), .A4(new_n620), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n722), .A2(new_n574), .ZN(new_n729));
  INV_X1    g0529(.A(new_n724), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n729), .A2(new_n730), .A3(KEYINPUT30), .A4(new_n721), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n672), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n719), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n683), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n740), .B(new_n673), .C1(new_n644), .C2(new_n651), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n715), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n700), .B1(new_n743), .B2(G1), .ZN(G364));
  INV_X1    g0544(.A(new_n684), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n696), .B1(new_n666), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n694), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(new_n683), .B2(new_n681), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n222), .B1(G20), .B2(new_n315), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n240), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n310), .A2(new_n693), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n286), .B2(new_n698), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n757), .A2(G45), .B1(KEYINPUT91), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(KEYINPUT91), .B2(new_n760), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n330), .B(new_n693), .C1(KEYINPUT90), .C2(G355), .ZN(new_n763));
  OR2_X1    g0563(.A1(G355), .A2(KEYINPUT90), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n763), .A2(new_n764), .B1(new_n355), .B2(new_n693), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n756), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n754), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n221), .A2(G179), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n260), .B1(new_n769), .B2(new_n382), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n221), .A2(new_n372), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n454), .A2(G190), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n454), .A2(new_n370), .A3(new_n771), .ZN(new_n773));
  INV_X1    g0573(.A(G68), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n202), .A2(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n221), .A2(new_n370), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n454), .A2(new_n372), .A3(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n770), .B(new_n775), .C1(new_n432), .C2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n454), .A2(G20), .A3(new_n370), .A4(new_n372), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT92), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G77), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n768), .A2(new_n370), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n221), .B1(new_n789), .B2(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n788), .A2(G107), .B1(new_n791), .B2(G97), .ZN(new_n792));
  NOR4_X1   g0592(.A1(new_n221), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G159), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT32), .Z(new_n795));
  NAND4_X1  g0595(.A1(new_n779), .A2(new_n786), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT33), .B(G317), .Z(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n777), .B1(new_n773), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n772), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(G326), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n260), .B1(G329), .B2(new_n793), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(new_n787), .ZN(new_n804));
  INV_X1    g0604(.A(G303), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n769), .A2(new_n805), .B1(new_n790), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n801), .B(new_n808), .C1(new_n784), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n767), .B1(new_n796), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n748), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n766), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n753), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n681), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n750), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n562), .A2(new_n672), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n560), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n564), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n658), .A2(new_n673), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n673), .B(new_n823), .C1(new_n644), .C2(new_n651), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n652), .A2(new_n673), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n822), .B(KEYINPUT95), .Z(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(new_n739), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n748), .B1(new_n827), .B2(new_n739), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n767), .A2(new_n752), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n748), .B1(G77), .B2(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n803), .A2(new_n773), .B1(new_n772), .B2(new_n805), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G294), .B2(new_n778), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n382), .A2(new_n787), .B1(new_n769), .B2(new_n247), .ZN(new_n835));
  INV_X1    g0635(.A(new_n793), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n330), .B1(new_n836), .B2(new_n809), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n835), .B(new_n837), .C1(G97), .C2(new_n791), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n834), .B(new_n838), .C1(new_n355), .C2(new_n784), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G150), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n840), .A2(new_n772), .B1(new_n773), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT93), .ZN(new_n843));
  INV_X1    g0643(.A(G143), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n844), .B2(new_n777), .C1(new_n475), .C2(new_n784), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT34), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n787), .A2(new_n774), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n432), .B2(new_n791), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n202), .B2(new_n769), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n317), .B(new_n850), .C1(G132), .C2(new_n793), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n845), .B2(new_n846), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n839), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n832), .B1(new_n853), .B2(new_n754), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n752), .B2(new_n823), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT94), .Z(new_n856));
  NOR2_X1   g0656(.A1(new_n830), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR3_X1   g0658(.A1(new_n222), .A2(new_n221), .A3(new_n355), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n267), .B(KEYINPUT96), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT35), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT36), .ZN(new_n865));
  OAI211_X1 g0665(.A(G77), .B(new_n698), .C1(new_n207), .C2(new_n463), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n202), .A2(G68), .ZN(new_n867));
  AOI211_X1 g0667(.A(G13), .B(new_n395), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n670), .B(KEYINPUT98), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n656), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n824), .A2(new_n821), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT97), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n535), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT97), .B(new_n518), .C1(new_n532), .C2(new_n534), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n518), .A2(new_n672), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n538), .B2(new_n539), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n532), .A2(new_n534), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n540), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n876), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n872), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n482), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT7), .B1(new_n310), .B2(G20), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n774), .B1(new_n468), .B2(new_n248), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n476), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n278), .B1(new_n888), .B2(KEYINPUT16), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n471), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n885), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n501), .B1(new_n892), .B2(new_n670), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n495), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n483), .A2(new_n870), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n497), .A2(new_n896), .A3(new_n897), .A4(new_n501), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT99), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT99), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n895), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n892), .A2(new_n670), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n507), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n900), .A2(KEYINPUT38), .A3(new_n902), .A4(new_n904), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n871), .B1(new_n884), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n874), .A2(new_n875), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(new_n672), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n497), .A2(new_n896), .A3(new_n501), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(new_n897), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n896), .B1(new_n656), .B2(new_n660), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n906), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT100), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n908), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(new_n907), .B2(new_n908), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n908), .A2(new_n917), .A3(new_n919), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT100), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n913), .B(new_n920), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n910), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n740), .B1(new_n713), .B2(new_n673), .ZN(new_n926));
  INV_X1    g0726(.A(new_n741), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n632), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n664), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n925), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n735), .A2(new_n736), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n675), .B2(new_n716), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n882), .A2(new_n823), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n908), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n899), .A2(KEYINPUT99), .B1(new_n507), .B2(new_n903), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n936), .B2(new_n902), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT40), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n908), .A2(new_n917), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n941), .A3(KEYINPUT40), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n632), .A2(new_n738), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n682), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n944), .B2(new_n943), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n930), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n395), .B2(new_n666), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n930), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n869), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT101), .Z(G367));
  NAND2_X1  g0751(.A1(new_n283), .A2(new_n672), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n323), .B(new_n952), .C1(new_n339), .C2(new_n341), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n646), .A2(new_n672), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n688), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n953), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n646), .B1(new_n627), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT102), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n672), .B1(new_n958), .B2(KEYINPUT102), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n956), .A2(KEYINPUT42), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT103), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n956), .B2(KEYINPUT42), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n956), .A2(new_n962), .A3(KEYINPUT42), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n636), .A2(new_n404), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n672), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n633), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n639), .B2(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT43), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n685), .A2(new_n955), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n956), .A2(new_n962), .A3(KEYINPUT42), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n963), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n978), .A2(new_n971), .A3(new_n970), .A4(new_n961), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n974), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n976), .B1(new_n974), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n694), .B(KEYINPUT41), .Z(new_n983));
  OAI21_X1  g0783(.A(new_n676), .B1(new_n717), .B2(new_n718), .ZN(new_n984));
  INV_X1    g0784(.A(new_n674), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n985), .A3(new_n687), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT105), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n688), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AOI211_X1 g0789(.A(KEYINPUT105), .B(new_n687), .C1(new_n630), .C2(new_n625), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n684), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n745), .B(new_n990), .C1(new_n986), .C2(new_n988), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n742), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT44), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n691), .B2(new_n955), .ZN(new_n996));
  INV_X1    g0796(.A(new_n955), .ZN(new_n997));
  OAI211_X1 g0797(.A(KEYINPUT44), .B(new_n997), .C1(new_n688), .C2(new_n690), .ZN(new_n998));
  INV_X1    g0798(.A(new_n687), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n717), .B2(new_n718), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(new_n689), .A3(new_n955), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1000), .A2(KEYINPUT45), .A3(new_n689), .A4(new_n955), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n996), .A2(new_n998), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n686), .B1(new_n1005), .B2(KEYINPUT104), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1000), .A2(new_n689), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT44), .B1(new_n1007), .B2(new_n997), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n998), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT45), .B1(new_n691), .B2(new_n955), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1004), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1008), .A2(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT104), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n1013), .A3(new_n685), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n994), .A2(new_n1006), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n983), .B1(new_n1015), .B2(new_n743), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n982), .B1(new_n1016), .B2(new_n747), .ZN(new_n1017));
  XOR2_X1   g0817(.A(KEYINPUT106), .B(G311), .Z(new_n1018));
  NOR2_X1   g0818(.A1(new_n769), .A2(new_n355), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n800), .A2(new_n1018), .B1(new_n1019), .B2(KEYINPUT46), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n806), .B2(new_n773), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n787), .A2(new_n264), .B1(new_n790), .B2(new_n247), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n310), .B(new_n1022), .C1(G317), .C2(new_n793), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n347), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1023), .B1(KEYINPUT46), .B2(new_n1019), .C1(new_n1024), .C2(new_n777), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1021), .B(new_n1025), .C1(G283), .C2(new_n785), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n785), .A2(G50), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G143), .A2(new_n800), .B1(new_n778), .B2(G150), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n475), .B2(new_n773), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n260), .B1(new_n769), .B2(new_n463), .C1(new_n836), .C2(new_n840), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n787), .A2(new_n268), .B1(new_n790), .B2(new_n774), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1026), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT47), .Z(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n754), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n970), .A2(new_n753), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n755), .B1(new_n224), .B2(new_n405), .C1(new_n759), .C2(new_n235), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n748), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1017), .A2(new_n1038), .ZN(G387));
  NOR2_X1   g0839(.A1(new_n992), .A2(new_n993), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT108), .B1(new_n1040), .B2(new_n743), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n994), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT108), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n742), .C1(new_n992), .C2(new_n993), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n694), .A4(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n260), .A2(new_n695), .A3(new_n224), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n232), .A2(new_n286), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n549), .A2(new_n202), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n695), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n286), .C1(new_n774), .C2(new_n268), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n758), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1046), .B1(G107), .B2(new_n224), .C1(new_n1047), .C2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n812), .B1(new_n1053), .B2(new_n755), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n268), .A2(new_n769), .B1(new_n787), .B2(new_n264), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n317), .B(new_n1055), .C1(G150), .C2(new_n793), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT107), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n419), .A2(new_n790), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G50), .B2(new_n778), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n475), .B2(new_n772), .C1(new_n479), .C2(new_n773), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1057), .B(new_n1060), .C1(G68), .C2(new_n785), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n773), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G322), .A2(new_n800), .B1(new_n1062), .B2(new_n1018), .ZN(new_n1063));
  INV_X1    g0863(.A(G317), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n777), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n785), .B2(new_n347), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT48), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT48), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n769), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1069), .A2(G294), .B1(new_n791), .B2(G283), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n310), .B1(G326), .B2(new_n793), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n355), .B2(new_n787), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1061), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1054), .B1(new_n1078), .B2(new_n767), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n677), .B2(new_n753), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n1040), .B2(new_n747), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1045), .A2(new_n1081), .ZN(G393));
  AND2_X1   g0882(.A1(new_n243), .A2(new_n758), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n755), .B1(new_n264), .B2(new_n224), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n260), .B1(G322), .B2(new_n793), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n247), .B2(new_n787), .C1(new_n803), .C2(new_n769), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n773), .A2(new_n1024), .B1(new_n355), .B2(new_n790), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(KEYINPUT110), .B2(new_n1087), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(KEYINPUT110), .B2(new_n1087), .C1(new_n806), .C2(new_n784), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n809), .A2(new_n777), .B1(new_n772), .B2(new_n1064), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT52), .Z(new_n1091));
  NOR2_X1   g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT111), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n785), .A2(new_n549), .B1(G50), .B2(new_n1062), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1094), .A2(KEYINPUT109), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(KEYINPUT109), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n841), .A2(new_n772), .B1(new_n777), .B2(new_n475), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT51), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n787), .A2(new_n382), .B1(new_n790), .B2(new_n268), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n310), .B1(new_n844), .B2(new_n836), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n473), .C2(new_n1069), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1093), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT112), .Z(new_n1104));
  OAI221_X1 g0904(.A(new_n748), .B1(new_n1083), .B2(new_n1084), .C1(new_n1104), .C2(new_n767), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n753), .B2(new_n997), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1005), .B(new_n685), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n747), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1015), .B(new_n694), .C1(new_n1107), .C2(new_n994), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(G390));
  INV_X1    g0910(.A(new_n694), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n941), .A2(new_n912), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n713), .A2(new_n673), .A3(new_n820), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n821), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1112), .B1(new_n882), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n343), .A2(new_n378), .A3(new_n425), .A4(new_n673), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n630), .B2(new_n625), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n683), .B(new_n823), .C1(new_n1118), .C2(new_n931), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n883), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n920), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n922), .A2(KEYINPUT100), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n909), .A2(KEYINPUT39), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n912), .B1(new_n872), .B2(new_n883), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1116), .B(new_n1121), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n920), .B1(new_n921), .B2(new_n923), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1115), .B1(new_n1129), .B2(new_n1126), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n822), .B1(new_n878), .B2(new_n881), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n738), .A2(G330), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1128), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(G330), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n719), .B2(new_n737), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT114), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n826), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(G330), .C1(new_n1118), .C2(new_n931), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n883), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1113), .B(new_n821), .C1(new_n1119), .C2(new_n883), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1119), .A2(new_n883), .ZN(new_n1144));
  AOI221_X4 g0944(.A(KEYINPUT113), .B1(new_n821), .B2(new_n824), .C1(new_n1144), .C2(new_n1132), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT113), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1132), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n824), .A2(new_n821), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1143), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1135), .A2(new_n632), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n928), .A2(new_n664), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1111), .B1(new_n1133), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT113), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1147), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1152), .B1(new_n1159), .B2(new_n1143), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n1128), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1155), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1129), .A2(new_n751), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n748), .B1(new_n433), .B2(new_n831), .ZN(new_n1164));
  INV_X1    g0964(.A(G125), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n260), .B1(new_n475), .B2(new_n790), .C1(new_n836), .C2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n769), .A2(new_n841), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1166), .B(new_n1169), .C1(G50), .C2(new_n788), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1171), .A2(new_n772), .B1(new_n773), .B2(new_n840), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G132), .B2(new_n778), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT54), .B(G143), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1170), .B(new_n1173), .C1(new_n784), .C2(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n330), .B1(new_n769), .B2(new_n382), .C1(new_n836), .C2(new_n806), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n848), .B(new_n1176), .C1(G77), .C2(new_n791), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n247), .A2(new_n773), .B1(new_n777), .B2(new_n355), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G283), .B2(new_n800), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(new_n264), .C2(new_n784), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1164), .B1(new_n1181), .B2(new_n754), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1163), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1133), .B2(new_n746), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1162), .A2(new_n1185), .ZN(G378));
  AOI211_X1 g0986(.A(new_n1120), .B(new_n1115), .C1(new_n1129), .C2(new_n1126), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1129), .A2(new_n1126), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1132), .B1(new_n1188), .B2(new_n1116), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1152), .B1(new_n1190), .B2(new_n1150), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1131), .B1(new_n1118), .B2(new_n931), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n907), .B2(new_n908), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n942), .B(G330), .C1(new_n1193), .C2(KEYINPUT40), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n462), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n440), .A2(new_n670), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n462), .B1(new_n440), .B2(new_n670), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1194), .A2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n940), .A2(G330), .A3(new_n942), .A4(new_n1204), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n925), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n924), .A4(new_n910), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(KEYINPUT57), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n694), .B1(new_n1191), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1153), .B1(new_n1133), .B2(new_n1154), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1214), .B2(new_n1211), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n746), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1205), .A2(new_n751), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n748), .B1(G50), .B2(new_n831), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n791), .A2(G150), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n769), .B2(new_n1174), .C1(new_n772), .C2(new_n1165), .ZN(new_n1221));
  INV_X1    g1021(.A(G132), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1171), .A2(new_n777), .B1(new_n773), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(new_n785), .C2(G137), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT59), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n788), .A2(G159), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n317), .B2(new_n288), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n264), .A2(new_n773), .B1(new_n772), .B2(new_n355), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n317), .B(new_n288), .C1(new_n777), .C2(new_n247), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n836), .A2(new_n803), .B1(new_n774), .B2(new_n790), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n268), .A2(new_n769), .B1(new_n787), .B2(new_n463), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1235), .B(new_n1238), .C1(new_n784), .C2(new_n419), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT58), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1232), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1230), .B(new_n1241), .C1(new_n1240), .C2(new_n1239), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1219), .B1(new_n1242), .B2(new_n754), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1218), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1217), .A2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1216), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(G375));
  INV_X1    g1048(.A(new_n983), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1143), .B(new_n1152), .C1(new_n1145), .C2(new_n1149), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1154), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT116), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n883), .A2(new_n751), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n748), .B1(G68), .B2(new_n831), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n260), .B(new_n1058), .C1(G77), .C2(new_n788), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n785), .A2(G107), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n355), .A2(new_n773), .B1(new_n777), .B2(new_n803), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G294), .B2(new_n800), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n836), .A2(new_n805), .B1(new_n769), .B2(new_n264), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT117), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1255), .A2(new_n1256), .A3(new_n1258), .A4(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n784), .A2(new_n841), .B1(new_n202), .B2(new_n790), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n1262), .B(KEYINPUT118), .Z(new_n1263));
  AOI22_X1  g1063(.A1(G132), .A2(new_n800), .B1(new_n778), .B2(G137), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n317), .B1(G128), .B2(new_n793), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(G159), .A2(new_n1069), .B1(new_n788), .B2(new_n432), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n773), .A2(new_n1174), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1261), .B1(new_n1263), .B2(new_n1268), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1269), .A2(KEYINPUT119), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n767), .B1(new_n1269), .B2(KEYINPUT119), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1254), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1150), .A2(new_n747), .B1(new_n1253), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1252), .A2(new_n1273), .ZN(G381));
  INV_X1    g1074(.A(G390), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1045), .A2(new_n816), .A3(new_n1081), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n857), .A3(new_n1277), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(G381), .A2(G378), .A3(new_n1278), .A4(G387), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1247), .A2(new_n1279), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1280), .B(KEYINPUT120), .Z(G407));
  AOI21_X1  g1081(.A(new_n1184), .B1(new_n1161), .B2(new_n1155), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n671), .A2(G213), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1247), .A2(new_n1282), .A3(new_n1284), .ZN(new_n1285));
  XOR2_X1   g1085(.A(new_n1285), .B(KEYINPUT121), .Z(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(G213), .A3(G407), .ZN(G409));
  AOI21_X1  g1087(.A(new_n816), .B1(new_n1045), .B2(new_n1081), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1277), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1017), .A2(new_n1038), .A3(G390), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G390), .B1(new_n1017), .B2(new_n1038), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1290), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(new_n1275), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1017), .A2(new_n1038), .A3(G390), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1289), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G378), .B(new_n1246), .C1(new_n1213), .C2(new_n1215), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1214), .A2(new_n1249), .A3(new_n1211), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1210), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1206), .A2(new_n1207), .B1(new_n924), .B2(new_n910), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n747), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(KEYINPUT122), .A3(new_n1244), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT122), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1217), .B2(new_n1245), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1299), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1282), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1298), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1111), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1250), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1159), .A2(KEYINPUT60), .A3(new_n1152), .A4(new_n1143), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1309), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT123), .B1(new_n1313), .B2(new_n1273), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(KEYINPUT123), .A3(new_n1273), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1315), .A2(G384), .A3(new_n1316), .ZN(new_n1317));
  AND4_X1   g1117(.A1(KEYINPUT123), .A2(new_n1313), .A3(new_n857), .A4(new_n1273), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1308), .A2(new_n1283), .A3(new_n1320), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1321), .A2(KEYINPUT62), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(KEYINPUT62), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1322), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1313), .A2(KEYINPUT123), .A3(new_n1273), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(new_n1326), .A2(new_n1314), .A3(new_n857), .ZN(new_n1327));
  OAI21_X1  g1127(.A(KEYINPUT125), .B1(new_n1327), .B2(new_n1318), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1284), .A2(G2897), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT125), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1317), .A2(new_n1319), .A3(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1328), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1308), .A2(new_n1283), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1330), .B1(new_n1328), .B2(new_n1332), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1297), .B1(new_n1325), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT127), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1284), .B1(new_n1298), .B2(new_n1307), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(KEYINPUT63), .A3(new_n1320), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1293), .A2(new_n1296), .A3(new_n1323), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(KEYINPUT126), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT126), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1293), .A2(new_n1296), .A3(new_n1344), .A4(new_n1323), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1341), .B(new_n1346), .C1(new_n1335), .C2(new_n1336), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT63), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1321), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(KEYINPUT124), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT124), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1321), .A2(new_n1352), .A3(new_n1349), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1351), .A2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1339), .B1(new_n1348), .B2(new_n1354), .ZN(new_n1355));
  AOI211_X1 g1155(.A(KEYINPUT124), .B(KEYINPUT63), .C1(new_n1340), .C2(new_n1320), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1352), .B1(new_n1321), .B2(new_n1349), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  NOR3_X1   g1158(.A1(new_n1358), .A2(new_n1347), .A3(KEYINPUT127), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1338), .B1(new_n1355), .B2(new_n1359), .ZN(G405));
  NOR2_X1   g1160(.A1(new_n1247), .A2(G378), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1298), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1320), .ZN(new_n1363));
  OR3_X1    g1163(.A1(new_n1361), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1363), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1364), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1297), .ZN(new_n1367));
  XNOR2_X1  g1167(.A(new_n1366), .B(new_n1367), .ZN(G402));
endmodule


