//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT24), .B(G110), .Z(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n189), .A2(KEYINPUT23), .A3(G128), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT23), .B1(new_n189), .B2(G128), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n188), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G110), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT16), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  OR3_X1    g016(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(G146), .A3(new_n203), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n199), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT71), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n197), .A2(new_n198), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n191), .B2(new_n192), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n200), .A2(new_n205), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n207), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(KEYINPUT22), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(G137), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n214), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n218), .B(KEYINPUT72), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT25), .B1(new_n223), .B2(G902), .ZN(new_n224));
  INV_X1    g038(.A(G217), .ZN(new_n225));
  INV_X1    g039(.A(G902), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(G234), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n222), .A2(new_n228), .A3(new_n226), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n227), .A2(G902), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n231), .B(KEYINPUT73), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n237));
  INV_X1    g051(.A(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G137), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(G137), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n238), .B2(G137), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT11), .A3(G134), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n244), .A2(new_n246), .A3(new_n247), .A4(new_n239), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n205), .A2(G143), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(G146), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n205), .A2(KEYINPUT64), .A3(G143), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n187), .B1(new_n250), .B2(KEYINPUT1), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(G146), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n250), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G128), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n249), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n250), .A2(new_n259), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n252), .A2(G146), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT64), .B1(new_n205), .B2(G143), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n251), .A2(new_n252), .A3(G146), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n265), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT67), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n275), .B(new_n265), .C1(new_n269), .C2(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n244), .A2(new_n239), .A3(new_n246), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G131), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n248), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n263), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(G116), .B(G119), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT2), .B(G113), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n284), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(G101), .ZN(new_n291));
  NOR2_X1   g105(.A1(G237), .A2(G953), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G210), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n291), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n279), .A2(new_n248), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(new_n273), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n258), .A2(new_n262), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n248), .A3(new_n242), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n255), .A2(new_n271), .B1(new_n264), .B2(new_n260), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n280), .A3(KEYINPUT65), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n303), .B1(new_n302), .B2(new_n304), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT68), .B1(new_n281), .B2(KEYINPUT30), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n296), .B1(new_n274), .B2(new_n276), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n309));
  NOR4_X1   g123(.A1(new_n308), .A2(new_n309), .A3(new_n304), .A4(new_n263), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n305), .A2(new_n306), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n289), .B(new_n294), .C1(new_n311), .C2(new_n288), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n237), .B1(new_n312), .B2(KEYINPUT31), .ZN(new_n313));
  INV_X1    g127(.A(new_n289), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n300), .A2(new_n280), .A3(KEYINPUT65), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT65), .B1(new_n300), .B2(new_n280), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(new_n263), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT66), .B1(new_n317), .B2(KEYINPUT30), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n255), .A2(new_n271), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n275), .B1(new_n320), .B2(new_n265), .ZN(new_n321));
  INV_X1    g135(.A(new_n276), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n280), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT30), .A3(new_n299), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n309), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n281), .A2(KEYINPUT68), .A3(KEYINPUT30), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n318), .A2(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n314), .B1(new_n327), .B2(new_n287), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n328), .A2(KEYINPUT69), .A3(new_n329), .A4(new_n294), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n313), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n289), .B(KEYINPUT28), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n288), .B2(new_n317), .ZN(new_n333));
  INV_X1    g147(.A(new_n294), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n312), .A2(KEYINPUT31), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(G472), .A2(G902), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT32), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n236), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n312), .A2(KEYINPUT31), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n333), .A2(new_n334), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n313), .B2(new_n330), .ZN(new_n344));
  INV_X1    g158(.A(new_n337), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(KEYINPUT32), .A3(new_n337), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n340), .B1(new_n348), .B2(new_n236), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n328), .A2(new_n334), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n333), .A2(new_n294), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n287), .B1(new_n308), .B2(new_n263), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n332), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n294), .A2(KEYINPUT29), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n226), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G472), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n235), .B1(new_n349), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n273), .A2(G125), .ZN(new_n359));
  OR2_X1    g173(.A1(new_n359), .A2(KEYINPUT82), .ZN(new_n360));
  INV_X1    g174(.A(new_n298), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n202), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(KEYINPUT82), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n215), .A2(G224), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(KEYINPUT83), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n364), .B(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G104), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G107), .ZN(new_n369));
  INV_X1    g183(.A(G107), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G104), .ZN(new_n371));
  OAI21_X1  g185(.A(G101), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n371), .B1(new_n373), .B2(new_n369), .ZN(new_n374));
  INV_X1    g188(.A(G101), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n368), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT75), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(KEYINPUT75), .B(KEYINPUT3), .C1(new_n368), .C2(G107), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n374), .A2(new_n375), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n380), .A2(new_n381), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n372), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT77), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n378), .A2(new_n379), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(KEYINPUT76), .A3(new_n375), .A4(new_n374), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n380), .A2(new_n381), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n372), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n189), .A3(G116), .ZN(new_n393));
  OAI211_X1 g207(.A(G113), .B(new_n393), .C1(new_n283), .C2(new_n392), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n285), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n385), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n386), .A2(new_n374), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G101), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(new_n287), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(G110), .B(G122), .Z(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n404), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n397), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  AND4_X1   g224(.A1(new_n409), .A2(new_n403), .A3(new_n410), .A4(new_n404), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n406), .B1(new_n397), .B2(new_n402), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n412), .B2(new_n410), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n367), .B(new_n408), .C1(new_n411), .C2(new_n413), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n404), .B(KEYINPUT8), .Z(new_n415));
  INV_X1    g229(.A(new_n397), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n396), .B1(new_n389), .B2(new_n372), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT84), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n362), .A2(new_n359), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n365), .A2(KEYINPUT7), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n364), .A2(KEYINPUT7), .A3(new_n365), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n407), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n425), .B(new_n415), .C1(new_n416), .C2(new_n417), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n419), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n414), .A2(new_n226), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G210), .B1(G237), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n414), .A2(new_n226), .A3(new_n429), .A4(new_n427), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G214), .B1(G237), .B2(G902), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT9), .B(G234), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n226), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G221), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT74), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n400), .A2(new_n401), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n277), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n262), .B1(new_n260), .B2(new_n256), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n389), .A2(new_n372), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT10), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n385), .A2(KEYINPUT10), .A3(new_n298), .A4(new_n391), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n280), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n442), .A2(new_n296), .A3(new_n446), .A4(new_n448), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G140), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n215), .A2(G227), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n452), .B(new_n453), .Z(new_n454));
  AND3_X1   g268(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n390), .B1(new_n389), .B2(new_n372), .ZN(new_n456));
  INV_X1    g270(.A(new_n372), .ZN(new_n457));
  AOI211_X1 g271(.A(KEYINPUT77), .B(new_n457), .C1(new_n387), .C2(new_n388), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n361), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT79), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n461), .B(new_n361), .C1(new_n456), .C2(new_n458), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n444), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n296), .A2(KEYINPUT78), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n463), .A2(KEYINPUT12), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT12), .B1(new_n463), .B2(new_n464), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n451), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n454), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n440), .B(new_n455), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n451), .A2(new_n454), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n464), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n463), .A2(KEYINPUT12), .A3(new_n464), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n454), .B1(new_n450), .B2(new_n451), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n440), .B(new_n226), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT80), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n470), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n465), .B2(new_n466), .ZN(new_n481));
  INV_X1    g295(.A(new_n476), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT80), .A3(new_n440), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n469), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n440), .A2(new_n226), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI211_X1 g301(.A(new_n435), .B(new_n439), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G475), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n368), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT85), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n200), .A2(new_n492), .A3(KEYINPUT19), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT19), .B1(new_n200), .B2(new_n492), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n205), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT86), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n200), .A2(new_n492), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT19), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n493), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(new_n205), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n292), .A2(G143), .A3(G214), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(G143), .B1(new_n292), .B2(G214), .ZN(new_n506));
  OAI21_X1  g320(.A(G131), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n247), .A3(new_n504), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n497), .A2(new_n503), .A3(new_n207), .A4(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n200), .B(new_n205), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n504), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(new_n247), .ZN(new_n515));
  OAI221_X1 g329(.A(new_n512), .B1(new_n513), .B2(new_n515), .C1(new_n514), .C2(new_n507), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n491), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n507), .A2(new_n509), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(KEYINPUT17), .A3(G131), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n206), .A4(new_n207), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n516), .A3(new_n491), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n489), .B(new_n226), .C1(new_n517), .C2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(G146), .B1(new_n500), .B2(new_n493), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n207), .B(new_n510), .C1(new_n527), .C2(new_n502), .ZN(new_n528));
  INV_X1    g342(.A(new_n503), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n516), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n491), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n522), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n533), .A2(KEYINPUT87), .A3(new_n489), .A4(new_n226), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(new_n534), .A3(KEYINPUT20), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT20), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n524), .A2(new_n525), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n491), .B1(new_n521), .B2(new_n516), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n226), .B1(new_n523), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G475), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n535), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n535), .A2(new_n537), .A3(KEYINPUT88), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G478), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n549));
  XNOR2_X1  g363(.A(G128), .B(G143), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n252), .A2(G128), .ZN(new_n553));
  OAI21_X1  g367(.A(G134), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n549), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n551), .A2(new_n553), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n550), .A2(new_n551), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n556), .A2(KEYINPUT90), .A3(G134), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n550), .A2(new_n238), .ZN(new_n560));
  XNOR2_X1  g374(.A(G116), .B(G122), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G107), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n550), .B(new_n238), .ZN(new_n567));
  INV_X1    g381(.A(G116), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(KEYINPUT14), .A3(G122), .ZN(new_n569));
  INV_X1    g383(.A(new_n561), .ZN(new_n570));
  OAI211_X1 g384(.A(G107), .B(new_n569), .C1(new_n570), .C2(KEYINPUT14), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n567), .B(new_n571), .C1(G107), .C2(new_n570), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n562), .B1(new_n555), .B2(new_n558), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT91), .A3(new_n560), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n566), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n436), .A2(G217), .A3(new_n215), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(KEYINPUT92), .Z(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n566), .A2(new_n579), .A3(new_n572), .A4(new_n574), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n548), .B1(new_n581), .B2(new_n226), .ZN(new_n582));
  AOI211_X1 g396(.A(G902), .B(new_n547), .C1(new_n578), .C2(new_n580), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n215), .A2(G952), .ZN(new_n585));
  NAND2_X1  g399(.A1(G234), .A2(G237), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT21), .B(G898), .Z(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(G902), .A3(G953), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n545), .A2(new_n584), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n358), .A2(new_n488), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT93), .B(G101), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G3));
  AOI21_X1  g408(.A(new_n439), .B1(new_n485), .B2(new_n487), .ZN(new_n595));
  INV_X1    g409(.A(new_n235), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n545), .ZN(new_n598));
  AOI21_X1  g412(.A(G478), .B1(new_n581), .B2(new_n226), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n573), .A2(KEYINPUT91), .A3(new_n560), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT91), .B1(new_n573), .B2(new_n560), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT95), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT94), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n577), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n602), .A2(new_n603), .A3(new_n572), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n575), .B2(KEYINPUT95), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n580), .A2(KEYINPUT95), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT33), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n581), .A2(KEYINPUT33), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n599), .B1(new_n613), .B2(G478), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n598), .A2(new_n615), .A3(KEYINPUT96), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n545), .B2(new_n614), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n434), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n431), .B2(new_n432), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n590), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n336), .B2(new_n226), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n336), .B2(new_n337), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n597), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  NOR3_X1   g443(.A1(new_n622), .A2(new_n584), .A3(new_n541), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n597), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  XNOR2_X1  g447(.A(new_n214), .B(KEYINPUT97), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n221), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n233), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n230), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n626), .A2(KEYINPUT98), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n344), .B2(G902), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n638), .A3(new_n338), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n488), .A2(new_n591), .A3(new_n639), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT37), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n198), .ZN(G12));
  AOI21_X1  g460(.A(KEYINPUT32), .B1(new_n336), .B2(new_n337), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n339), .B(new_n345), .C1(new_n331), .C2(new_n335), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n236), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n650), .A3(new_n357), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n587), .B1(new_n589), .B2(G900), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n541), .A2(new_n584), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT99), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n655), .A2(new_n638), .A3(new_n621), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n595), .A2(new_n651), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  XOR2_X1   g472(.A(new_n433), .B(KEYINPUT38), .Z(new_n659));
  XOR2_X1   g473(.A(new_n652), .B(KEYINPUT39), .Z(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n595), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n659), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n328), .A2(new_n334), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n289), .A2(new_n334), .A3(new_n353), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n226), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n649), .A2(new_n650), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT100), .ZN(new_n672));
  INV_X1    g486(.A(new_n638), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n545), .A2(new_n620), .A3(new_n584), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT101), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n666), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  AOI21_X1  g492(.A(new_n673), .B1(new_n349), .B2(new_n357), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n545), .A2(new_n614), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n680), .B1(new_n681), .B2(new_n652), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n545), .A2(new_n614), .A3(KEYINPUT102), .A4(new_n653), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n679), .A2(new_n488), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT103), .B1(new_n483), .B2(new_n440), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n473), .A2(new_n474), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n476), .B1(new_n690), .B2(new_n480), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n689), .B(G469), .C1(new_n691), .C2(G902), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n479), .A2(new_n484), .ZN(new_n694));
  INV_X1    g508(.A(new_n439), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n358), .A2(new_n687), .A3(new_n623), .A4(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n623), .A2(new_n696), .A3(new_n651), .A4(new_n596), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT41), .Z(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(G113), .Z(G15));
  NAND3_X1  g516(.A1(new_n358), .A2(new_n630), .A3(new_n696), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  AND4_X1   g518(.A1(new_n621), .A2(new_n693), .A3(new_n694), .A4(new_n695), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n651), .A2(new_n705), .A3(new_n591), .A4(new_n638), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n189), .ZN(G21));
  AOI22_X1  g521(.A1(new_n313), .A2(new_n330), .B1(new_n334), .B2(new_n354), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n345), .B1(new_n708), .B2(new_n341), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n235), .A2(new_n625), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n674), .A2(new_n433), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n696), .A2(new_n590), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NOR3_X1   g527(.A1(new_n673), .A2(new_n625), .A3(new_n709), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n696), .A2(new_n684), .A3(new_n621), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  NOR2_X1   g530(.A1(new_n439), .A2(new_n620), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n431), .A2(new_n432), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n486), .B(KEYINPUT105), .Z(new_n719));
  AOI21_X1  g533(.A(new_n718), .B1(new_n485), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n684), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT107), .B1(new_n647), .B2(new_n648), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n346), .A2(new_n723), .A3(new_n347), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n724), .A3(new_n357), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n725), .A2(KEYINPUT108), .A3(new_n596), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT108), .B1(new_n725), .B2(new_n596), .ZN(new_n727));
  OAI211_X1 g541(.A(KEYINPUT42), .B(new_n721), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n720), .A2(new_n651), .A3(new_n596), .A4(new_n684), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n729), .A2(KEYINPUT106), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT106), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  NAND3_X1  g548(.A1(new_n358), .A2(new_n655), .A3(new_n720), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT109), .B(G134), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G36));
  NAND2_X1  g551(.A1(new_n615), .A2(new_n545), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT43), .ZN(new_n739));
  OR3_X1    g553(.A1(new_n739), .A2(new_n626), .A3(new_n673), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT112), .Z(new_n743));
  NOR2_X1   g557(.A1(new_n433), .A2(new_n620), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n741), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n455), .B1(new_n467), .B2(new_n468), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(G469), .A3(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(new_n719), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n751));
  OR3_X1    g565(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT46), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n750), .B2(KEYINPUT46), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n719), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n694), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(KEYINPUT110), .A3(new_n694), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n752), .A2(new_n753), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n695), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n660), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n759), .A2(KEYINPUT47), .A3(new_n695), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n684), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n651), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n767), .A2(new_n235), .A3(new_n744), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  AND2_X1   g585(.A1(new_n693), .A2(new_n694), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n596), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n774), .A2(new_n620), .A3(new_n439), .A4(new_n738), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT113), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n672), .B1(new_n773), .B2(new_n772), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n659), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n726), .A2(new_n727), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n587), .ZN(new_n781));
  INV_X1    g595(.A(new_n718), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n772), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n739), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT122), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT48), .Z(new_n787));
  NOR3_X1   g601(.A1(new_n672), .A2(new_n235), .A3(new_n783), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n545), .A3(new_n614), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n710), .A2(new_n781), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n739), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n620), .A3(new_n659), .A4(new_n696), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n792), .A2(KEYINPUT50), .B1(new_n784), .B2(new_n714), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n789), .B(new_n793), .C1(KEYINPUT50), .C2(new_n792), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n772), .A2(new_n439), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n765), .A2(new_n766), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n791), .A2(new_n744), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT121), .Z(new_n798));
  AOI21_X1  g612(.A(new_n794), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(KEYINPUT51), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n585), .B1(new_n799), .B2(KEYINPUT51), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n672), .A2(new_n235), .A3(new_n619), .A4(new_n783), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n787), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n673), .A2(KEYINPUT116), .A3(new_n652), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n638), .B2(new_n653), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n671), .A2(new_n807), .A3(new_n711), .A4(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n485), .A2(new_n719), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n439), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n806), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n715), .A2(new_n657), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n715), .B2(new_n657), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n813), .B(new_n685), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n595), .A2(new_n651), .A3(new_n621), .A4(new_n638), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n657), .B(new_n715), .C1(new_n819), .C2(new_n768), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n671), .A2(new_n807), .A3(new_n711), .A4(new_n809), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n439), .A3(new_n811), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n818), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n817), .A2(KEYINPUT118), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT118), .B1(new_n817), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n584), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n545), .A2(KEYINPUT114), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT114), .B1(new_n545), .B2(new_n614), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n545), .A2(new_n827), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n622), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n595), .A3(new_n596), .A4(new_n626), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n592), .A2(new_n644), .A3(new_n712), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n706), .B1(new_n697), .B2(new_n699), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n625), .A2(new_n709), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n720), .A2(new_n684), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n827), .A2(new_n653), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n595), .A2(new_n651), .A3(new_n744), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n839), .B2(new_n541), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n638), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n834), .A2(new_n835), .A3(new_n703), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n733), .A2(new_n735), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n805), .B1(new_n826), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT52), .B1(new_n820), .B2(new_n822), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n715), .A2(new_n657), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n810), .A2(new_n812), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n806), .A4(new_n685), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n842), .A2(new_n843), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT53), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n804), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n844), .B(KEYINPUT53), .C1(new_n825), .C2(new_n824), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n825), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n817), .A2(KEYINPUT118), .A3(new_n823), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(KEYINPUT120), .A3(KEYINPUT53), .A4(new_n844), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n852), .B2(KEYINPUT53), .ZN(new_n863));
  INV_X1    g677(.A(new_n843), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n834), .A2(new_n703), .A3(new_n835), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n847), .A2(new_n850), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n841), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(KEYINPUT119), .A3(new_n805), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n857), .A2(new_n861), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n854), .B1(new_n869), .B2(new_n804), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n791), .A2(new_n705), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n803), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n778), .B1(new_n872), .B2(new_n873), .ZN(G75));
  OAI21_X1  g688(.A(new_n408), .B1(new_n411), .B2(new_n413), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n367), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT55), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(G210), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n869), .A2(new_n879), .A3(new_n226), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n880), .B2(KEYINPUT56), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n857), .A2(new_n861), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n863), .A2(new_n868), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(G902), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n882), .B(new_n877), .C1(new_n886), .C2(new_n879), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n215), .A2(G952), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n881), .A2(new_n887), .A3(new_n889), .ZN(G51));
  XOR2_X1   g704(.A(new_n719), .B(KEYINPUT57), .Z(new_n891));
  AND3_X1   g705(.A1(new_n883), .A2(new_n804), .A3(new_n884), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n804), .B1(new_n883), .B2(new_n884), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n691), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n886), .A2(new_n749), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n888), .B1(new_n896), .B2(new_n897), .ZN(G54));
  NAND4_X1  g712(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n522), .A3(new_n532), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n869), .A2(new_n226), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .A4(new_n533), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n900), .A2(new_n902), .A3(new_n889), .ZN(G60));
  INV_X1    g717(.A(new_n611), .ZN(new_n904));
  INV_X1    g718(.A(new_n612), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(G478), .A2(G902), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT59), .Z(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n870), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n906), .ZN(new_n910));
  INV_X1    g724(.A(new_n908), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n910), .B(new_n911), .C1(new_n892), .C2(new_n893), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n909), .A2(new_n912), .A3(new_n889), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n223), .B1(new_n869), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT124), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n883), .B2(new_n884), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n636), .B(KEYINPUT123), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n888), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n921), .B(new_n223), .C1(new_n869), .C2(new_n915), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n917), .A2(new_n920), .A3(KEYINPUT61), .A4(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n915), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n885), .A2(new_n924), .A3(new_n919), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n916), .A3(new_n889), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n928), .ZN(G66));
  AOI21_X1  g743(.A(new_n215), .B1(new_n588), .B2(G224), .ZN(new_n930));
  INV_X1    g744(.A(new_n865), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(new_n215), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n875), .B1(G898), .B2(new_n215), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n932), .B(new_n933), .Z(G69));
  NAND2_X1  g748(.A1(G227), .A2(G900), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(G953), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n501), .B(KEYINPUT125), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n311), .B(new_n937), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n815), .A2(new_n816), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n939), .A2(new_n685), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n677), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT62), .ZN(new_n942));
  INV_X1    g756(.A(new_n831), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n663), .A2(new_n358), .A3(new_n744), .A4(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n770), .A2(new_n762), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n938), .B1(new_n948), .B2(G953), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n215), .A2(G900), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n761), .A2(new_n711), .A3(new_n780), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n770), .A2(new_n762), .A3(new_n735), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n940), .A2(new_n733), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n951), .B(new_n952), .C1(new_n956), .C2(G953), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n936), .B(new_n949), .C1(new_n958), .C2(new_n938), .ZN(new_n959));
  OAI211_X1 g773(.A(G953), .B(new_n935), .C1(new_n957), .C2(new_n938), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(G72));
  NOR3_X1   g775(.A1(new_n942), .A2(new_n947), .A3(new_n931), .ZN(new_n962));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n667), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n350), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n954), .A2(new_n931), .A3(new_n955), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n846), .A2(new_n853), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n967), .A2(new_n667), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n964), .A3(new_n971), .ZN(new_n972));
  AND4_X1   g786(.A1(new_n889), .A2(new_n966), .A3(new_n969), .A4(new_n972), .ZN(G57));
endmodule


