//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT70), .ZN(new_n207));
  INV_X1    g006(.A(G134gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT69), .ZN(new_n209));
  XNOR2_X1  g008(.A(G113gat), .B(G120gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n211));
  INV_X1    g010(.A(G120gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G113gat), .ZN(new_n213));
  INV_X1    g012(.A(G113gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G120gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n208), .ZN(new_n218));
  INV_X1    g017(.A(G127gat), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n211), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(new_n211), .B2(new_n218), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n207), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n209), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(new_n216), .B2(new_n217), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n210), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n225));
  OAI21_X1  g024(.A(G127gat), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n218), .A3(new_n219), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(KEYINPUT70), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G141gat), .B(G148gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT77), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT77), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT77), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(G155gat), .A3(G162gat), .ZN(new_n236));
  INV_X1    g035(.A(G155gat), .ZN(new_n237));
  INV_X1    g036(.A(G162gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n242));
  AND2_X1   g041(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n243), .A2(new_n244), .A3(new_n238), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n242), .B1(new_n245), .B2(new_n230), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT78), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n237), .ZN(new_n248));
  NAND2_X1  g047(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(G162gat), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT79), .A3(KEYINPUT2), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n229), .B1(new_n233), .B2(new_n239), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n241), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n222), .A2(new_n228), .A3(new_n254), .A4(KEYINPUT4), .ZN(new_n255));
  INV_X1    g054(.A(new_n229), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n233), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n246), .B2(new_n251), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT3), .B1(new_n259), .B2(new_n241), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n220), .A2(new_n221), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n250), .A2(KEYINPUT79), .A3(KEYINPUT2), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT79), .B1(new_n250), .B2(KEYINPUT2), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n253), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g064(.A(new_n241), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n260), .A2(new_n261), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G225gat), .A2(G233gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n255), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n266), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT80), .B1(new_n272), .B2(new_n261), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT80), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n226), .A2(new_n227), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n254), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n271), .A2(new_n279), .A3(KEYINPUT81), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT81), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT4), .B1(new_n273), .B2(new_n276), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n281), .B1(new_n270), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT82), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n254), .A2(new_n275), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n286), .B1(new_n273), .B2(new_n276), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n287), .B2(new_n269), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n261), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n254), .A2(new_n274), .A3(new_n275), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n274), .B1(new_n254), .B2(new_n275), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n269), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(KEYINPUT82), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n288), .A2(new_n294), .A3(KEYINPUT5), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT83), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n269), .B1(new_n277), .B2(new_n289), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(KEYINPUT82), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(KEYINPUT83), .A3(new_n288), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n284), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n222), .A2(new_n228), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n278), .B1(new_n303), .B2(new_n272), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n268), .B(new_n304), .C1(new_n277), .C2(new_n278), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n305), .A2(KEYINPUT5), .A3(new_n293), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n206), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n280), .A2(new_n283), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT83), .B1(new_n300), .B2(new_n288), .ZN(new_n309));
  AND4_X1   g108(.A1(KEYINPUT83), .A2(new_n288), .A3(new_n294), .A4(KEYINPUT5), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n206), .ZN(new_n312));
  INV_X1    g111(.A(new_n306), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT6), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n307), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(KEYINPUT6), .B(new_n206), .C1(new_n302), .C2(new_n306), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319));
  AND2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(G169gat), .ZN(new_n321));
  INV_X1    g120(.A(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n320), .B1(new_n323), .B2(KEYINPUT26), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(KEYINPUT26), .B2(new_n323), .ZN(new_n325));
  NAND2_X1  g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(G183gat), .ZN(new_n327));
  OR3_X1    g126(.A1(new_n327), .A2(KEYINPUT68), .A3(KEYINPUT27), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G183gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT68), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(KEYINPUT27), .ZN(new_n332));
  NOR2_X1   g131(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n328), .A2(new_n331), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n330), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT28), .B1(new_n335), .B2(G190gat), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n325), .A2(new_n326), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n320), .B1(new_n323), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n339), .A2(G169gat), .ZN(new_n347));
  AND2_X1   g146(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n340), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT66), .B1(new_n341), .B2(KEYINPUT67), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n354), .A2(new_n326), .ZN(new_n355));
  NAND3_X1  g154(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT67), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT24), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n344), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n352), .B1(new_n360), .B2(KEYINPUT23), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n340), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n353), .A2(KEYINPUT65), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n351), .A2(new_n364), .A3(new_n352), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n338), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n319), .B1(new_n366), .B2(KEYINPUT29), .ZN(new_n367));
  XNOR2_X1  g166(.A(G197gat), .B(G204gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT22), .ZN(new_n369));
  INV_X1    g168(.A(G211gat), .ZN(new_n370));
  INV_X1    g169(.A(G218gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G211gat), .B(G218gat), .Z(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT75), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n368), .A2(new_n372), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(KEYINPUT75), .A3(new_n374), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n353), .A2(KEYINPUT65), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n359), .A2(new_n362), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n365), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n337), .ZN(new_n383));
  INV_X1    g182(.A(new_n319), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n367), .A2(new_n379), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n379), .B1(new_n367), .B2(new_n385), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n386), .A2(new_n387), .ZN(new_n393));
  INV_X1    g192(.A(new_n391), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT30), .A3(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n388), .B2(new_n391), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n392), .A2(new_n395), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT76), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n318), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n267), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n379), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n267), .A2(KEYINPUT86), .A3(new_n406), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n265), .B1(new_n410), .B2(KEYINPUT29), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(new_n272), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT87), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n412), .A2(new_n415), .A3(KEYINPUT87), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n379), .B1(new_n267), .B2(new_n406), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n373), .A2(new_n374), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n406), .B1(new_n373), .B2(new_n374), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n265), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n272), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n421), .B2(new_n422), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n413), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n420), .A2(KEYINPUT88), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n412), .A2(new_n415), .A3(KEYINPUT87), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT87), .B1(new_n412), .B2(new_n415), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT31), .B(G50gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT84), .ZN(new_n438));
  XOR2_X1   g237(.A(G78gat), .B(G106gat), .Z(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  AOI21_X1  g239(.A(new_n431), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n440), .ZN(new_n442));
  AOI211_X1 g241(.A(G22gat), .B(new_n442), .C1(new_n434), .C2(new_n435), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n430), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT88), .B1(new_n420), .B2(new_n429), .ZN(new_n445));
  OAI21_X1  g244(.A(G22gat), .B1(new_n445), .B2(new_n442), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n436), .A2(new_n431), .A3(new_n440), .ZN(new_n447));
  INV_X1    g246(.A(new_n430), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT71), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n383), .B2(new_n303), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n366), .A2(KEYINPUT71), .A3(new_n228), .A4(new_n222), .ZN(new_n452));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n383), .A2(new_n303), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n455), .A2(KEYINPUT73), .A3(KEYINPUT34), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT34), .B1(new_n455), .B2(KEYINPUT73), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n460));
  INV_X1    g259(.A(new_n453), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G15gat), .B(G43gat), .Z(new_n465));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT32), .ZN(new_n469));
  AOI211_X1 g268(.A(KEYINPUT72), .B(new_n469), .C1(new_n460), .C2(new_n461), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT72), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n462), .B2(KEYINPUT32), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n468), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n469), .B1(new_n460), .B2(new_n461), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(KEYINPUT33), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n459), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n464), .B(new_n467), .C1(new_n471), .C2(new_n474), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n458), .B(new_n476), .C1(new_n479), .C2(new_n470), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n444), .A2(new_n449), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT35), .B1(new_n405), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT74), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n480), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n485), .B2(KEYINPUT74), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n396), .A2(new_n400), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT35), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n444), .A2(new_n449), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n486), .A2(new_n318), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n444), .A2(new_n449), .ZN(new_n493));
  INV_X1    g292(.A(new_n307), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT39), .B1(new_n292), .B2(new_n293), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n305), .A2(new_n293), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n497), .A2(KEYINPUT39), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n312), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n499), .A2(KEYINPUT40), .A3(new_n312), .A4(new_n500), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n493), .B1(new_n494), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n391), .B1(new_n393), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n393), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT91), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n393), .A2(new_n512), .A3(new_n509), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT38), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n514), .A2(new_n515), .B1(new_n394), .B2(new_n393), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n316), .A2(new_n517), .A3(new_n317), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n518), .B2(KEYINPUT92), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n316), .A2(new_n517), .A3(new_n520), .A4(new_n317), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n506), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n484), .ZN(new_n523));
  INV_X1    g322(.A(new_n480), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n462), .A2(KEYINPUT32), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n474), .A2(new_n471), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n526), .A2(new_n467), .A3(new_n527), .A4(new_n464), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n458), .B1(new_n528), .B2(new_n476), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT74), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT36), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n485), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n403), .B1(new_n316), .B2(new_n317), .ZN(new_n534));
  OAI22_X1  g333(.A1(new_n531), .A2(new_n533), .B1(new_n493), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n492), .B1(new_n522), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT103), .ZN(new_n537));
  INV_X1    g336(.A(G92gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n203), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(KEYINPUT103), .A2(G85gat), .A3(G92gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n539), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G99gat), .ZN(new_n543));
  INV_X1    g342(.A(G106gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT8), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n203), .A2(new_n538), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT104), .ZN(new_n548));
  XOR2_X1   g347(.A(G99gat), .B(G106gat), .Z(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n549), .A2(new_n548), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n542), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n542), .B2(new_n550), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G43gat), .B(G50gat), .Z(new_n555));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G43gat), .B(G50gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT15), .ZN(new_n559));
  OR3_X1    g358(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n557), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G29gat), .A2(G36gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT95), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(G29gat), .A3(G36gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT96), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n560), .A2(KEYINPUT94), .A3(new_n561), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n573), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n572), .A2(new_n574), .A3(new_n567), .A4(new_n565), .ZN(new_n575));
  INV_X1    g374(.A(new_n559), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n554), .A2(new_n578), .B1(KEYINPUT41), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n571), .A2(KEYINPUT17), .A3(new_n577), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n552), .A2(new_n553), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G134gat), .B(G162gat), .Z(new_n587));
  AND2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n590));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n588), .B2(new_n589), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n597), .A2(KEYINPUT99), .ZN(new_n598));
  XOR2_X1   g397(.A(G57gat), .B(G64gat), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(KEYINPUT99), .ZN(new_n600));
  XNOR2_X1  g399(.A(G71gat), .B(G78gat), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT100), .ZN(new_n603));
  INV_X1    g402(.A(new_n601), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT9), .B1(new_n599), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n611));
  XOR2_X1   g410(.A(G127gat), .B(G155gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n617));
  XNOR2_X1  g416(.A(G15gat), .B(G22gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT16), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(G1gat), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(G1gat), .B2(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(G8gat), .ZN(new_n622));
  INV_X1    g421(.A(G8gat), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n620), .B(new_n623), .C1(G1gat), .C2(new_n618), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G231gat), .ZN(new_n626));
  INV_X1    g425(.A(G233gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n617), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n617), .B2(new_n625), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n616), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n615), .A3(new_n630), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n614), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G183gat), .B(G211gat), .Z(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  NAND3_X1  g439(.A1(new_n633), .A2(new_n614), .A3(new_n635), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n636), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n596), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n609), .A2(new_n584), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n603), .B(new_n608), .C1(new_n553), .C2(new_n552), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n647), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n648), .A2(new_n656), .A3(new_n649), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n610), .A2(new_n554), .A3(KEYINPUT10), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(KEYINPUT105), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n661));
  AOI211_X1 g460(.A(new_n661), .B(new_n655), .C1(new_n657), .C2(new_n658), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n654), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g464(.A(KEYINPUT106), .B(new_n654), .C1(new_n660), .C2(new_n662), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n653), .B1(new_n659), .B2(new_n650), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n646), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n622), .A2(new_n624), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n578), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n563), .A2(new_n570), .B1(new_n576), .B2(new_n575), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n625), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(G229gat), .A2(G233gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT13), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n578), .A2(new_n672), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n583), .A2(new_n625), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n677), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(KEYINPUT18), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n582), .A2(new_n625), .A3(new_n583), .ZN(new_n688));
  INV_X1    g487(.A(new_n686), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n688), .A2(new_n677), .A3(new_n681), .A4(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n680), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT93), .ZN(new_n692));
  XNOR2_X1  g491(.A(G113gat), .B(G141gat), .ZN(new_n693));
  INV_X1    g492(.A(G197gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT11), .B(G169gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT12), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n691), .A2(new_n692), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n691), .B2(new_n692), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n671), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n536), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n318), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g508(.A1(new_n705), .A2(new_n488), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT42), .B1(new_n710), .B2(new_n623), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT107), .B(KEYINPUT16), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G8gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  MUX2_X1   g513(.A(KEYINPUT42), .B(new_n711), .S(new_n714), .Z(G1325gat));
  INV_X1    g514(.A(G15gat), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n483), .B1(new_n478), .B2(new_n480), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n532), .B1(new_n717), .B2(new_n484), .ZN(new_n718));
  INV_X1    g517(.A(new_n533), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n486), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n716), .B2(new_n722), .ZN(G1326gat));
  NOR2_X1   g522(.A1(new_n705), .A2(new_n493), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT43), .B(G22gat), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1327gat));
  NAND2_X1  g525(.A1(new_n536), .A2(new_n596), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n642), .A2(new_n645), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(new_n702), .A3(new_n670), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n318), .A2(G29gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT108), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(new_n735), .A3(new_n732), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n734), .A2(new_n736), .A3(KEYINPUT45), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n734), .B2(new_n736), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(G29gat), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT110), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT110), .B1(new_n594), .B2(new_n595), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n536), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n596), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n518), .A2(KEYINPUT92), .ZN(new_n748));
  INV_X1    g547(.A(new_n516), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n521), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n506), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n493), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n718), .A2(new_n719), .B1(new_n405), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n747), .B1(new_n755), .B2(new_n492), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n746), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT109), .B1(new_n700), .B2(new_n701), .ZN(new_n759));
  INV_X1    g558(.A(new_n698), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n680), .A2(new_n687), .A3(new_n690), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(KEYINPUT93), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(new_n763), .A3(new_n699), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n766), .A2(new_n728), .A3(new_n669), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT111), .B1(new_n758), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n757), .B1(new_n536), .B2(new_n596), .ZN(new_n770));
  INV_X1    g569(.A(new_n745), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n755), .B2(new_n492), .ZN(new_n772));
  OAI211_X1 g571(.A(KEYINPUT111), .B(new_n767), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n318), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n739), .B1(new_n740), .B2(new_n774), .ZN(G1328gat));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  INV_X1    g575(.A(G36gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n731), .A2(new_n777), .A3(new_n487), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(KEYINPUT46), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(KEYINPUT46), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n778), .A2(new_n776), .A3(KEYINPUT46), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n488), .B1(new_n769), .B2(new_n773), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n781), .B(new_n782), .C1(new_n783), .C2(new_n777), .ZN(G1329gat));
  NAND2_X1  g583(.A1(new_n758), .A2(new_n767), .ZN(new_n785));
  OAI21_X1  g584(.A(G43gat), .B1(new_n785), .B2(new_n720), .ZN(new_n786));
  INV_X1    g585(.A(new_n486), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(G43gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n731), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(KEYINPUT47), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n789), .ZN(new_n791));
  INV_X1    g590(.A(new_n720), .ZN(new_n792));
  INV_X1    g591(.A(new_n773), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n768), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n794), .B2(G43gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n790), .B1(new_n795), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g595(.A(G50gat), .B1(new_n785), .B2(new_n493), .ZN(new_n797));
  NOR4_X1   g596(.A1(new_n727), .A2(G50gat), .A3(new_n493), .A4(new_n730), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(KEYINPUT48), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n753), .B1(new_n768), .B2(new_n793), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n798), .B1(new_n801), .B2(G50gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n802), .B2(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g602(.A1(new_n646), .A2(new_n669), .A3(new_n766), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n536), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n318), .ZN(new_n806));
  XOR2_X1   g605(.A(KEYINPUT113), .B(G57gat), .Z(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1332gat));
  NOR2_X1   g607(.A1(new_n805), .A2(new_n488), .ZN(new_n809));
  NOR2_X1   g608(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n810));
  AND2_X1   g609(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n809), .B2(new_n810), .ZN(G1333gat));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n805), .A2(new_n787), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT114), .ZN(new_n816));
  INV_X1    g615(.A(G71gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n805), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n817), .B1(new_n819), .B2(new_n792), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n814), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g621(.A(KEYINPUT50), .B(new_n820), .C1(new_n816), .C2(new_n817), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(G1334gat));
  NAND2_X1  g623(.A1(new_n819), .A2(new_n753), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g625(.A1(new_n729), .A2(new_n766), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n670), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n758), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n707), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G85gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n727), .A2(new_n827), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n707), .A2(new_n203), .A3(new_n669), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(G1336gat));
  NAND3_X1  g635(.A1(new_n758), .A2(new_n487), .A3(new_n828), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(G92gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n669), .A2(new_n538), .A3(new_n487), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n838), .B(new_n842), .C1(new_n834), .C2(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1337gat));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n792), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G99gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n486), .A2(new_n543), .A3(new_n669), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n834), .B2(new_n847), .ZN(G1338gat));
  NAND3_X1  g647(.A1(new_n758), .A2(new_n753), .A3(new_n828), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G106gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n493), .A2(G106gat), .A3(new_n670), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT115), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n834), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT53), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n850), .B(new_n855), .C1(new_n834), .C2(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1339gat));
  NAND3_X1  g656(.A1(new_n646), .A2(new_n670), .A3(new_n766), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n657), .A2(new_n658), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT54), .B1(new_n860), .B2(new_n647), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n647), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n661), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n659), .A2(KEYINPUT105), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n653), .B1(new_n862), .B2(KEYINPUT54), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT55), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n866), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n660), .A2(new_n662), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n861), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n765), .A2(new_n872), .A3(new_n667), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n688), .A2(new_n681), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n676), .A2(new_n679), .B1(new_n874), .B2(new_n677), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n761), .A2(new_n698), .B1(new_n875), .B2(new_n697), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n669), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n744), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n867), .A2(new_n871), .B1(new_n665), .B2(new_n666), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n743), .A3(new_n876), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n859), .B1(new_n882), .B2(new_n729), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n318), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n787), .A2(new_n753), .A3(new_n487), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G113gat), .B1(new_n887), .B2(new_n703), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n883), .A2(new_n481), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n318), .A2(new_n487), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT116), .Z(new_n892));
  NAND2_X1  g691(.A1(new_n765), .A2(new_n214), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(G1340gat));
  OAI21_X1  g693(.A(G120gat), .B1(new_n887), .B2(new_n670), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n669), .A2(new_n212), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n892), .B2(new_n896), .ZN(G1341gat));
  XOR2_X1   g696(.A(KEYINPUT69), .B(G127gat), .Z(new_n898));
  NAND3_X1  g697(.A1(new_n886), .A2(new_n728), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  INV_X1    g701(.A(new_n891), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n898), .B1(new_n903), .B2(new_n728), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(G1342gat));
  INV_X1    g704(.A(new_n481), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n747), .A2(new_n487), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n884), .A2(new_n208), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT56), .Z(new_n909));
  OAI21_X1  g708(.A(G134gat), .B1(new_n887), .B2(new_n747), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1343gat));
  AOI22_X1  g710(.A1(new_n880), .A2(new_n702), .B1(new_n669), .B2(new_n876), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n881), .B1(new_n912), .B2(new_n596), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n859), .B1(new_n913), .B2(new_n729), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT57), .B1(new_n914), .B2(new_n493), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n720), .A2(new_n890), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n743), .B1(new_n873), .B2(new_n877), .ZN(new_n918));
  INV_X1    g717(.A(new_n881), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n729), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n858), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n753), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(KEYINPUT57), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(G141gat), .B1(new_n925), .B2(new_n703), .ZN(new_n926));
  INV_X1    g725(.A(new_n922), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n916), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(G141gat), .A3(new_n703), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(KEYINPUT58), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT58), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n924), .A2(new_n765), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n929), .B1(new_n933), .B2(G141gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n932), .B2(new_n934), .ZN(G1344gat));
  INV_X1    g734(.A(new_n928), .ZN(new_n936));
  INV_X1    g735(.A(G148gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n937), .A3(new_n669), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(KEYINPUT59), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(new_n925), .B2(new_n670), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT118), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n916), .B(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT57), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n671), .A2(new_n702), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n880), .A2(new_n596), .A3(new_n876), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n947), .B1(new_n912), .B2(new_n596), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(new_n729), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n949), .B2(new_n493), .ZN(new_n950));
  AOI211_X1 g749(.A(new_n945), .B(new_n493), .C1(new_n920), .C2(new_n858), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n922), .A2(KEYINPUT120), .A3(new_n945), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n669), .B(new_n944), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n937), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n942), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n938), .B1(new_n941), .B2(new_n959), .ZN(G1345gat));
  NAND2_X1  g759(.A1(new_n936), .A2(new_n728), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n248), .A2(new_n249), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n729), .A2(new_n962), .ZN(new_n963));
  AOI22_X1  g762(.A1(new_n961), .A2(new_n962), .B1(new_n924), .B2(new_n963), .ZN(G1346gat));
  OAI21_X1  g763(.A(G162gat), .B1(new_n925), .B2(new_n744), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n922), .A2(new_n792), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n966), .A2(new_n238), .A3(new_n707), .A4(new_n907), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1347gat));
  NOR2_X1   g767(.A1(new_n707), .A2(new_n488), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n889), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n321), .A3(new_n765), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT122), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n787), .A2(new_n707), .A3(new_n488), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n974), .A2(new_n493), .A3(new_n921), .A4(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(G169gat), .B1(new_n976), .B2(new_n703), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n972), .A2(new_n977), .ZN(G1348gat));
  NAND2_X1  g777(.A1(new_n970), .A2(new_n669), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n322), .ZN(new_n980));
  OR3_X1    g779(.A1(new_n670), .A2(new_n349), .A3(new_n348), .ZN(new_n981));
  OAI22_X1  g780(.A1(new_n980), .A2(KEYINPUT124), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n982), .B1(KEYINPUT124), .B2(new_n980), .ZN(G1349gat));
  OAI21_X1  g782(.A(G183gat), .B1(new_n976), .B2(new_n729), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n729), .A2(new_n335), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n986), .A2(KEYINPUT125), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n986), .A2(KEYINPUT125), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g789(.A1(new_n970), .A2(new_n343), .A3(new_n743), .ZN(new_n991));
  OAI21_X1  g790(.A(G190gat), .B1(new_n976), .B2(new_n747), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n992), .A2(KEYINPUT61), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n992), .A2(KEYINPUT61), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(G1351gat));
  NAND2_X1  g794(.A1(new_n966), .A2(new_n969), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n996), .A2(G197gat), .A3(new_n766), .ZN(new_n997));
  XOR2_X1   g796(.A(new_n997), .B(KEYINPUT126), .Z(new_n998));
  OR2_X1    g797(.A1(new_n953), .A2(new_n954), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n720), .A2(new_n969), .ZN(new_n1000));
  INV_X1    g799(.A(new_n1000), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n1002), .A2(new_n702), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n998), .B1(new_n1003), .B2(new_n694), .ZN(G1352gat));
  NOR3_X1   g803(.A1(new_n996), .A2(G204gat), .A3(new_n670), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT62), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n999), .A2(new_n669), .A3(new_n1001), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(G204gat), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1006), .A2(new_n1008), .ZN(G1353gat));
  INV_X1    g808(.A(new_n996), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1010), .A2(new_n370), .A3(new_n728), .ZN(new_n1011));
  OAI211_X1 g810(.A(new_n728), .B(new_n1001), .C1(new_n953), .C2(new_n954), .ZN(new_n1012));
  AND3_X1   g811(.A1(new_n1012), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1013));
  AOI21_X1  g812(.A(KEYINPUT63), .B1(new_n1012), .B2(G211gat), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g816(.A(KEYINPUT127), .B(new_n1011), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1017), .A2(new_n1018), .ZN(G1354gat));
  AOI21_X1  g818(.A(G218gat), .B1(new_n1010), .B2(new_n743), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n747), .A2(new_n371), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1020), .B1(new_n1002), .B2(new_n1021), .ZN(G1355gat));
endmodule


