//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155, new_n1156;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n464), .B1(new_n466), .B2(G101), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n460), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n460), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n478), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n461), .B2(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n488), .B(new_n491), .C1(new_n462), .C2(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n460), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n481), .A2(G126), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n493), .B2(new_n498), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G50), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n504), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n502), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n506), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  NAND2_X1  g093(.A1(new_n505), .A2(G51), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT69), .B(G89), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n521), .A2(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n503), .A2(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n527), .A2(G90), .B1(new_n505), .B2(G52), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(new_n512), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n516), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n536), .B1(new_n535), .B2(new_n534), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n530), .A2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  AOI22_X1  g114(.A1(new_n527), .A2(G81), .B1(new_n505), .B2(G43), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT73), .Z(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n532), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n516), .B1(new_n544), .B2(KEYINPUT72), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n545), .B1(KEYINPUT72), .B2(new_n544), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n505), .A2(G53), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OR3_X1    g135(.A1(new_n513), .A2(KEYINPUT75), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT75), .B1(new_n513), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n532), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n561), .A2(new_n562), .B1(G651), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n559), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  OAI21_X1  g144(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(new_n505), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n527), .A2(G87), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G288));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n505), .A2(new_n577), .A3(G48), .ZN(new_n578));
  INV_X1    g153(.A(new_n504), .ZN(new_n579));
  NOR2_X1   g154(.A1(KEYINPUT6), .A2(G651), .ZN(new_n580));
  OAI211_X1 g155(.A(G48), .B(G543), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT77), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n578), .A2(new_n582), .B1(G86), .B2(new_n527), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n510), .B2(new_n511), .ZN(new_n585));
  AND2_X1   g160(.A1(G73), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n583), .B1(new_n589), .B2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n505), .A2(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n513), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n516), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(new_n527), .A2(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT10), .Z(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n532), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n505), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G284));
  OAI21_X1  g183(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  XNOR2_X1  g187(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g188(.A(new_n605), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n547), .A2(new_n606), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n605), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n475), .A2(new_n466), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  XOR2_X1   g197(.A(KEYINPUT79), .B(KEYINPUT13), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT80), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n477), .A2(G135), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n481), .A2(G123), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n460), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2096), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n624), .B2(new_n625), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n627), .A2(new_n634), .ZN(G156));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT82), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2451), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n640), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2454), .Z(new_n649));
  OR2_X1    g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT83), .Z(new_n655));
  NOR2_X1   g230(.A1(G2072), .A2(G2078), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n445), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(KEYINPUT17), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n653), .B(new_n654), .C1(new_n445), .C2(new_n656), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n655), .A3(new_n653), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n625), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(G2096), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n665), .B(new_n666), .Z(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n672), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT20), .Z(new_n676));
  AOI211_X1 g251(.A(new_n674), .B(new_n676), .C1(new_n669), .C2(new_n673), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G32), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n466), .A2(G105), .ZN(new_n686));
  NAND3_X1  g261(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT26), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n475), .A2(G2105), .ZN(new_n689));
  INV_X1    g264(.A(G129), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI211_X1 g266(.A(new_n686), .B(new_n691), .C1(G141), .C2(new_n477), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n685), .B1(new_n692), .B2(new_n684), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT27), .B(G1996), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT25), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n698), .A2(new_n460), .ZN(new_n699));
  AOI211_X1 g274(.A(new_n697), .B(new_n699), .C1(G139), .C2(new_n477), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G29), .ZN(new_n701));
  NOR2_X1   g276(.A1(G29), .A2(G33), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT87), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(new_n443), .ZN(new_n705));
  INV_X1    g280(.A(G34), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(KEYINPUT24), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(KEYINPUT24), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(KEYINPUT88), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(KEYINPUT88), .B2(new_n708), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT89), .Z(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G29), .B2(G160), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n695), .B(new_n705), .C1(G2084), .C2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT96), .B(G1956), .Z(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G20), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT23), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n611), .B2(new_n716), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n714), .A2(KEYINPUT90), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n684), .A2(G35), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n684), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G2090), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n720), .B1(KEYINPUT95), .B2(new_n725), .C1(new_n715), .C2(new_n719), .ZN(new_n726));
  NOR2_X1   g301(.A1(G168), .A2(new_n716), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n716), .B2(G21), .ZN(new_n728));
  INV_X1    g303(.A(G1966), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G1348), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n605), .A2(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n716), .A2(G4), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n732), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n733), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n684), .A2(G27), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G164), .B2(new_n684), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT94), .B(G2078), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n725), .A2(KEYINPUT95), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n743), .B(new_n744), .C1(new_n714), .C2(KEYINPUT90), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n693), .A2(new_n694), .B1(new_n728), .B2(new_n729), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n684), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n477), .A2(G140), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n481), .A2(G128), .ZN(new_n750));
  OR2_X1    g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n751), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(new_n684), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n746), .B1(G2067), .B2(new_n755), .C1(G2084), .C2(new_n712), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT92), .B(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n758), .B2(KEYINPUT30), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(KEYINPUT93), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(KEYINPUT93), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(KEYINPUT30), .B2(new_n758), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n757), .B1(new_n760), .B2(new_n762), .C1(new_n632), .C2(new_n684), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G2067), .B2(new_n755), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n730), .B2(new_n731), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n756), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n716), .A2(G19), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n548), .B2(new_n716), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(G1341), .ZN(new_n769));
  NAND2_X1  g344(.A1(G301), .A2(G16), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n716), .A2(G5), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n768), .A2(G1341), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n772), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n775), .A2(G1961), .B1(new_n723), .B2(G2090), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n766), .A2(new_n769), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n726), .A2(new_n745), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n716), .A2(G24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n597), .B2(new_n716), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1986), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n481), .A2(G119), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n460), .A2(G107), .ZN(new_n783));
  OAI21_X1  g358(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G131), .B2(new_n477), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT85), .Z(new_n787));
  MUX2_X1   g362(.A(G25), .B(new_n787), .S(G29), .Z(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT35), .B(G1991), .Z(new_n790));
  AOI21_X1  g365(.A(new_n781), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n716), .A2(G22), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G166), .B2(new_n716), .ZN(new_n793));
  INV_X1    g368(.A(G1971), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n716), .A2(G6), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G305), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT32), .B(G1981), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n716), .A2(G23), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n575), .B2(new_n716), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n797), .A2(new_n799), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n795), .A2(new_n800), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n791), .B1(KEYINPUT34), .B2(new_n806), .C1(new_n789), .C2(new_n790), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(KEYINPUT34), .B2(new_n806), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT86), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n812));
  OR3_X1    g387(.A1(new_n808), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n778), .A2(new_n811), .A3(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  NAND2_X1  g390(.A1(new_n505), .A2(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n513), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n516), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n548), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n547), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n605), .A2(new_n615), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n825), .B(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n830));
  INV_X1    g405(.A(G860), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n821), .A2(new_n831), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(G145));
  XNOR2_X1  g411(.A(new_n692), .B(new_n700), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n481), .A2(G130), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n460), .A2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G142), .B2(new_n477), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(new_n622), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n837), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n492), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n491), .B1(new_n475), .B2(new_n488), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n495), .A2(new_n497), .ZN(new_n848));
  INV_X1    g423(.A(G126), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n689), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n753), .B(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n787), .B(new_n852), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n844), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n632), .B(KEYINPUT98), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n485), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G160), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT99), .Z(new_n860));
  AOI21_X1  g435(.A(G37), .B1(new_n855), .B2(new_n858), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g438(.A1(new_n823), .A2(new_n606), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n825), .B(KEYINPUT100), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n618), .ZN(new_n866));
  XNOR2_X1  g441(.A(G299), .B(new_n614), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n867), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n870), .B(KEYINPUT101), .C1(new_n871), .C2(new_n866), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(KEYINPUT101), .B2(new_n870), .ZN(new_n873));
  XNOR2_X1  g448(.A(G305), .B(G303), .ZN(new_n874));
  XNOR2_X1  g449(.A(G288), .B(new_n597), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n876), .A2(KEYINPUT102), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(KEYINPUT102), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n874), .B2(new_n877), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT103), .Z(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  MUX2_X1   g457(.A(new_n880), .B(new_n882), .S(KEYINPUT42), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n873), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n864), .B1(new_n884), .B2(new_n606), .ZN(G295));
  OAI21_X1  g460(.A(new_n864), .B1(new_n884), .B2(new_n606), .ZN(G331));
  OAI21_X1  g461(.A(G168), .B1(G301), .B2(KEYINPUT104), .ZN(new_n887));
  NAND2_X1  g462(.A1(G301), .A2(KEYINPUT104), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(new_n825), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n825), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n893), .A2(new_n867), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n894), .A2(new_n869), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(G37), .B1(new_n896), .B2(new_n881), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(new_n895), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n890), .A2(new_n893), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n871), .A2(KEYINPUT106), .A3(KEYINPUT41), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n899), .B(new_n900), .C1(new_n869), .C2(KEYINPUT106), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n898), .B1(new_n901), .B2(KEYINPUT107), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(KEYINPUT107), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n882), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n896), .A2(new_n881), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT43), .B1(new_n908), .B2(new_n897), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT44), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n906), .B1(new_n908), .B2(new_n897), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n913), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g489(.A(new_n473), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n468), .B(KEYINPUT67), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n915), .A2(G40), .A3(new_n463), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(G1384), .B1(new_n493), .B2(new_n498), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT45), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G1996), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n692), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT109), .ZN(new_n923));
  INV_X1    g498(.A(G2067), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n753), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n921), .B2(new_n692), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n790), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n787), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n754), .A2(new_n924), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n920), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n919), .A2(new_n921), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT125), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n920), .B1(new_n925), .B2(new_n692), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n934), .B2(new_n933), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n939), .B(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n787), .B(new_n790), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n942), .A2(KEYINPUT110), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(KEYINPUT110), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n919), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n927), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1986), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n597), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT108), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(new_n920), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT48), .Z(new_n952));
  AOI211_X1 g527(.A(new_n932), .B(new_n941), .C1(new_n947), .C2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT124), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n950), .B1(new_n948), .B2(new_n597), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n919), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n947), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1981), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n583), .C1(new_n589), .C2(new_n590), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n578), .A2(new_n582), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n527), .A2(G86), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n587), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(G1981), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n847), .B2(new_n850), .ZN(new_n968));
  OAI21_X1  g543(.A(G8), .B1(new_n968), .B2(new_n917), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G40), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n470), .A2(new_n473), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n918), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT113), .A3(G8), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n966), .A2(KEYINPUT49), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n964), .A2(new_n965), .A3(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1976), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n575), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n959), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n971), .A2(new_n975), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(G166), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n989));
  OAI22_X1  g564(.A1(G166), .A2(new_n985), .B1(KEYINPUT112), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n967), .B1(new_n499), .B2(new_n500), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n918), .A2(KEYINPUT45), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n917), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n992), .A2(new_n996), .A3(new_n993), .ZN(new_n999));
  AOI21_X1  g574(.A(G1971), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G2090), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n917), .B1(new_n918), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT68), .B1(new_n847), .B2(new_n850), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1001), .B(new_n1003), .C1(new_n1006), .C2(new_n1002), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(G8), .B(new_n991), .C1(new_n1000), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n575), .A2(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT113), .B1(new_n974), .B2(G8), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n970), .B(new_n985), .C1(new_n918), .C2(new_n973), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n976), .A2(new_n978), .B1(KEYINPUT52), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n980), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1010), .B(new_n1015), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n983), .A2(KEYINPUT114), .A3(new_n1010), .A4(new_n1015), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n984), .B1(new_n1009), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT63), .ZN(new_n1023));
  INV_X1    g598(.A(new_n991), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n973), .B1(new_n918), .B2(new_n1002), .ZN(new_n1025));
  AOI211_X1 g600(.A(G2090), .B(new_n1025), .C1(new_n1006), .C2(new_n1002), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n997), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n973), .A3(new_n999), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1026), .B1(new_n1028), .B2(new_n794), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1024), .B1(new_n1029), .B2(new_n985), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1030), .A2(new_n1009), .A3(new_n1020), .A4(new_n1014), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n973), .B1(new_n918), .B2(KEYINPUT45), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT116), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT45), .B(new_n967), .C1(new_n499), .C2(new_n500), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1036), .B(new_n973), .C1(new_n918), .C2(KEYINPUT45), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1032), .B1(new_n1038), .B2(G1966), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n973), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(KEYINPUT50), .B2(new_n992), .ZN(new_n1041));
  INV_X1    g616(.A(G2084), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT117), .A3(new_n729), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1039), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(G8), .A3(G168), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1023), .B1(new_n1031), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1047), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1008), .B1(new_n1028), .B2(new_n794), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1050), .A2(new_n985), .A3(new_n1024), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n1021), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1000), .B2(new_n1008), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1023), .B1(new_n1053), .B2(new_n1024), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1022), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G2078), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1003), .B1(new_n1006), .B2(new_n1002), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1038), .A2(new_n1058), .B1(new_n773), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1027), .A2(new_n444), .A3(new_n999), .A4(new_n973), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1057), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G171), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1031), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G168), .A2(new_n985), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1046), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1066), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(new_n1069), .B2(KEYINPUT122), .ZN(new_n1070));
  OAI211_X1 g645(.A(G8), .B(new_n1070), .C1(new_n1046), .C2(G286), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1045), .A2(new_n1043), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT117), .B1(new_n1044), .B2(new_n729), .ZN(new_n1073));
  OAI21_X1  g648(.A(G8), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1070), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1067), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1065), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g654(.A(KEYINPUT62), .B(new_n1067), .C1(new_n1076), .C2(new_n1071), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1056), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1067), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n995), .A2(new_n1058), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(new_n1033), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1059), .B2(new_n773), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1062), .A2(G301), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT54), .B1(new_n1064), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(new_n1031), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1060), .A2(new_n1062), .A3(G301), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1086), .A2(new_n1033), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1041), .B2(G1961), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1092), .B(KEYINPUT54), .C1(G301), .C2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1085), .A2(new_n1091), .A3(KEYINPUT123), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1062), .A2(G301), .A3(new_n1088), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1102), .A2(new_n1052), .A3(new_n1096), .A4(new_n1030), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1098), .B1(new_n1103), .B2(new_n1077), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT57), .B(new_n566), .C1(new_n557), .C2(new_n558), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n566), .A2(new_n555), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT119), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1105), .A2(KEYINPUT119), .A3(new_n1108), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1025), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1027), .A2(new_n973), .A3(new_n999), .A4(new_n1114), .ZN(new_n1115));
  AOI211_X1 g690(.A(new_n1109), .B(new_n1110), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1041), .A2(G1348), .B1(G2067), .B2(new_n974), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1117), .A2(new_n614), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1113), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1116), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT120), .B(G1996), .Z(new_n1122));
  INV_X1    g697(.A(new_n974), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT58), .B(G1341), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n1028), .A2(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n548), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1129));
  OR3_X1    g704(.A1(new_n1117), .A2(KEYINPUT60), .A3(new_n605), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1117), .A2(new_n614), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT60), .B1(new_n1118), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1115), .A2(new_n1113), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(new_n1119), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1120), .A2(KEYINPUT61), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1135), .A2(KEYINPUT61), .B1(new_n1116), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1121), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1097), .A2(new_n1104), .A3(new_n1138), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n954), .B(new_n957), .C1(new_n1082), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(new_n1142), .A3(new_n1065), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n1143), .A3(new_n1056), .ZN(new_n1144));
  INV_X1    g719(.A(new_n957), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT124), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n953), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT127), .B(new_n953), .C1(new_n1140), .C2(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g726(.A(G227), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n1153), .A2(G319), .ZN(new_n1154));
  NOR3_X1   g728(.A1(G229), .A2(G401), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n862), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g730(.A1(new_n913), .A2(new_n1156), .ZN(G308));
  OR2_X1    g731(.A1(new_n913), .A2(new_n1156), .ZN(G225));
endmodule


