

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759;

  XNOR2_X1 U370 ( .A(G146), .B(G125), .ZN(n466) );
  INV_X1 U371 ( .A(G128), .ZN(n405) );
  INV_X4 U372 ( .A(G953), .ZN(n752) );
  NAND2_X1 U373 ( .A1(n689), .A2(KEYINPUT76), .ZN(n369) );
  AND2_X2 U374 ( .A1(n751), .A2(n739), .ZN(n689) );
  XNOR2_X1 U375 ( .A(n459), .B(KEYINPUT71), .ZN(n527) );
  XOR2_X1 U376 ( .A(n594), .B(KEYINPUT80), .Z(n348) );
  XNOR2_X2 U377 ( .A(n589), .B(KEYINPUT35), .ZN(n637) );
  XNOR2_X2 U378 ( .A(n501), .B(n407), .ZN(n750) );
  AND2_X1 U379 ( .A1(n651), .A2(n650), .ZN(n653) );
  INV_X1 U380 ( .A(n532), .ZN(n671) );
  OR2_X2 U381 ( .A1(n620), .A2(G902), .ZN(n427) );
  AND2_X2 U382 ( .A1(n616), .A2(n615), .ZN(n654) );
  NAND2_X1 U383 ( .A1(n367), .A2(n365), .ZN(n616) );
  NAND2_X1 U384 ( .A1(n356), .A2(n366), .ZN(n365) );
  NAND2_X1 U385 ( .A1(n399), .A2(n398), .ZN(n612) );
  AND2_X1 U386 ( .A1(n526), .A2(n693), .ZN(n685) );
  XNOR2_X1 U387 ( .A(n574), .B(KEYINPUT32), .ZN(n636) );
  OR2_X1 U388 ( .A1(n582), .A2(n592), .ZN(n584) );
  XNOR2_X1 U389 ( .A(n602), .B(n388), .ZN(n592) );
  BUF_X1 U390 ( .A(n501), .Z(n502) );
  BUF_X1 U391 ( .A(n654), .Z(n644) );
  XNOR2_X2 U392 ( .A(n464), .B(G134), .ZN(n501) );
  XNOR2_X2 U393 ( .A(n426), .B(n413), .ZN(n638) );
  XNOR2_X1 U394 ( .A(n685), .B(KEYINPUT79), .ZN(n364) );
  NAND2_X1 U395 ( .A1(KEYINPUT44), .A2(KEYINPUT64), .ZN(n397) );
  AND2_X1 U396 ( .A1(n634), .A2(n608), .ZN(n393) );
  NAND2_X1 U397 ( .A1(n372), .A2(n420), .ZN(n371) );
  NOR2_X1 U398 ( .A1(n677), .A2(n362), .ZN(n555) );
  NAND2_X1 U399 ( .A1(n387), .A2(n349), .ZN(n362) );
  NAND2_X1 U400 ( .A1(n382), .A2(n504), .ZN(n381) );
  AND2_X1 U401 ( .A1(n550), .A2(n629), .ZN(n363) );
  NAND2_X1 U402 ( .A1(n400), .A2(n591), .ZN(n399) );
  NAND2_X1 U403 ( .A1(n393), .A2(n392), .ZN(n391) );
  AND2_X1 U404 ( .A1(n634), .A2(n389), .ZN(n395) );
  INV_X1 U405 ( .A(KEYINPUT101), .ZN(n416) );
  XNOR2_X1 U406 ( .A(n490), .B(n489), .ZN(n648) );
  XNOR2_X1 U407 ( .A(n571), .B(n355), .ZN(n573) );
  AND2_X1 U408 ( .A1(n573), .A2(n575), .ZN(n593) );
  INV_X1 U409 ( .A(KEYINPUT6), .ZN(n388) );
  NOR2_X1 U410 ( .A1(n390), .A2(n396), .ZN(n389) );
  INV_X1 U411 ( .A(KEYINPUT64), .ZN(n396) );
  XNOR2_X1 U412 ( .A(KEYINPUT65), .B(G101), .ZN(n465) );
  XNOR2_X1 U413 ( .A(G113), .B(G143), .ZN(n358) );
  AND2_X1 U414 ( .A1(n739), .A2(n377), .ZN(n357) );
  INV_X1 U415 ( .A(KEYINPUT76), .ZN(n366) );
  XNOR2_X1 U416 ( .A(n465), .B(n466), .ZN(n378) );
  OR2_X2 U417 ( .A1(n383), .A2(n380), .ZN(n596) );
  NAND2_X1 U418 ( .A1(n385), .A2(n384), .ZN(n383) );
  AND2_X1 U419 ( .A1(n353), .A2(n374), .ZN(n373) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n539) );
  XNOR2_X1 U421 ( .A(n491), .B(G475), .ZN(n359) );
  OR2_X1 U422 ( .A1(n648), .A2(G902), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n524), .ZN(n526) );
  NAND2_X1 U424 ( .A1(n555), .A2(n529), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n402), .B(KEYINPUT72), .ZN(n401) );
  NOR2_X1 U426 ( .A1(n572), .A2(n352), .ZN(n402) );
  NAND2_X1 U427 ( .A1(n348), .A2(n696), .ZN(n634) );
  AND2_X1 U428 ( .A1(n595), .A2(n350), .ZN(n349) );
  AND2_X1 U429 ( .A1(n522), .A2(n707), .ZN(n350) );
  NAND2_X1 U430 ( .A1(n580), .A2(n579), .ZN(n351) );
  NAND2_X1 U431 ( .A1(n693), .A2(n595), .ZN(n352) );
  AND2_X1 U432 ( .A1(n525), .A2(n458), .ZN(n353) );
  AND2_X1 U433 ( .A1(n364), .A2(n363), .ZN(n354) );
  XOR2_X1 U434 ( .A(KEYINPUT68), .B(KEYINPUT22), .Z(n355) );
  INV_X1 U435 ( .A(n614), .ZN(n377) );
  NOR2_X1 U436 ( .A1(n752), .A2(G952), .ZN(n659) );
  NAND2_X1 U437 ( .A1(n357), .A2(n751), .ZN(n356) );
  XNOR2_X1 U438 ( .A(n358), .B(G122), .ZN(n484) );
  NAND2_X1 U439 ( .A1(n368), .A2(n377), .ZN(n367) );
  NAND2_X1 U440 ( .A1(n369), .A2(n613), .ZN(n368) );
  NAND2_X1 U441 ( .A1(n371), .A2(n370), .ZN(n375) );
  NAND2_X1 U442 ( .A1(n576), .A2(n376), .ZN(n370) );
  INV_X1 U443 ( .A(n576), .ZN(n372) );
  NAND2_X1 U444 ( .A1(n375), .A2(n373), .ZN(n459) );
  NAND2_X1 U445 ( .A1(n419), .A2(n534), .ZN(n374) );
  NAND2_X1 U446 ( .A1(n420), .A2(n707), .ZN(n376) );
  XNOR2_X2 U447 ( .A(n596), .B(n416), .ZN(n576) );
  AND2_X1 U448 ( .A1(n689), .A2(KEYINPUT2), .ZN(n690) );
  XNOR2_X1 U449 ( .A(n464), .B(n378), .ZN(n473) );
  XNOR2_X2 U450 ( .A(n379), .B(n405), .ZN(n464) );
  XNOR2_X2 U451 ( .A(G143), .B(KEYINPUT74), .ZN(n379) );
  NAND2_X1 U452 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U453 ( .A1(n394), .A2(n391), .ZN(n398) );
  XNOR2_X2 U454 ( .A(n410), .B(n409), .ZN(n461) );
  NOR2_X1 U455 ( .A1(n638), .A2(n381), .ZN(n380) );
  INV_X1 U456 ( .A(n415), .ZN(n382) );
  NAND2_X1 U457 ( .A1(n415), .A2(G902), .ZN(n384) );
  NAND2_X1 U458 ( .A1(n638), .A2(n415), .ZN(n385) );
  INV_X1 U459 ( .A(n508), .ZN(n554) );
  XNOR2_X2 U460 ( .A(n386), .B(KEYINPUT39), .ZN(n508) );
  NAND2_X1 U461 ( .A1(n527), .A2(n706), .ZN(n386) );
  INV_X1 U462 ( .A(n592), .ZN(n387) );
  INV_X1 U463 ( .A(n608), .ZN(n390) );
  NAND2_X1 U464 ( .A1(n609), .A2(n397), .ZN(n392) );
  NAND2_X1 U465 ( .A1(n395), .A2(n637), .ZN(n394) );
  NAND2_X1 U466 ( .A1(n351), .A2(n590), .ZN(n400) );
  NAND2_X1 U467 ( .A1(n573), .A2(n401), .ZN(n574) );
  AND2_X1 U468 ( .A1(n619), .A2(n650), .ZN(G63) );
  XNOR2_X1 U469 ( .A(KEYINPUT59), .B(n648), .ZN(n404) );
  INV_X1 U470 ( .A(KEYINPUT46), .ZN(n520) );
  XNOR2_X1 U471 ( .A(n521), .B(n520), .ZN(n551) );
  INV_X1 U472 ( .A(KEYINPUT2), .ZN(n613) );
  INV_X1 U473 ( .A(n690), .ZN(n615) );
  XNOR2_X1 U474 ( .A(n477), .B(n476), .ZN(n533) );
  BUF_X1 U475 ( .A(n533), .Z(n558) );
  NAND2_X1 U476 ( .A1(n593), .A2(n577), .ZN(n630) );
  XNOR2_X1 U477 ( .A(KEYINPUT66), .B(G131), .ZN(n479) );
  XNOR2_X1 U478 ( .A(KEYINPUT4), .B(G137), .ZN(n406) );
  XNOR2_X1 U479 ( .A(n479), .B(n406), .ZN(n407) );
  XNOR2_X1 U480 ( .A(n465), .B(G146), .ZN(n408) );
  XNOR2_X2 U481 ( .A(n750), .B(n408), .ZN(n426) );
  XNOR2_X2 U482 ( .A(G116), .B(G113), .ZN(n410) );
  XNOR2_X2 U483 ( .A(KEYINPUT3), .B(G119), .ZN(n409) );
  NOR2_X1 U484 ( .A1(G953), .A2(G237), .ZN(n482) );
  NAND2_X1 U485 ( .A1(n482), .A2(G210), .ZN(n411) );
  XNOR2_X1 U486 ( .A(n411), .B(KEYINPUT5), .ZN(n412) );
  XNOR2_X1 U487 ( .A(n461), .B(n412), .ZN(n413) );
  INV_X1 U488 ( .A(KEYINPUT91), .ZN(n414) );
  XNOR2_X1 U489 ( .A(n414), .B(G472), .ZN(n415) );
  INV_X1 U490 ( .A(G902), .ZN(n504) );
  INV_X1 U491 ( .A(G237), .ZN(n417) );
  NAND2_X1 U492 ( .A1(n504), .A2(n417), .ZN(n475) );
  NAND2_X1 U493 ( .A1(n475), .A2(G214), .ZN(n707) );
  INV_X1 U494 ( .A(KEYINPUT105), .ZN(n418) );
  XNOR2_X1 U495 ( .A(n418), .B(KEYINPUT30), .ZN(n419) );
  INV_X1 U496 ( .A(n419), .ZN(n420) );
  XNOR2_X1 U497 ( .A(G107), .B(G104), .ZN(n421) );
  XNOR2_X1 U498 ( .A(n421), .B(G110), .ZN(n463) );
  XOR2_X1 U499 ( .A(KEYINPUT86), .B(G140), .Z(n423) );
  NAND2_X1 U500 ( .A1(n752), .A2(G227), .ZN(n422) );
  XNOR2_X1 U501 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U502 ( .A(n463), .B(n424), .ZN(n425) );
  XNOR2_X1 U503 ( .A(n426), .B(n425), .ZN(n620) );
  XNOR2_X2 U504 ( .A(n427), .B(G469), .ZN(n525) );
  XNOR2_X1 U505 ( .A(KEYINPUT75), .B(KEYINPUT8), .ZN(n429) );
  NAND2_X1 U506 ( .A1(G234), .A2(n752), .ZN(n428) );
  XNOR2_X1 U507 ( .A(n429), .B(n428), .ZN(n498) );
  NAND2_X1 U508 ( .A1(n498), .A2(G221), .ZN(n434) );
  XNOR2_X1 U509 ( .A(G119), .B(G128), .ZN(n430) );
  XNOR2_X1 U510 ( .A(n430), .B(KEYINPUT67), .ZN(n432) );
  XNOR2_X1 U511 ( .A(KEYINPUT88), .B(KEYINPUT23), .ZN(n431) );
  XNOR2_X1 U512 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U513 ( .A(n434), .B(n433), .ZN(n440) );
  XNOR2_X1 U514 ( .A(KEYINPUT10), .B(G140), .ZN(n435) );
  XNOR2_X1 U515 ( .A(n466), .B(n435), .ZN(n748) );
  XNOR2_X1 U516 ( .A(G137), .B(KEYINPUT24), .ZN(n437) );
  XNOR2_X1 U517 ( .A(G110), .B(KEYINPUT87), .ZN(n436) );
  XNOR2_X1 U518 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U519 ( .A(n748), .B(n438), .ZN(n439) );
  XNOR2_X1 U520 ( .A(n440), .B(n439), .ZN(n645) );
  OR2_X1 U521 ( .A1(n645), .A2(G902), .ZN(n444) );
  XNOR2_X1 U522 ( .A(G902), .B(KEYINPUT15), .ZN(n614) );
  NAND2_X1 U523 ( .A1(n614), .A2(G234), .ZN(n441) );
  XNOR2_X1 U524 ( .A(n441), .B(KEYINPUT20), .ZN(n445) );
  AND2_X1 U525 ( .A1(n445), .A2(G217), .ZN(n442) );
  XNOR2_X1 U526 ( .A(n442), .B(KEYINPUT25), .ZN(n443) );
  XNOR2_X1 U527 ( .A(n444), .B(n443), .ZN(n696) );
  INV_X1 U528 ( .A(n445), .ZN(n447) );
  INV_X1 U529 ( .A(G221), .ZN(n446) );
  OR2_X1 U530 ( .A1(n447), .A2(n446), .ZN(n451) );
  XOR2_X1 U531 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n449) );
  INV_X1 U532 ( .A(KEYINPUT89), .ZN(n448) );
  XNOR2_X1 U533 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U534 ( .A(n451), .B(n450), .ZN(n695) );
  NAND2_X1 U535 ( .A1(G234), .A2(G237), .ZN(n452) );
  XNOR2_X1 U536 ( .A(n452), .B(KEYINPUT14), .ZN(n722) );
  OR2_X1 U537 ( .A1(n752), .A2(G902), .ZN(n453) );
  AND2_X1 U538 ( .A1(n722), .A2(n453), .ZN(n565) );
  INV_X1 U539 ( .A(G952), .ZN(n454) );
  NAND2_X1 U540 ( .A1(n752), .A2(n454), .ZN(n563) );
  NAND2_X1 U541 ( .A1(G953), .A2(G900), .ZN(n455) );
  AND2_X1 U542 ( .A1(n563), .A2(n455), .ZN(n456) );
  AND2_X1 U543 ( .A1(n565), .A2(n456), .ZN(n457) );
  AND2_X1 U544 ( .A1(n695), .A2(n457), .ZN(n522) );
  AND2_X1 U545 ( .A1(n696), .A2(n522), .ZN(n458) );
  XNOR2_X1 U546 ( .A(KEYINPUT16), .B(G122), .ZN(n460) );
  XNOR2_X1 U547 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U548 ( .A(n463), .B(n462), .ZN(n736) );
  XNOR2_X1 U549 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n468) );
  XNOR2_X1 U550 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n467) );
  XNOR2_X1 U551 ( .A(n468), .B(n467), .ZN(n471) );
  NAND2_X1 U552 ( .A1(n752), .A2(G224), .ZN(n469) );
  XNOR2_X1 U553 ( .A(n469), .B(KEYINPUT83), .ZN(n470) );
  XNOR2_X1 U554 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U555 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U556 ( .A(n736), .B(n474), .ZN(n656) );
  NAND2_X1 U557 ( .A1(n656), .A2(n614), .ZN(n477) );
  NAND2_X1 U558 ( .A1(n475), .A2(G210), .ZN(n476) );
  XNOR2_X1 U559 ( .A(KEYINPUT70), .B(KEYINPUT38), .ZN(n478) );
  XNOR2_X1 U560 ( .A(n558), .B(n478), .ZN(n706) );
  XOR2_X1 U561 ( .A(KEYINPUT94), .B(G104), .Z(n480) );
  XNOR2_X1 U562 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U563 ( .A(n481), .B(n748), .ZN(n490) );
  AND2_X1 U564 ( .A1(n482), .A2(G214), .ZN(n483) );
  XNOR2_X1 U565 ( .A(n484), .B(n483), .ZN(n488) );
  XOR2_X1 U566 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n486) );
  XNOR2_X1 U567 ( .A(KEYINPUT93), .B(KEYINPUT95), .ZN(n485) );
  XNOR2_X1 U568 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U569 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U570 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n491) );
  XOR2_X1 U571 ( .A(KEYINPUT98), .B(G107), .Z(n493) );
  XNOR2_X1 U572 ( .A(G116), .B(G122), .ZN(n492) );
  XNOR2_X1 U573 ( .A(n493), .B(n492), .ZN(n497) );
  XOR2_X1 U574 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n495) );
  XNOR2_X1 U575 ( .A(KEYINPUT97), .B(KEYINPUT99), .ZN(n494) );
  XNOR2_X1 U576 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U577 ( .A(n497), .B(n496), .ZN(n500) );
  NAND2_X1 U578 ( .A1(n498), .A2(G217), .ZN(n499) );
  XNOR2_X1 U579 ( .A(n500), .B(n499), .ZN(n503) );
  XNOR2_X1 U580 ( .A(n503), .B(n502), .ZN(n617) );
  NAND2_X1 U581 ( .A1(n617), .A2(n504), .ZN(n506) );
  INV_X1 U582 ( .A(G478), .ZN(n505) );
  XNOR2_X1 U583 ( .A(n506), .B(n505), .ZN(n515) );
  INV_X1 U584 ( .A(n515), .ZN(n538) );
  OR2_X1 U585 ( .A1(n539), .A2(n538), .ZN(n541) );
  INV_X1 U586 ( .A(n541), .ZN(n507) );
  NAND2_X2 U587 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X2 U588 ( .A(n509), .B(KEYINPUT40), .ZN(n635) );
  INV_X1 U589 ( .A(n522), .ZN(n510) );
  NOR2_X1 U590 ( .A1(n696), .A2(n510), .ZN(n511) );
  NAND2_X1 U591 ( .A1(n576), .A2(n511), .ZN(n512) );
  XNOR2_X1 U592 ( .A(n512), .B(KEYINPUT28), .ZN(n514) );
  INV_X1 U593 ( .A(n525), .ZN(n513) );
  OR2_X1 U594 ( .A1(n514), .A2(n513), .ZN(n532) );
  NAND2_X1 U595 ( .A1(n706), .A2(n707), .ZN(n711) );
  NAND2_X1 U596 ( .A1(n539), .A2(n515), .ZN(n710) );
  OR2_X1 U597 ( .A1(n711), .A2(n710), .ZN(n518) );
  INV_X1 U598 ( .A(KEYINPUT106), .ZN(n516) );
  XNOR2_X1 U599 ( .A(n516), .B(KEYINPUT41), .ZN(n517) );
  XNOR2_X1 U600 ( .A(n518), .B(n517), .ZN(n726) );
  OR2_X1 U601 ( .A1(n532), .A2(n726), .ZN(n519) );
  XNOR2_X1 U602 ( .A(n519), .B(KEYINPUT42), .ZN(n631) );
  NAND2_X1 U603 ( .A1(n635), .A2(n631), .ZN(n521) );
  XOR2_X1 U604 ( .A(KEYINPUT103), .B(n541), .Z(n677) );
  INV_X1 U605 ( .A(n696), .ZN(n595) );
  INV_X1 U606 ( .A(n596), .ZN(n602) );
  INV_X1 U607 ( .A(n558), .ZN(n529) );
  XOR2_X1 U608 ( .A(KEYINPUT107), .B(KEYINPUT36), .Z(n523) );
  XNOR2_X1 U609 ( .A(n523), .B(KEYINPUT81), .ZN(n524) );
  XNOR2_X2 U610 ( .A(n525), .B(KEYINPUT1), .ZN(n693) );
  INV_X1 U611 ( .A(n527), .ZN(n531) );
  INV_X1 U612 ( .A(n539), .ZN(n528) );
  AND2_X1 U613 ( .A1(n528), .A2(n538), .ZN(n587) );
  NAND2_X1 U614 ( .A1(n587), .A2(n529), .ZN(n530) );
  OR2_X1 U615 ( .A1(n531), .A2(n530), .ZN(n629) );
  INV_X1 U616 ( .A(n533), .ZN(n535) );
  INV_X1 U617 ( .A(n707), .ZN(n534) );
  NAND2_X1 U618 ( .A1(n535), .A2(n707), .ZN(n537) );
  INV_X1 U619 ( .A(KEYINPUT19), .ZN(n536) );
  XNOR2_X2 U620 ( .A(n537), .B(n536), .ZN(n669) );
  NAND2_X1 U621 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U622 ( .A(n540), .B(KEYINPUT100), .ZN(n682) );
  AND2_X1 U623 ( .A1(n682), .A2(n541), .ZN(n712) );
  OR2_X1 U624 ( .A1(n712), .A2(KEYINPUT69), .ZN(n542) );
  NOR2_X1 U625 ( .A1(n669), .A2(n542), .ZN(n543) );
  NAND2_X1 U626 ( .A1(n671), .A2(n543), .ZN(n545) );
  INV_X1 U627 ( .A(KEYINPUT47), .ZN(n544) );
  XNOR2_X1 U628 ( .A(n545), .B(n544), .ZN(n549) );
  NAND2_X1 U629 ( .A1(n712), .A2(KEYINPUT69), .ZN(n546) );
  NOR2_X1 U630 ( .A1(n546), .A2(n669), .ZN(n547) );
  NAND2_X1 U631 ( .A1(n547), .A2(n671), .ZN(n548) );
  AND2_X1 U632 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U633 ( .A1(n551), .A2(n354), .ZN(n553) );
  INV_X1 U634 ( .A(KEYINPUT48), .ZN(n552) );
  XNOR2_X1 U635 ( .A(n553), .B(n552), .ZN(n561) );
  OR2_X1 U636 ( .A1(n554), .A2(n682), .ZN(n687) );
  XNOR2_X1 U637 ( .A(n555), .B(KEYINPUT104), .ZN(n556) );
  INV_X1 U638 ( .A(n693), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n556), .A2(n575), .ZN(n557) );
  XNOR2_X1 U640 ( .A(n557), .B(KEYINPUT43), .ZN(n559) );
  NAND2_X1 U641 ( .A1(n559), .A2(n558), .ZN(n632) );
  AND2_X1 U642 ( .A1(n687), .A2(n632), .ZN(n560) );
  AND2_X2 U643 ( .A1(n561), .A2(n560), .ZN(n751) );
  NAND2_X1 U644 ( .A1(G953), .A2(G898), .ZN(n562) );
  AND2_X1 U645 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U646 ( .A1(n565), .A2(n564), .ZN(n566) );
  OR2_X2 U647 ( .A1(n669), .A2(n566), .ZN(n568) );
  INV_X1 U648 ( .A(KEYINPUT0), .ZN(n567) );
  XNOR2_X2 U649 ( .A(n568), .B(n567), .ZN(n598) );
  INV_X1 U650 ( .A(n695), .ZN(n569) );
  NOR2_X1 U651 ( .A1(n710), .A2(n569), .ZN(n570) );
  NAND2_X1 U652 ( .A1(n598), .A2(n570), .ZN(n571) );
  XNOR2_X1 U653 ( .A(n592), .B(KEYINPUT73), .ZN(n572) );
  AND2_X1 U654 ( .A1(n372), .A2(n595), .ZN(n577) );
  NAND2_X1 U655 ( .A1(n636), .A2(n630), .ZN(n580) );
  INV_X1 U656 ( .A(KEYINPUT44), .ZN(n578) );
  OR2_X1 U657 ( .A1(n578), .A2(KEYINPUT64), .ZN(n579) );
  INV_X1 U658 ( .A(n598), .ZN(n581) );
  XNOR2_X1 U659 ( .A(n581), .B(KEYINPUT85), .ZN(n601) );
  AND2_X1 U660 ( .A1(n696), .A2(n695), .ZN(n692) );
  NAND2_X1 U661 ( .A1(n693), .A2(n692), .ZN(n582) );
  XNOR2_X1 U662 ( .A(KEYINPUT102), .B(KEYINPUT33), .ZN(n583) );
  XNOR2_X2 U663 ( .A(n584), .B(n583), .ZN(n728) );
  NAND2_X1 U664 ( .A1(n601), .A2(n728), .ZN(n586) );
  INV_X1 U665 ( .A(KEYINPUT34), .ZN(n585) );
  XNOR2_X1 U666 ( .A(n586), .B(n585), .ZN(n588) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n589) );
  INV_X1 U668 ( .A(n637), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n578), .A2(KEYINPUT64), .ZN(n591) );
  AND2_X1 U670 ( .A1(n596), .A2(n692), .ZN(n597) );
  AND2_X1 U671 ( .A1(n693), .A2(n597), .ZN(n702) );
  NAND2_X1 U672 ( .A1(n598), .A2(n702), .ZN(n600) );
  XOR2_X1 U673 ( .A(KEYINPUT92), .B(KEYINPUT31), .Z(n599) );
  XNOR2_X1 U674 ( .A(n600), .B(n599), .ZN(n681) );
  INV_X1 U675 ( .A(n601), .ZN(n605) );
  AND2_X1 U676 ( .A1(n525), .A2(n692), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  OR2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n665) );
  NAND2_X1 U679 ( .A1(n681), .A2(n665), .ZN(n607) );
  INV_X1 U680 ( .A(n712), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n608) );
  AND2_X1 U682 ( .A1(n630), .A2(n636), .ZN(n609) );
  INV_X1 U683 ( .A(KEYINPUT77), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT45), .ZN(n611) );
  XNOR2_X2 U685 ( .A(n612), .B(n611), .ZN(n739) );
  NAND2_X1 U686 ( .A1(n644), .A2(G478), .ZN(n618) );
  XNOR2_X1 U687 ( .A(n618), .B(n617), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n654), .A2(G469), .ZN(n624) );
  XOR2_X1 U689 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n621) );
  XNOR2_X1 U690 ( .A(n621), .B(KEYINPUT58), .ZN(n622) );
  XNOR2_X1 U691 ( .A(n620), .B(n622), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n624), .B(n623), .ZN(n625) );
  NOR2_X2 U693 ( .A1(n625), .A2(n659), .ZN(n627) );
  INV_X1 U694 ( .A(KEYINPUT123), .ZN(n626) );
  XNOR2_X1 U695 ( .A(n627), .B(n626), .ZN(G54) );
  XOR2_X1 U696 ( .A(G143), .B(KEYINPUT111), .Z(n628) );
  XNOR2_X1 U697 ( .A(n629), .B(n628), .ZN(G45) );
  XNOR2_X1 U698 ( .A(n630), .B(G110), .ZN(G12) );
  XNOR2_X1 U699 ( .A(n631), .B(G137), .ZN(G39) );
  XNOR2_X1 U700 ( .A(n632), .B(G140), .ZN(G42) );
  XNOR2_X1 U701 ( .A(G101), .B(KEYINPUT108), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(G3) );
  XNOR2_X1 U703 ( .A(n635), .B(G131), .ZN(G33) );
  XNOR2_X1 U704 ( .A(n636), .B(G119), .ZN(G21) );
  XOR2_X1 U705 ( .A(n637), .B(G122), .Z(G24) );
  NAND2_X1 U706 ( .A1(n654), .A2(G472), .ZN(n640) );
  XNOR2_X1 U707 ( .A(n638), .B(KEYINPUT62), .ZN(n639) );
  XNOR2_X1 U708 ( .A(n640), .B(n639), .ZN(n641) );
  NOR2_X2 U709 ( .A1(n641), .A2(n659), .ZN(n643) );
  XOR2_X1 U710 ( .A(KEYINPUT82), .B(KEYINPUT63), .Z(n642) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(G57) );
  NAND2_X1 U712 ( .A1(n644), .A2(G217), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X1 U714 ( .A1(n647), .A2(n659), .ZN(G66) );
  NAND2_X1 U715 ( .A1(n654), .A2(G475), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n649), .B(n404), .ZN(n651) );
  INV_X1 U717 ( .A(n659), .ZN(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n652) );
  XNOR2_X1 U719 ( .A(n653), .B(n652), .ZN(G60) );
  NAND2_X1 U720 ( .A1(n654), .A2(G210), .ZN(n658) );
  XNOR2_X1 U721 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n655) );
  XNOR2_X1 U722 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U723 ( .A(n658), .B(n657), .ZN(n660) );
  NOR2_X2 U724 ( .A1(n660), .A2(n659), .ZN(n662) );
  XNOR2_X1 U725 ( .A(KEYINPUT78), .B(KEYINPUT56), .ZN(n661) );
  XNOR2_X1 U726 ( .A(n662), .B(n661), .ZN(G51) );
  NOR2_X1 U727 ( .A1(n665), .A2(n677), .ZN(n664) );
  XNOR2_X1 U728 ( .A(G104), .B(KEYINPUT109), .ZN(n663) );
  XNOR2_X1 U729 ( .A(n664), .B(n663), .ZN(G6) );
  NOR2_X1 U730 ( .A1(n665), .A2(n682), .ZN(n667) );
  XNOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n666) );
  XNOR2_X1 U732 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U733 ( .A(G107), .B(n668), .ZN(G9) );
  XOR2_X1 U734 ( .A(KEYINPUT29), .B(KEYINPUT110), .Z(n673) );
  INV_X1 U735 ( .A(n669), .ZN(n670) );
  NAND2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n675) );
  OR2_X1 U737 ( .A1(n675), .A2(n682), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U739 ( .A(G128), .B(n674), .ZN(G30) );
  NOR2_X1 U740 ( .A1(n675), .A2(n677), .ZN(n676) );
  XOR2_X1 U741 ( .A(G146), .B(n676), .Z(G48) );
  NOR2_X1 U742 ( .A1(n681), .A2(n677), .ZN(n679) );
  XNOR2_X1 U743 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n678) );
  XNOR2_X1 U744 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U745 ( .A(G113), .B(n680), .ZN(G15) );
  NOR2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U747 ( .A(KEYINPUT114), .B(n683), .Z(n684) );
  XNOR2_X1 U748 ( .A(G116), .B(n684), .ZN(G18) );
  XNOR2_X1 U749 ( .A(G125), .B(n685), .ZN(n686) );
  XNOR2_X1 U750 ( .A(n686), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U751 ( .A(G134), .B(n687), .Z(n688) );
  XNOR2_X1 U752 ( .A(n688), .B(KEYINPUT115), .ZN(G36) );
  XOR2_X1 U753 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n735) );
  NOR2_X1 U754 ( .A1(n689), .A2(KEYINPUT2), .ZN(n691) );
  NOR2_X1 U755 ( .A1(n691), .A2(n690), .ZN(n732) );
  NOR2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U757 ( .A(n694), .B(KEYINPUT50), .ZN(n700) );
  NOR2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U759 ( .A(n697), .B(KEYINPUT49), .ZN(n698) );
  NAND2_X1 U760 ( .A1(n602), .A2(n698), .ZN(n699) );
  NOR2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U762 ( .A(n701), .B(KEYINPUT116), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U764 ( .A(KEYINPUT51), .B(n704), .Z(n705) );
  NOR2_X1 U765 ( .A1(n726), .A2(n705), .ZN(n720) );
  NOR2_X1 U766 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U767 ( .A(KEYINPUT117), .B(n708), .Z(n709) );
  NOR2_X1 U768 ( .A1(n710), .A2(n709), .ZN(n715) );
  NOR2_X1 U769 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U770 ( .A(n713), .B(KEYINPUT118), .ZN(n714) );
  NOR2_X1 U771 ( .A1(n715), .A2(n714), .ZN(n717) );
  INV_X1 U772 ( .A(n728), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U774 ( .A(KEYINPUT119), .B(n718), .Z(n719) );
  NOR2_X1 U775 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U776 ( .A(KEYINPUT52), .B(n721), .ZN(n724) );
  NAND2_X1 U777 ( .A1(G952), .A2(n722), .ZN(n723) );
  NOR2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U779 ( .A1(G953), .A2(n725), .ZN(n730) );
  INV_X1 U780 ( .A(n726), .ZN(n727) );
  NAND2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n733), .B(KEYINPUT120), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n735), .B(n734), .ZN(G75) );
  XNOR2_X1 U786 ( .A(n736), .B(G101), .ZN(n738) );
  NOR2_X1 U787 ( .A1(n752), .A2(G898), .ZN(n737) );
  NOR2_X1 U788 ( .A1(n738), .A2(n737), .ZN(n747) );
  AND2_X1 U789 ( .A1(n739), .A2(n752), .ZN(n745) );
  INV_X1 U790 ( .A(G898), .ZN(n743) );
  NAND2_X1 U791 ( .A1(G224), .A2(G953), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n740), .B(KEYINPUT125), .ZN(n741) );
  XNOR2_X1 U793 ( .A(n741), .B(KEYINPUT61), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U795 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U796 ( .A(n747), .B(n746), .Z(G69) );
  XNOR2_X1 U797 ( .A(n748), .B(KEYINPUT126), .ZN(n749) );
  XNOR2_X1 U798 ( .A(n750), .B(n749), .ZN(n754) );
  XOR2_X1 U799 ( .A(n754), .B(n751), .Z(n753) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n759) );
  XNOR2_X1 U801 ( .A(G227), .B(n754), .ZN(n755) );
  NAND2_X1 U802 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U803 ( .A1(G953), .A2(n756), .ZN(n757) );
  XOR2_X1 U804 ( .A(KEYINPUT127), .B(n757), .Z(n758) );
  NAND2_X1 U805 ( .A1(n759), .A2(n758), .ZN(G72) );
endmodule

