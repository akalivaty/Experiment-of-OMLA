//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  NAND2_X1  g0021(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n219), .A2(new_n221), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(new_n209), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n212), .B1(new_n214), .B2(new_n215), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G68), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT67), .B(G50), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G1), .A2(G13), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n207), .A2(new_n249), .A3(KEYINPUT71), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT71), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G20), .B2(G33), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G50), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n207), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n256), .A2(new_n257), .B1(new_n207), .B2(G68), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n248), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT11), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT73), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT72), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n206), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n261), .B1(new_n266), .B2(new_n248), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n265), .ZN(new_n268));
  INV_X1    g0068(.A(new_n248), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(KEYINPUT73), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(G68), .C1(G1), .C2(new_n207), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT12), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n266), .B2(new_n202), .ZN(new_n274));
  INV_X1    g0074(.A(G13), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G1), .ZN(new_n276));
  AND4_X1   g0076(.A1(new_n273), .A2(new_n276), .A3(G20), .A4(new_n202), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n260), .B(new_n272), .C1(new_n274), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G226), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n230), .A2(G1698), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G97), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n285), .A2(KEYINPUT75), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT75), .B1(new_n285), .B2(new_n286), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G1), .A3(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT68), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT68), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n294), .B(new_n206), .C1(G41), .C2(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n213), .B2(new_n289), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G238), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT69), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n206), .B(KEYINPUT69), .C1(G41), .C2(G45), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n290), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n299), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT13), .B1(new_n291), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n302), .A2(new_n290), .A3(new_n303), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(G238), .B1(new_n298), .B2(new_n296), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT13), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n247), .B1(G33), .B2(G41), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n281), .A2(new_n282), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT3), .B(G33), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n311), .A2(new_n312), .B1(G33), .B2(G97), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n310), .B1(new_n313), .B2(KEYINPUT75), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n308), .B(new_n309), .C1(new_n314), .C2(new_n287), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n306), .A2(KEYINPUT76), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  INV_X1    g0117(.A(new_n291), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT76), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(new_n309), .A4(new_n308), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n316), .A2(new_n317), .A3(G169), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT77), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n316), .A2(G169), .A3(new_n320), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT14), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n306), .A2(G179), .A3(new_n315), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n321), .A2(KEYINPUT77), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n278), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n315), .A2(G190), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n278), .B1(new_n306), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n316), .A2(G200), .A3(new_n320), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G150), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n253), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT8), .B(G58), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n256), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n248), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n262), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n248), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n254), .B1(new_n206), .B2(G20), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n340), .A2(new_n341), .B1(new_n254), .B2(new_n339), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT9), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n338), .A2(KEYINPUT9), .A3(new_n342), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT74), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT10), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n347), .A2(KEYINPUT10), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(KEYINPUT3), .A2(G33), .ZN(new_n353));
  NAND2_X1  g0153(.A1(KEYINPUT3), .A2(G33), .ZN(new_n354));
  AOI21_X1  g0154(.A(G1698), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n283), .A2(new_n284), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n355), .A2(G222), .B1(new_n356), .B2(G77), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT70), .B(G223), .Z(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(G1698), .A3(new_n312), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n290), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n299), .B1(new_n279), .B2(new_n304), .ZN(new_n361));
  OAI21_X1  g0161(.A(G200), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n360), .A2(new_n361), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G190), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n350), .A2(new_n352), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT73), .B1(new_n268), .B2(new_n269), .ZN(new_n366));
  AOI211_X1 g0166(.A(new_n261), .B(new_n248), .C1(new_n264), .C2(new_n265), .ZN(new_n367));
  OAI221_X1 g0167(.A(G77), .B1(G1), .B2(new_n207), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G20), .A2(G77), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n369), .B1(new_n256), .B2(new_n370), .C1(new_n253), .C2(new_n336), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n248), .B1(new_n257), .B2(new_n266), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n307), .A2(G244), .ZN(new_n374));
  NOR2_X1   g0174(.A1(G232), .A2(G1698), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n280), .A2(G238), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n312), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n377), .B(new_n310), .C1(G107), .C2(new_n312), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(new_n378), .A3(new_n299), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n379), .A2(G179), .ZN(new_n380));
  INV_X1    g0180(.A(G169), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n373), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(G200), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n374), .A2(new_n378), .A3(G190), .A4(new_n299), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n384), .A2(new_n368), .A3(new_n372), .A4(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n364), .B1(new_n388), .B2(new_n363), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n351), .B1(new_n389), .B2(new_n349), .ZN(new_n390));
  INV_X1    g0190(.A(G179), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n363), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n381), .B1(new_n360), .B2(new_n361), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n343), .A3(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n365), .A2(new_n387), .A3(new_n390), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n312), .B2(G20), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n356), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n202), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(G58), .B(G68), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G20), .ZN(new_n402));
  INV_X1    g0202(.A(G159), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n402), .B1(new_n253), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n356), .B2(new_n207), .ZN(new_n406));
  NOR4_X1   g0206(.A1(new_n283), .A2(new_n284), .A3(new_n397), .A4(G20), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n250), .A2(new_n252), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(G159), .B1(new_n401), .B2(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(KEYINPUT16), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n405), .A2(new_n411), .A3(new_n248), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n336), .B1(new_n206), .B2(G20), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n340), .B1(new_n339), .B2(new_n336), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n279), .B2(G1698), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n312), .B1(G33), .B2(G87), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT78), .B1(new_n418), .B2(new_n290), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n279), .A2(G1698), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n420), .B1(G223), .B2(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G87), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT78), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n310), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n302), .A2(G232), .A3(new_n290), .A4(new_n303), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n299), .A2(new_n391), .A3(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n299), .B(new_n427), .C1(new_n418), .C2(new_n290), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n426), .A2(new_n428), .B1(new_n429), .B2(new_n381), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n415), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT18), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n388), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n419), .A2(new_n425), .ZN(new_n434));
  INV_X1    g0234(.A(G190), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n299), .A2(new_n435), .A3(new_n427), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n433), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n412), .A3(new_n414), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n437), .A2(KEYINPUT17), .A3(new_n412), .A4(new_n414), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n415), .A2(new_n430), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n432), .A2(new_n440), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n395), .A2(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n328), .A2(new_n332), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT84), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n257), .B1(new_n250), .B2(new_n252), .ZN(new_n448));
  XNOR2_X1  g0248(.A(G97), .B(G107), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT6), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G107), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n452), .A2(KEYINPUT6), .A3(G97), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n448), .B1(new_n455), .B2(G20), .ZN(new_n456));
  OAI211_X1 g0256(.A(KEYINPUT79), .B(G107), .C1(new_n406), .C2(new_n407), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n452), .B1(new_n398), .B2(new_n399), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n248), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n262), .A2(G97), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n206), .A2(G33), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n340), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  INV_X1    g0269(.A(G41), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT5), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(KEYINPUT80), .B2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(G45), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G1), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n476), .A2(new_n297), .A3(new_n310), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n476), .A2(G257), .A3(new_n290), .ZN(new_n478));
  OAI211_X1 g0278(.A(G244), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n312), .A2(KEYINPUT4), .A3(G244), .A4(new_n280), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  OAI211_X1 g0283(.A(G250), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  AOI211_X1 g0285(.A(new_n477), .B(new_n478), .C1(new_n485), .C2(new_n310), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n461), .A2(new_n468), .B1(new_n486), .B2(new_n391), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n483), .B(new_n484), .C1(new_n479), .C2(new_n480), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT4), .B1(new_n355), .B2(G244), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n310), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n298), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n491));
  INV_X1    g0291(.A(new_n478), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n381), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n490), .A2(new_n435), .A3(new_n491), .A4(new_n492), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n486), .B2(G200), .ZN(new_n496));
  OAI21_X1  g0296(.A(G107), .B1(new_n406), .B2(new_n407), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT79), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(new_n457), .A3(new_n456), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n467), .B1(new_n500), .B2(new_n248), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n487), .A2(new_n494), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT19), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n207), .B1(new_n286), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G87), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n466), .A3(new_n452), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n207), .B(G68), .C1(new_n283), .C2(new_n284), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n503), .B1(new_n256), .B2(new_n466), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(new_n248), .B1(new_n266), .B2(new_n370), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n340), .A2(G87), .A3(new_n464), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n290), .A2(G274), .A3(new_n475), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n206), .A2(G45), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n290), .A2(G250), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT81), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(G116), .ZN(new_n518));
  INV_X1    g0318(.A(G116), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(KEYINPUT81), .ZN(new_n520));
  OAI21_X1  g0320(.A(G33), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G238), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n522));
  OAI211_X1 g0322(.A(G244), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n516), .B1(new_n524), .B2(new_n310), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n511), .B(new_n512), .C1(new_n525), .C2(new_n388), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT83), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n525), .B2(G190), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(new_n527), .A3(G190), .ZN(new_n530));
  AOI211_X1 g0330(.A(G179), .B(new_n516), .C1(new_n310), .C2(new_n524), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n524), .A2(new_n310), .ZN(new_n532));
  INV_X1    g0332(.A(new_n516), .ZN(new_n533));
  AOI21_X1  g0333(.A(G169), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT82), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n465), .B2(new_n370), .ZN(new_n537));
  INV_X1    g0337(.A(new_n370), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n340), .A2(KEYINPUT82), .A3(new_n538), .A4(new_n464), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n511), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n529), .A2(new_n530), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n447), .B1(new_n502), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n486), .A2(new_n391), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n453), .B1(new_n449), .B2(new_n450), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n544), .A2(new_n207), .B1(new_n257), .B2(new_n253), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(KEYINPUT79), .B2(new_n459), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n269), .B1(new_n546), .B2(new_n499), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n543), .B(new_n494), .C1(new_n547), .C2(new_n467), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n496), .A2(new_n501), .ZN(new_n549));
  AND4_X1   g0349(.A1(new_n447), .A2(new_n541), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n542), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT81), .B(G116), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n552), .A2(G20), .A3(new_n249), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT86), .B1(new_n207), .B2(G107), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT23), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(KEYINPUT86), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n207), .B(G87), .C1(new_n283), .C2(new_n284), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT22), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n312), .A2(new_n563), .A3(new_n207), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n560), .B1(new_n559), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n248), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n262), .A2(G107), .ZN(new_n569));
  XNOR2_X1  g0369(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n465), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(G107), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G257), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n574));
  OAI211_X1 g0374(.A(G250), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G294), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n310), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n476), .A2(G264), .A3(new_n290), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n491), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n476), .A2(new_n290), .ZN(new_n582));
  AOI22_X1  g0382(.A1(G264), .A2(new_n582), .B1(new_n577), .B2(new_n310), .ZN(new_n583));
  AOI21_X1  g0383(.A(G200), .B1(new_n583), .B2(new_n491), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n568), .B(new_n573), .C1(new_n581), .C2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n264), .A2(new_n552), .A3(new_n265), .ZN(new_n586));
  AOI21_X1  g0386(.A(G20), .B1(G33), .B2(G283), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n249), .A2(G97), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n588), .B1(new_n246), .B2(new_n247), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n519), .A2(KEYINPUT81), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n517), .A2(G116), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n591), .A3(G20), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT20), .B1(new_n589), .B2(new_n592), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n586), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n519), .B1(new_n206), .B2(G33), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n271), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n476), .A2(G270), .A3(new_n290), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n598), .A2(new_n491), .ZN(new_n599));
  OAI211_X1 g0399(.A(G264), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n600));
  OAI211_X1 g0400(.A(G257), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n353), .A2(G303), .A3(new_n354), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n310), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G200), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n597), .B(new_n606), .C1(new_n435), .C2(new_n605), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n585), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT85), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(G169), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n597), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n596), .B1(new_n366), .B2(new_n367), .ZN(new_n613));
  INV_X1    g0413(.A(new_n594), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n592), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n586), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n605), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(G179), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n610), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n381), .B1(new_n599), .B2(new_n604), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n612), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n583), .A2(new_n391), .A3(new_n491), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n580), .A2(new_n381), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n568), .B2(new_n573), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n608), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n446), .A2(new_n551), .A3(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n394), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n432), .A2(new_n443), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n321), .A2(KEYINPUT77), .ZN(new_n632));
  INV_X1    g0432(.A(new_n325), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n323), .B2(KEYINPUT14), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n322), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n383), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n635), .A2(new_n278), .B1(new_n332), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n440), .A2(new_n441), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n631), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n365), .A2(new_n390), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n630), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n446), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n388), .B1(new_n532), .B2(new_n533), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n510), .A2(new_n248), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n266), .A2(new_n370), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n512), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n532), .A2(G190), .A3(new_n533), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n535), .A2(new_n540), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n548), .A2(new_n549), .A3(new_n649), .A4(new_n585), .ZN(new_n650));
  INV_X1    g0450(.A(new_n623), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n568), .A2(new_n573), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n624), .A2(new_n625), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n650), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n648), .A2(KEYINPUT83), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n532), .A2(new_n533), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G200), .ZN(new_n658));
  INV_X1    g0458(.A(new_n646), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n656), .A2(new_n658), .A3(new_n659), .A4(new_n530), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n525), .A2(new_n391), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n540), .B(new_n661), .C1(G169), .C2(new_n525), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT26), .B1(new_n548), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n649), .A2(new_n665), .A3(new_n487), .A4(new_n494), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n655), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n641), .B1(new_n642), .B2(new_n668), .ZN(G369));
  NAND2_X1  g0469(.A1(new_n276), .A2(new_n207), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n652), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n627), .B1(new_n585), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n654), .A2(new_n675), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n675), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n623), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n654), .B2(new_n675), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT88), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT88), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n597), .A2(new_n680), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n623), .B(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(new_n607), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n679), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(G399));
  NAND2_X1  g0492(.A1(new_n210), .A2(new_n470), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n206), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n506), .A2(G116), .ZN(new_n696));
  INV_X1    g0496(.A(new_n215), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n695), .A2(new_n696), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n490), .A2(new_n492), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n604), .A2(G179), .A3(new_n491), .A4(new_n598), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT89), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n583), .A2(new_n704), .A3(new_n525), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n704), .B1(new_n583), .B2(new_n525), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n703), .B(KEYINPUT30), .C1(new_n705), .C2(new_n706), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n618), .A2(G179), .A3(new_n525), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n493), .A3(new_n580), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n675), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT31), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n716), .A3(new_n675), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n628), .B(new_n680), .C1(new_n542), .C2(new_n550), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n700), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n680), .B1(new_n655), .B2(new_n667), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND4_X1   g0523(.A1(new_n548), .A2(new_n549), .A3(new_n649), .A4(new_n585), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT91), .B1(new_n623), .B2(new_n627), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n619), .A2(new_n622), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT91), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n654), .A4(new_n612), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n662), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n661), .B1(G169), .B2(new_n525), .ZN(new_n731));
  INV_X1    g0531(.A(new_n540), .ZN(new_n732));
  INV_X1    g0532(.A(new_n648), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n731), .A2(new_n732), .B1(new_n733), .B2(new_n526), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT90), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n548), .A2(new_n734), .A3(new_n735), .A4(new_n665), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n665), .B1(new_n548), .B2(new_n663), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT90), .ZN(new_n738));
  INV_X1    g0538(.A(new_n548), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT26), .A3(new_n649), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n736), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT29), .B(new_n680), .C1(new_n730), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n720), .B1(new_n723), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n699), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n275), .A2(G20), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G45), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT92), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n695), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n210), .A2(new_n312), .ZN(new_n750));
  INV_X1    g0550(.A(G355), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n750), .A2(new_n751), .B1(G116), .B2(new_n210), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n241), .A2(G45), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n210), .A2(new_n356), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n474), .B2(new_n697), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n213), .B1(new_n207), .B2(G169), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT93), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT93), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n749), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n207), .A2(new_n391), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n768), .A2(new_n435), .A3(G200), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n356), .B1(new_n769), .B2(G58), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n207), .A2(G179), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(new_n435), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G179), .A2(G200), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n207), .B1(new_n774), .B2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n773), .A2(G107), .B1(new_n776), .B2(G97), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n767), .A2(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n770), .B(new_n777), .C1(new_n202), .C2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n774), .A2(G20), .A3(new_n435), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n778), .A2(new_n435), .ZN(new_n785));
  AOI22_X1  g0585(.A1(KEYINPUT32), .A2(new_n784), .B1(new_n785), .B2(G50), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n771), .A2(G190), .A3(G200), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n786), .B1(KEYINPUT32), .B2(new_n784), .C1(new_n505), .C2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT94), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n789), .A2(KEYINPUT94), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n781), .B(new_n788), .C1(G77), .C2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n789), .A2(G311), .B1(G329), .B2(new_n783), .ZN(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  INV_X1    g0597(.A(new_n769), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n356), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n787), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G303), .B1(new_n773), .B2(G283), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT33), .B(G317), .Z(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(new_n802), .B2(new_n775), .C1(new_n780), .C2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n785), .B(KEYINPUT95), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n799), .B(new_n804), .C1(G326), .C2(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n795), .A2(new_n807), .A3(KEYINPUT96), .ZN(new_n808));
  INV_X1    g0608(.A(new_n760), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(KEYINPUT96), .B1(new_n795), .B2(new_n807), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n766), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n763), .B(KEYINPUT97), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n688), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n689), .A2(new_n748), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n688), .A2(G330), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT98), .Z(G396));
  AOI21_X1  g0618(.A(new_n680), .B1(new_n368), .B2(new_n372), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n819), .A2(KEYINPUT100), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n386), .B1(new_n819), .B2(KEYINPUT100), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n383), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n383), .A2(new_n675), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n721), .B(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n720), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT101), .Z(new_n830));
  AOI21_X1  g0630(.A(new_n749), .B1(new_n827), .B2(new_n828), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n760), .A2(new_n761), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n748), .B1(new_n833), .B2(new_n257), .ZN(new_n834));
  INV_X1    g0634(.A(new_n826), .ZN(new_n835));
  INV_X1    g0635(.A(G283), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n780), .A2(new_n836), .B1(new_n452), .B2(new_n787), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n798), .A2(new_n802), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n312), .B(new_n838), .C1(G311), .C2(new_n783), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n773), .A2(G87), .B1(new_n776), .B2(G97), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n839), .B(new_n840), .C1(new_n793), .C2(new_n552), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n837), .B(new_n841), .C1(G303), .C2(new_n785), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n769), .A2(G143), .B1(new_n785), .B2(G137), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n843), .B1(new_n333), .B2(new_n780), .C1(new_n793), .C2(new_n403), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n312), .B1(new_n782), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT99), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n800), .A2(G50), .B1(new_n776), .B2(G58), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n849), .B(new_n850), .C1(new_n202), .C2(new_n772), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n844), .B2(new_n845), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n842), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n834), .B1(new_n835), .B2(new_n762), .C1(new_n809), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n832), .A2(new_n854), .ZN(G384));
  NOR2_X1   g0655(.A1(new_n745), .A2(new_n206), .ZN(new_n856));
  INV_X1    g0656(.A(new_n673), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n415), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n431), .A2(new_n858), .A3(new_n438), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n431), .A2(new_n858), .A3(new_n861), .A4(new_n438), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(KEYINPUT103), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n858), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n444), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT103), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n859), .A2(new_n866), .A3(KEYINPUT37), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n863), .A2(new_n865), .A3(KEYINPUT38), .A4(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT104), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n871), .A2(new_n866), .B1(new_n444), .B2(new_n864), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n872), .B2(new_n863), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n863), .A2(new_n865), .A3(new_n867), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(KEYINPUT104), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT39), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT106), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n860), .A2(new_n862), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n865), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n868), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n879), .A2(new_n880), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n875), .A2(new_n876), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n869), .A3(new_n868), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n886), .B1(new_n890), .B2(new_n877), .ZN(new_n891));
  INV_X1    g0691(.A(new_n887), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT106), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n328), .A2(new_n675), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n888), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n721), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n824), .B1(new_n896), .B2(new_n835), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n278), .A2(new_n675), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n328), .A2(new_n332), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n332), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n278), .B(new_n675), .C1(new_n635), .C2(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n874), .A2(new_n878), .ZN(new_n904));
  INV_X1    g0704(.A(new_n631), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n903), .A2(new_n904), .B1(new_n905), .B2(new_n673), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n895), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n742), .A2(new_n446), .A3(new_n723), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n641), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n826), .B1(new_n899), .B2(new_n901), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n718), .A2(new_n719), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(new_n885), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT40), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n890), .A2(new_n916), .A3(new_n877), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n446), .A2(new_n912), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n700), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n856), .B1(new_n910), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n910), .B2(new_n921), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n214), .A2(new_n519), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT102), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n926), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT36), .Z(new_n930));
  OAI21_X1  g0730(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n215), .A2(new_n931), .B1(G50), .B2(new_n202), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(G1), .A3(new_n275), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n923), .A2(new_n930), .A3(new_n933), .ZN(G367));
  INV_X1    g0734(.A(new_n691), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n675), .B1(new_n547), .B2(new_n467), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n502), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT109), .Z(new_n938));
  NOR2_X1   g0738(.A1(new_n548), .A2(new_n680), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT110), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n675), .A2(new_n646), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT107), .Z(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n649), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT108), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT108), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n945), .A2(new_n662), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n943), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n739), .B1(new_n938), .B2(new_n627), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n675), .ZN(new_n956));
  INV_X1    g0756(.A(new_n681), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n941), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n956), .B1(new_n958), .B2(KEYINPUT42), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(KEYINPUT42), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n952), .B2(new_n951), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n954), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n693), .B(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n685), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT45), .B1(new_n685), .B2(new_n941), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n683), .A2(new_n684), .A3(new_n940), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT44), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n972), .A3(new_n691), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n935), .B1(new_n968), .B2(new_n971), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n679), .B1(new_n623), .B2(new_n680), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n957), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n689), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n973), .A2(new_n974), .A3(new_n743), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n965), .B1(new_n978), .B2(new_n743), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n747), .A2(G1), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n962), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n764), .B1(new_n210), .B2(new_n370), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n236), .A2(new_n754), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n749), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(G137), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n312), .B1(new_n782), .B2(new_n985), .C1(new_n798), .C2(new_n333), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n800), .A2(G58), .B1(new_n773), .B2(G77), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n202), .B2(new_n775), .C1(new_n403), .C2(new_n780), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n986), .B(new_n988), .C1(G50), .C2(new_n794), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n806), .A2(G143), .ZN(new_n990));
  XNOR2_X1  g0790(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n991));
  INV_X1    g0791(.A(new_n552), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n991), .B1(new_n800), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n783), .A2(G317), .ZN(new_n994));
  INV_X1    g0794(.A(G303), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n356), .B(new_n994), .C1(new_n798), .C2(new_n995), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n993), .B(new_n996), .C1(new_n794), .C2(G283), .ZN(new_n997));
  NAND2_X1  g0797(.A1(KEYINPUT46), .A2(G116), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n787), .A2(new_n998), .B1(new_n775), .B2(new_n452), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n780), .A2(new_n802), .B1(new_n772), .B2(new_n466), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n806), .C2(G311), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n989), .A2(new_n990), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT47), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n809), .B1(new_n1002), .B2(KEYINPUT47), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n984), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n813), .B2(new_n950), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n981), .A2(new_n1006), .ZN(G387));
  OR2_X1    g0807(.A1(new_n679), .A2(new_n813), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n750), .A2(new_n696), .B1(G107), .B2(new_n210), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n233), .A2(new_n474), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n696), .ZN(new_n1011));
  AOI211_X1 g0811(.A(G45), .B(new_n1011), .C1(G68), .C2(G77), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n336), .A2(G50), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n754), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1009), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n749), .B1(new_n1016), .B2(new_n765), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n789), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1018), .A2(new_n202), .B1(new_n333), .B2(new_n782), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n356), .B(new_n1019), .C1(G50), .C2(new_n769), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n800), .A2(G77), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n336), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n779), .A2(new_n1022), .B1(new_n538), .B2(new_n776), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n785), .A2(G159), .B1(new_n773), .B2(G97), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n312), .B1(new_n783), .B2(G326), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n787), .A2(new_n802), .B1(new_n775), .B2(new_n836), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT113), .Z(new_n1028));
  AOI22_X1  g0828(.A1(G317), .A2(new_n769), .B1(new_n779), .B2(G311), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n805), .B2(new_n797), .C1(new_n793), .C2(new_n995), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1026), .B1(new_n552), .B2(new_n772), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1025), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1017), .B1(new_n1037), .B2(new_n760), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n977), .A2(new_n980), .B1(new_n1008), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n977), .A2(new_n743), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n694), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n977), .A2(new_n743), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(G393));
  INV_X1    g0843(.A(new_n973), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n974), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1040), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n694), .A3(new_n978), .ZN(new_n1047));
  AND3_X1   g0847(.A1(new_n244), .A2(new_n210), .A3(new_n356), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n764), .B1(new_n466), .B2(new_n210), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n356), .B1(new_n783), .B2(G143), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n505), .B2(new_n772), .C1(new_n793), .C2(new_n336), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n775), .A2(new_n257), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n780), .A2(new_n254), .B1(new_n202), .B2(new_n787), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n769), .A2(G159), .B1(new_n785), .B2(G150), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT51), .Z(new_n1056));
  AOI22_X1  g0856(.A1(new_n769), .A2(G311), .B1(new_n785), .B2(G317), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  OAI221_X1 g0858(.A(new_n356), .B1(new_n782), .B2(new_n797), .C1(new_n1018), .C2(new_n802), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n787), .A2(new_n836), .B1(new_n775), .B2(new_n552), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n780), .A2(new_n995), .B1(new_n772), .B2(new_n452), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1054), .A2(new_n1056), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n749), .B1(new_n1048), .B2(new_n1049), .C1(new_n1063), .C2(new_n809), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n940), .B2(new_n763), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n980), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1047), .A2(new_n1067), .ZN(G390));
  NAND3_X1  g0868(.A1(new_n912), .A2(G330), .A3(new_n835), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n902), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n899), .A2(new_n901), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n720), .A3(new_n835), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n680), .B(new_n823), .C1(new_n730), .C2(new_n741), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1073), .A2(new_n825), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1070), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n902), .A2(new_n1069), .B1(new_n911), .B2(new_n720), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1075), .B1(new_n1076), .B2(new_n897), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n332), .A2(new_n636), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n638), .B1(new_n328), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n640), .B1(new_n1079), .B2(new_n905), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n720), .A2(new_n446), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n908), .A2(new_n1080), .A3(new_n1081), .A4(new_n394), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT114), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n641), .A2(KEYINPUT114), .A3(new_n908), .A4(new_n1081), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1077), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n880), .B1(new_n879), .B2(new_n887), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT106), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1087), .A2(new_n1088), .B1(new_n894), .B2(new_n903), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1074), .A2(new_n902), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n885), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1090), .A2(new_n894), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1072), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n903), .A2(new_n894), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n888), .B2(new_n893), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1072), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n1092), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1086), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1089), .A2(new_n1072), .A3(new_n1093), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1097), .B1(new_n1096), .B2(new_n1092), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1086), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1099), .A2(new_n694), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1100), .A2(new_n1101), .A3(new_n980), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n761), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n356), .B1(new_n783), .B2(G125), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT54), .B(G143), .Z(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT115), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1107), .B1(new_n847), .B2(new_n798), .C1(new_n793), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n800), .A2(G150), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT53), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n780), .A2(new_n985), .B1(new_n775), .B2(new_n403), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n785), .ZN(new_n1115));
  INV_X1    g0915(.A(G128), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1115), .A2(new_n1116), .B1(new_n772), .B2(new_n254), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .A4(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT116), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1115), .A2(new_n836), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1052), .B(new_n1120), .C1(G107), .C2(new_n779), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n356), .B1(new_n782), .B2(new_n802), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n202), .A2(new_n772), .B1(new_n787), .B2(new_n505), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(G116), .C2(new_n769), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1121), .B(new_n1124), .C1(new_n466), .C2(new_n793), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT117), .Z(new_n1126));
  AOI21_X1  g0926(.A(new_n809), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n748), .B(new_n1127), .C1(new_n336), .C2(new_n833), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1106), .A2(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1105), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1104), .A2(new_n1130), .ZN(G378));
  INV_X1    g0931(.A(new_n917), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n915), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1132), .A2(new_n1133), .B1(new_n913), .B2(KEYINPUT40), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n640), .A2(new_n394), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n343), .A2(new_n857), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1137), .B(new_n1138), .Z(new_n1139));
  NOR3_X1   g0939(.A1(new_n1134), .A2(new_n700), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1139), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n918), .B2(G330), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n907), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1139), .B1(new_n1134), .B2(new_n700), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n918), .A2(G330), .A3(new_n1141), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n1145), .A3(new_n895), .A4(new_n906), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n980), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1115), .A2(new_n519), .B1(new_n772), .B2(new_n201), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G97), .B2(new_n779), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n356), .A2(new_n470), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G283), .B2(new_n783), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n538), .A2(new_n789), .B1(new_n769), .B2(G107), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n800), .A2(G77), .B1(new_n776), .B2(G68), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT58), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G50), .B1(new_n249), .B2(new_n470), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1155), .A2(new_n1156), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1116), .A2(new_n798), .B1(new_n1018), .B2(new_n985), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G132), .B2(new_n779), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n785), .A2(G125), .B1(G150), .B2(new_n776), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n787), .C2(new_n1110), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n773), .A2(G159), .ZN(new_n1164));
  AOI211_X1 g0964(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1158), .B1(new_n1156), .B2(new_n1155), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n760), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n748), .B1(new_n833), .B2(new_n254), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(new_n1141), .C2(new_n762), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1148), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT118), .Z(new_n1174));
  NAND2_X1  g0974(.A1(new_n1103), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1176), .A2(KEYINPUT119), .A3(new_n895), .A4(new_n906), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT119), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1143), .A2(new_n1178), .A3(new_n1146), .ZN(new_n1179));
  AND4_X1   g0979(.A1(KEYINPUT57), .A2(new_n1175), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1103), .A2(new_n1174), .B1(new_n1146), .B2(new_n1143), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n694), .B1(new_n1181), .B2(KEYINPUT57), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1172), .B1(new_n1180), .B2(new_n1182), .ZN(G375));
  AND3_X1   g0983(.A1(new_n1070), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n897), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n1173), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1086), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(new_n965), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT120), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1077), .A2(new_n980), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n794), .A2(G107), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1115), .A2(new_n802), .B1(new_n787), .B2(new_n466), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n992), .B2(new_n779), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n356), .B1(new_n782), .B2(new_n995), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n769), .B2(G283), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n773), .A2(G77), .B1(new_n776), .B2(new_n538), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1192), .A2(new_n1194), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n312), .B1(new_n772), .B2(new_n201), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT121), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n798), .A2(new_n985), .B1(new_n1116), .B2(new_n782), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G150), .B2(new_n789), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1115), .A2(new_n847), .B1(new_n787), .B2(new_n403), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G50), .B2(new_n776), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n780), .C2(new_n1110), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1198), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n760), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n748), .B1(new_n833), .B2(new_n202), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n1071), .C2(new_n762), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1191), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1190), .A2(new_n1211), .ZN(G381));
  OR3_X1    g1012(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT122), .Z(new_n1215));
  NOR2_X1   g1015(.A1(G375), .A2(G378), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(G407));
  INV_X1    g1017(.A(new_n1216), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G407), .B(G213), .C1(G343), .C2(new_n1218), .ZN(G409));
  XOR2_X1   g1019(.A(G393), .B(G396), .Z(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n981), .A2(G390), .A3(new_n1006), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G390), .B1(new_n981), .B2(new_n1006), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1221), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G390), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G387), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n1220), .A3(new_n1222), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT61), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1225), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1230), .A2(KEYINPUT125), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n674), .A2(G213), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1175), .A2(new_n964), .A3(new_n1147), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1179), .A2(new_n1177), .A3(new_n980), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1104), .A2(new_n1130), .A3(new_n1171), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1232), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G375), .B2(G378), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT123), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1187), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n694), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1240), .B1(new_n1187), .B2(new_n1086), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1239), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1188), .A2(KEYINPUT60), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n693), .B1(new_n1187), .B2(new_n1240), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(KEYINPUT123), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G384), .B1(new_n1248), .B2(new_n1211), .ZN(new_n1249));
  INV_X1    g1049(.A(G384), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1250), .B(new_n1210), .C1(new_n1244), .C2(new_n1247), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1238), .A2(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT63), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1232), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(G2897), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1252), .A2(new_n1255), .A3(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(KEYINPUT124), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1242), .A2(new_n1239), .A3(new_n1243), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT123), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1211), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1250), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1248), .A2(G384), .A3(new_n1211), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1255), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1260), .A2(new_n1266), .A3(new_n1257), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1238), .B1(new_n1259), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1230), .A2(KEYINPUT125), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1231), .A2(new_n1254), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT126), .B1(new_n1268), .B2(KEYINPUT61), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  NOR4_X1   g1073(.A1(new_n1249), .A2(new_n1251), .A3(KEYINPUT124), .A4(new_n1257), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1258), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n1260), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1273), .B(new_n1229), .C1(new_n1276), .C2(new_n1238), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G375), .A2(G378), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1237), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1252), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1278), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1238), .A2(KEYINPUT62), .A3(new_n1252), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1272), .A2(new_n1277), .A3(KEYINPUT127), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1267), .A2(new_n1259), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1289), .B2(new_n1281), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1290), .A2(new_n1273), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT127), .B1(new_n1291), .B2(new_n1272), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1271), .B1(new_n1288), .B2(new_n1292), .ZN(G405));
  NAND2_X1  g1093(.A1(new_n1218), .A2(new_n1279), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1294), .B(new_n1282), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(new_n1287), .ZN(G402));
endmodule


