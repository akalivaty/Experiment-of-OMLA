

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581;

  INV_X1 U320 ( .A(KEYINPUT86), .ZN(n324) );
  XNOR2_X1 U321 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U322 ( .A(n368), .B(n422), .Z(n288) );
  XOR2_X1 U323 ( .A(n350), .B(n349), .Z(n289) );
  XOR2_X1 U324 ( .A(n345), .B(n379), .Z(n290) );
  INV_X1 U325 ( .A(KEYINPUT112), .ZN(n396) );
  XNOR2_X1 U326 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n294) );
  XNOR2_X1 U327 ( .A(n396), .B(KEYINPUT47), .ZN(n397) );
  XNOR2_X1 U328 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U329 ( .A(n398), .B(n397), .ZN(n403) );
  NOR2_X1 U330 ( .A1(n478), .A2(n574), .ZN(n467) );
  XNOR2_X1 U331 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U332 ( .A(n351), .B(n289), .ZN(n352) );
  NOR2_X1 U333 ( .A1(n461), .A2(n564), .ZN(n431) );
  INV_X1 U334 ( .A(G183GAT), .ZN(n447) );
  INV_X1 U335 ( .A(G29GAT), .ZN(n472) );
  XNOR2_X1 U336 ( .A(n447), .B(KEYINPUT122), .ZN(n448) );
  XNOR2_X1 U337 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U338 ( .A(n449), .B(n448), .ZN(G1350GAT) );
  XNOR2_X1 U339 ( .A(n475), .B(n474), .ZN(G1328GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n292) );
  XNOR2_X1 U341 ( .A(G64GAT), .B(G8GAT), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n309) );
  XNOR2_X1 U343 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n293), .B(KEYINPUT70), .ZN(n361) );
  XNOR2_X1 U345 ( .A(n294), .B(KEYINPUT13), .ZN(n345) );
  XNOR2_X1 U346 ( .A(n361), .B(n345), .ZN(n307) );
  XOR2_X1 U347 ( .A(G211GAT), .B(G78GAT), .Z(n296) );
  XNOR2_X1 U348 ( .A(G155GAT), .B(G22GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U350 ( .A(G183GAT), .B(G15GAT), .Z(n298) );
  XNOR2_X1 U351 ( .A(G127GAT), .B(G71GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U353 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U354 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n302) );
  NAND2_X1 U355 ( .A1(G231GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U357 ( .A(KEYINPUT15), .B(n303), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n574) );
  INV_X1 U361 ( .A(n574), .ZN(n545) );
  XNOR2_X1 U362 ( .A(G204GAT), .B(KEYINPUT88), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n310), .B(KEYINPUT21), .ZN(n311) );
  XOR2_X1 U364 ( .A(n311), .B(KEYINPUT87), .Z(n313) );
  XNOR2_X1 U365 ( .A(G218GAT), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n334) );
  XOR2_X1 U367 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n315) );
  XNOR2_X1 U368 ( .A(G197GAT), .B(KEYINPUT91), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U370 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n317) );
  XNOR2_X1 U371 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n329) );
  XOR2_X1 U374 ( .A(G141GAT), .B(G22GAT), .Z(n368) );
  XOR2_X1 U375 ( .A(G155GAT), .B(KEYINPUT3), .Z(n321) );
  XNOR2_X1 U376 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n422) );
  NAND2_X1 U378 ( .A1(G228GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n288), .B(n322), .ZN(n327) );
  XNOR2_X1 U380 ( .A(G148GAT), .B(G106GAT), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n323), .B(G78GAT), .ZN(n348) );
  XNOR2_X1 U382 ( .A(n348), .B(KEYINPUT85), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n334), .B(n330), .ZN(n450) );
  INV_X1 U385 ( .A(n450), .ZN(n461) );
  XOR2_X1 U386 ( .A(G92GAT), .B(G64GAT), .Z(n343) );
  XOR2_X1 U387 ( .A(n343), .B(KEYINPUT96), .Z(n332) );
  NAND2_X1 U388 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(n333), .ZN(n338) );
  XOR2_X1 U391 ( .A(G8GAT), .B(G197GAT), .Z(n369) );
  XOR2_X1 U392 ( .A(n369), .B(n334), .Z(n336) );
  XNOR2_X1 U393 ( .A(G36GAT), .B(G190GAT), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U396 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n340) );
  XNOR2_X1 U397 ( .A(KEYINPUT19), .B(G176GAT), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U399 ( .A(G183GAT), .B(n341), .Z(n445) );
  XNOR2_X1 U400 ( .A(n342), .B(n445), .ZN(n492) );
  INV_X1 U401 ( .A(n492), .ZN(n515) );
  XNOR2_X1 U402 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n405) );
  XNOR2_X1 U403 ( .A(G176GAT), .B(G204GAT), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n355) );
  XOR2_X1 U405 ( .A(G85GAT), .B(KEYINPUT73), .Z(n379) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n290), .B(n346), .ZN(n353) );
  XNOR2_X1 U408 ( .A(G120GAT), .B(G99GAT), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n347), .B(G71GAT), .ZN(n440) );
  XNOR2_X1 U410 ( .A(n440), .B(n348), .ZN(n351) );
  XOR2_X1 U411 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n350) );
  XNOR2_X1 U412 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n570) );
  XNOR2_X1 U414 ( .A(KEYINPUT41), .B(n570), .ZN(n553) );
  XOR2_X1 U415 ( .A(KEYINPUT66), .B(KEYINPUT64), .Z(n357) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n358), .B(KEYINPUT65), .Z(n363) );
  XOR2_X1 U419 ( .A(G169GAT), .B(G15GAT), .Z(n360) );
  XNOR2_X1 U420 ( .A(G113GAT), .B(G43GAT), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n433) );
  XNOR2_X1 U422 ( .A(n361), .B(n433), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U424 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n365) );
  XNOR2_X1 U425 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U427 ( .A(n367), .B(n366), .Z(n371) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n376) );
  XOR2_X1 U430 ( .A(KEYINPUT8), .B(G50GAT), .Z(n373) );
  XNOR2_X1 U431 ( .A(KEYINPUT7), .B(G36GAT), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U433 ( .A(G29GAT), .B(n374), .Z(n392) );
  INV_X1 U434 ( .A(n392), .ZN(n375) );
  XOR2_X1 U435 ( .A(n376), .B(n375), .Z(n538) );
  NOR2_X1 U436 ( .A1(n553), .A2(n538), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n377), .B(KEYINPUT46), .ZN(n378) );
  NOR2_X1 U438 ( .A1(n574), .A2(n378), .ZN(n395) );
  XOR2_X1 U439 ( .A(G99GAT), .B(G92GAT), .Z(n381) );
  XOR2_X1 U440 ( .A(G134GAT), .B(G190GAT), .Z(n432) );
  XNOR2_X1 U441 ( .A(n379), .B(n432), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U443 ( .A(n382), .B(G106GAT), .Z(n387) );
  XOR2_X1 U444 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n384) );
  XNOR2_X1 U445 ( .A(G162GAT), .B(G43GAT), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n385), .B(G218GAT), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U449 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n389) );
  NAND2_X1 U450 ( .A1(G232GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U452 ( .A(n391), .B(n390), .Z(n394) );
  XNOR2_X1 U453 ( .A(n392), .B(KEYINPUT11), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n560) );
  NAND2_X1 U455 ( .A1(n395), .A2(n560), .ZN(n398) );
  XOR2_X1 U456 ( .A(KEYINPUT36), .B(n560), .Z(n576) );
  NAND2_X1 U457 ( .A1(n576), .A2(n574), .ZN(n399) );
  XNOR2_X1 U458 ( .A(KEYINPUT45), .B(n399), .ZN(n400) );
  NOR2_X1 U459 ( .A1(n570), .A2(n400), .ZN(n401) );
  INV_X1 U460 ( .A(n538), .ZN(n566) );
  XNOR2_X1 U461 ( .A(KEYINPUT71), .B(n566), .ZN(n551) );
  NAND2_X1 U462 ( .A1(n401), .A2(n551), .ZN(n402) );
  NAND2_X1 U463 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n535) );
  NOR2_X1 U465 ( .A1(n515), .A2(n535), .ZN(n406) );
  XNOR2_X1 U466 ( .A(KEYINPUT54), .B(n406), .ZN(n429) );
  XOR2_X1 U467 ( .A(G1GAT), .B(G113GAT), .Z(n408) );
  XNOR2_X1 U468 ( .A(G148GAT), .B(G120GAT), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U470 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n410) );
  XNOR2_X1 U471 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U473 ( .A(n412), .B(n411), .Z(n419) );
  XOR2_X1 U474 ( .A(G127GAT), .B(KEYINPUT0), .Z(n414) );
  XNOR2_X1 U475 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n441) );
  XOR2_X1 U477 ( .A(G85GAT), .B(n441), .Z(n416) );
  XNOR2_X1 U478 ( .A(G29GAT), .B(G141GAT), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(G134GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n428) );
  XOR2_X1 U482 ( .A(KEYINPUT95), .B(KEYINPUT92), .Z(n421) );
  XNOR2_X1 U483 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n426) );
  XOR2_X1 U485 ( .A(n422), .B(KEYINPUT5), .Z(n424) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U488 ( .A(n426), .B(n425), .Z(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n471) );
  INV_X1 U490 ( .A(n471), .ZN(n513) );
  NAND2_X1 U491 ( .A1(n429), .A2(n513), .ZN(n564) );
  XNOR2_X1 U492 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n446) );
  XOR2_X1 U494 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U497 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n437) );
  XNOR2_X1 U498 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U500 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n524) );
  NAND2_X1 U504 ( .A1(n446), .A2(n524), .ZN(n559) );
  NOR2_X1 U505 ( .A1(n545), .A2(n559), .ZN(n449) );
  NAND2_X1 U506 ( .A1(n524), .A2(n492), .ZN(n451) );
  NAND2_X1 U507 ( .A1(n451), .A2(n450), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n452), .B(KEYINPUT25), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n453), .B(KEYINPUT98), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n515), .B(KEYINPUT27), .ZN(n460) );
  INV_X1 U511 ( .A(n524), .ZN(n517) );
  NAND2_X1 U512 ( .A1(n517), .A2(n461), .ZN(n454) );
  XNOR2_X1 U513 ( .A(KEYINPUT26), .B(n454), .ZN(n565) );
  NOR2_X1 U514 ( .A1(n460), .A2(n565), .ZN(n455) );
  NOR2_X1 U515 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U516 ( .A(KEYINPUT99), .B(n457), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n458), .A2(n513), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT100), .ZN(n465) );
  XNOR2_X1 U519 ( .A(n517), .B(KEYINPUT84), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n513), .A2(n460), .ZN(n537) );
  XOR2_X1 U521 ( .A(n461), .B(KEYINPUT28), .Z(n520) );
  NAND2_X1 U522 ( .A1(n537), .A2(n520), .ZN(n523) );
  XNOR2_X1 U523 ( .A(n523), .B(KEYINPUT97), .ZN(n462) );
  NAND2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U526 ( .A(KEYINPUT101), .B(n466), .ZN(n478) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT106), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n468), .A2(n576), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n469), .B(KEYINPUT37), .ZN(n512) );
  NOR2_X1 U530 ( .A1(n551), .A2(n570), .ZN(n482) );
  NAND2_X1 U531 ( .A1(n512), .A2(n482), .ZN(n470) );
  XOR2_X2 U532 ( .A(KEYINPUT38), .B(n470), .Z(n498) );
  NAND2_X1 U533 ( .A1(n498), .A2(n471), .ZN(n475) );
  XOR2_X1 U534 ( .A(KEYINPUT39), .B(KEYINPUT107), .Z(n473) );
  XOR2_X1 U535 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n477) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(n484) );
  BUF_X1 U538 ( .A(n478), .Z(n481) );
  NAND2_X1 U539 ( .A1(n560), .A2(n574), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT16), .B(n479), .ZN(n480) );
  NOR2_X1 U541 ( .A1(n481), .A2(n480), .ZN(n502) );
  NAND2_X1 U542 ( .A1(n482), .A2(n502), .ZN(n489) );
  NOR2_X1 U543 ( .A1(n513), .A2(n489), .ZN(n483) );
  XOR2_X1 U544 ( .A(n484), .B(n483), .Z(G1324GAT) );
  NOR2_X1 U545 ( .A1(n515), .A2(n489), .ZN(n485) );
  XOR2_X1 U546 ( .A(G8GAT), .B(n485), .Z(G1325GAT) );
  NOR2_X1 U547 ( .A1(n517), .A2(n489), .ZN(n487) );
  XNOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n520), .A2(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1327GAT) );
  NAND2_X1 U554 ( .A1(n498), .A2(n492), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(KEYINPUT108), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n498), .A2(n524), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n495), .B(KEYINPUT40), .ZN(n496) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  XOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT109), .Z(n500) );
  INV_X1 U561 ( .A(n520), .ZN(n497) );
  NAND2_X1 U562 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  NOR2_X1 U564 ( .A1(n566), .A2(n553), .ZN(n501) );
  XNOR2_X1 U565 ( .A(KEYINPUT110), .B(n501), .ZN(n511) );
  NAND2_X1 U566 ( .A1(n502), .A2(n511), .ZN(n507) );
  NOR2_X1 U567 ( .A1(n513), .A2(n507), .ZN(n503) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n503), .Z(n504) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n515), .A2(n507), .ZN(n505) );
  XOR2_X1 U571 ( .A(G64GAT), .B(n505), .Z(G1333GAT) );
  NOR2_X1 U572 ( .A1(n517), .A2(n507), .ZN(n506) );
  XOR2_X1 U573 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U574 ( .A1(n520), .A2(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U577 ( .A(G78GAT), .B(n510), .Z(G1335GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n519) );
  NOR2_X1 U579 ( .A1(n513), .A2(n519), .ZN(n514) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n519), .ZN(n516) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n519), .ZN(n518) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(n521), .Z(n522) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n535), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n532) );
  NOR2_X1 U590 ( .A1(n551), .A2(n532), .ZN(n526) );
  XOR2_X1 U591 ( .A(G113GAT), .B(n526), .Z(G1340GAT) );
  NOR2_X1 U592 ( .A1(n553), .A2(n532), .ZN(n528) );
  XNOR2_X1 U593 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(n529), .ZN(G1341GAT) );
  NOR2_X1 U596 ( .A1(n545), .A2(n532), .ZN(n530) );
  XOR2_X1 U597 ( .A(KEYINPUT50), .B(n530), .Z(n531) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  NOR2_X1 U599 ( .A1(n560), .A2(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  NOR2_X1 U602 ( .A1(n565), .A2(n535), .ZN(n536) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n548) );
  NOR2_X1 U604 ( .A1(n538), .A2(n548), .ZN(n540) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1344GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n542) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n553), .A2(n548), .ZN(n543) );
  XOR2_X1 U611 ( .A(n544), .B(n543), .Z(G1345GAT) );
  NOR2_X1 U612 ( .A1(n545), .A2(n548), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1346GAT) );
  NOR2_X1 U615 ( .A1(n560), .A2(n548), .ZN(n549) );
  XOR2_X1 U616 ( .A(KEYINPUT118), .B(n549), .Z(n550) );
  XNOR2_X1 U617 ( .A(G162GAT), .B(n550), .ZN(G1347GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n559), .ZN(n552) );
  XOR2_X1 U619 ( .A(G169GAT), .B(n552), .Z(G1348GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n559), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(KEYINPUT120), .B(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U627 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n577) );
  NAND2_X1 U632 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n572) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n577), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1355GAT) );
endmodule

