//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n645, new_n646, new_n649, new_n651, new_n652, new_n653, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G567), .ZN(new_n460));
  INV_X1    g035(.A(G2106), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n466), .A2(new_n468), .A3(G137), .A4(new_n464), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n477), .A2(new_n464), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g059(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G112), .B2(new_n464), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n480), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT68), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n464), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n489), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n464), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n477), .A2(new_n499), .A3(G138), .A4(new_n464), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n503), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT69), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n503), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n516), .A2(G88), .A3(new_n505), .A4(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(G50), .A3(G543), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n518), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n511), .B1(new_n521), .B2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  AOI211_X1 g099(.A(KEYINPUT71), .B(new_n504), .C1(new_n514), .C2(new_n515), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n516), .B2(new_n505), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n504), .B1(new_n514), .B2(new_n515), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(new_n517), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  AND2_X1   g108(.A1(KEYINPUT6), .A2(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(KEYINPUT6), .A2(G651), .ZN(new_n535));
  OAI21_X1  g110(.A(G543), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g113(.A(KEYINPUT72), .B(G543), .C1(new_n534), .C2(new_n535), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n533), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n529), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n532), .A2(G90), .B1(new_n540), .B2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n528), .B2(G64), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  OAI211_X1 g125(.A(KEYINPUT73), .B(new_n546), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n530), .A2(new_n526), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n553), .A2(G64), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n550), .B1(new_n555), .B2(new_n547), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n540), .A2(G52), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n558), .B2(new_n531), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n552), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n551), .A2(new_n560), .ZN(G171));
  AND3_X1   g136(.A1(new_n553), .A2(G56), .A3(new_n554), .ZN(new_n562));
  AND2_X1   g137(.A1(G68), .A2(G543), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n532), .A2(G81), .B1(new_n540), .B2(G43), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  OAI211_X1 g148(.A(G53), .B(G543), .C1(new_n534), .C2(new_n535), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT75), .B1(new_n574), .B2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n517), .A2(new_n576), .A3(G53), .A4(G543), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n574), .B2(KEYINPUT74), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n574), .A2(KEYINPUT74), .ZN(new_n582));
  AND4_X1   g157(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT9), .A4(new_n577), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT76), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n577), .A3(KEYINPUT9), .ZN(new_n585));
  INV_X1    g160(.A(new_n575), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n579), .A2(new_n581), .A3(new_n577), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G78), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G65), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n508), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n532), .A2(G91), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n591), .A2(new_n598), .ZN(G299));
  AND2_X1   g174(.A1(new_n551), .A2(new_n560), .ZN(G301));
  INV_X1    g175(.A(G168), .ZN(G286));
  NAND3_X1  g176(.A1(new_n530), .A2(G87), .A3(new_n517), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(G74), .B1(new_n553), .B2(new_n554), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n550), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(G288));
  NAND3_X1  g187(.A1(new_n516), .A2(G61), .A3(new_n505), .ZN(new_n613));
  NAND2_X1  g188(.A1(G73), .A2(G543), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G651), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n516), .A2(G86), .A3(new_n505), .A4(new_n517), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n616), .A2(new_n619), .ZN(G305));
  AOI22_X1  g195(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n621), .A2(new_n550), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n540), .A2(G47), .ZN(new_n624));
  INV_X1    g199(.A(G85), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n531), .ZN(new_n626));
  OR3_X1    g201(.A1(new_n622), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n623), .B1(new_n622), .B2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(G290));
  NAND4_X1  g204(.A1(new_n516), .A2(G92), .A3(new_n505), .A4(new_n517), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT79), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n530), .A2(new_n632), .A3(G92), .A4(new_n517), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n631), .A2(KEYINPUT10), .A3(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n540), .A2(G54), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n530), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n550), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(KEYINPUT10), .B1(new_n631), .B2(new_n633), .ZN(new_n639));
  NOR3_X1   g214(.A1(new_n635), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n641), .A2(G868), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g218(.A(new_n642), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g219(.A1(G286), .A2(G868), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n597), .B1(new_n584), .B2(new_n590), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(G868), .ZN(G297));
  OAI21_X1  g222(.A(new_n645), .B1(new_n646), .B2(G868), .ZN(G280));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n640), .B1(new_n649), .B2(G860), .ZN(G148));
  NOR2_X1   g225(.A1(new_n641), .A2(G559), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G868), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g229(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g230(.A1(new_n481), .A2(G2104), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT12), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT80), .B(KEYINPUT13), .Z(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n479), .A2(G123), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n481), .A2(G135), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n464), .A2(G111), .ZN(new_n664));
  OAI21_X1  g239(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n662), .B(new_n663), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT81), .B(G2096), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n660), .A2(new_n661), .A3(new_n668), .ZN(G156));
  XNOR2_X1  g244(.A(G2427), .B(G2438), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2430), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(KEYINPUT14), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1341), .B(G1348), .Z(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2451), .B(G2454), .Z(new_n680));
  XNOR2_X1  g255(.A(G2443), .B(G2446), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(G14), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT83), .ZN(G401));
  XOR2_X1   g261(.A(G2084), .B(G2090), .Z(new_n687));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  NOR2_X1   g263(.A1(G2072), .A2(G2078), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n687), .B(new_n688), .C1(new_n444), .C2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT18), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(KEYINPUT84), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n444), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n687), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(KEYINPUT17), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n694), .B(new_n695), .C1(new_n692), .C2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n696), .A2(new_n692), .A3(new_n687), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n691), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(G2100), .Z(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT85), .B(G2096), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G227));
  XOR2_X1   g278(.A(G1971), .B(G1976), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT19), .ZN(new_n705));
  XOR2_X1   g280(.A(G1956), .B(G2474), .Z(new_n706));
  XOR2_X1   g281(.A(G1961), .B(G1966), .Z(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT20), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n707), .ZN(new_n711));
  NOR3_X1   g286(.A1(new_n705), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n705), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1991), .B(G1996), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(G1981), .B(G1986), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(G229));
  XOR2_X1   g295(.A(KEYINPUT31), .B(G11), .Z(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n666), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT30), .B(G28), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n721), .B(new_n723), .C1(new_n722), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  NOR2_X1   g301(.A1(G168), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(G21), .ZN(new_n728));
  INV_X1    g303(.A(G1966), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n729), .B2(new_n728), .ZN(new_n731));
  NOR2_X1   g306(.A1(G5), .A2(G16), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT94), .Z(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G171), .B2(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G1961), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n726), .A2(G19), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n567), .B2(new_n726), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G1341), .Z(new_n741));
  NOR2_X1   g316(.A1(G4), .A2(G16), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT88), .Z(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n641), .B2(new_n726), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1348), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n722), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT28), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n479), .A2(G128), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n481), .A2(G140), .ZN(new_n749));
  OR2_X1    g324(.A1(G104), .A2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n750), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n747), .B1(new_n753), .B2(new_n722), .ZN(new_n754));
  INV_X1    g329(.A(G2067), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n741), .A2(new_n745), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT89), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  AND3_X1   g337(.A1(new_n481), .A2(KEYINPUT90), .A3(G139), .ZN(new_n763));
  AOI21_X1  g338(.A(KEYINPUT90), .B1(new_n481), .B2(G139), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n761), .B1(new_n464), .B2(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G33), .B(new_n765), .S(G29), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(new_n442), .ZN(new_n767));
  INV_X1    g342(.A(G34), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(KEYINPUT24), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(KEYINPUT24), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n722), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G160), .B2(new_n722), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT91), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G2084), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n481), .A2(G141), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n473), .A2(G105), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  INV_X1    g354(.A(G129), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n478), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(new_n722), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n722), .B2(G32), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT27), .B(G1996), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT92), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n767), .A2(new_n774), .A3(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT93), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n734), .A2(G1961), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(KEYINPUT93), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n722), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n722), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT29), .B(G2090), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n786), .B2(new_n784), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n773), .A2(G2084), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n722), .A2(G27), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT96), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n491), .A2(new_n493), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n495), .B1(new_n800), .B2(G2105), .ZN(new_n801));
  AND4_X1   g376(.A1(G126), .A2(new_n466), .A3(new_n468), .A4(G2105), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n498), .A2(new_n500), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(G29), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(new_n443), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n796), .A2(new_n797), .A3(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n789), .A2(new_n790), .A3(new_n791), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n726), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n646), .B2(new_n726), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1956), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n738), .A2(new_n758), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  MUX2_X1   g390(.A(G23), .B(new_n607), .S(G16), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT33), .ZN(new_n817));
  INV_X1    g392(.A(G1976), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G22), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G166), .B2(G16), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1971), .ZN(new_n822));
  MUX2_X1   g397(.A(G6), .B(G305), .S(G16), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT32), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1981), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n819), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n726), .A2(G24), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G290), .B2(G16), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT87), .B(G1986), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n722), .A2(G25), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT86), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n479), .A2(G119), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n481), .A2(G131), .ZN(new_n837));
  OR2_X1    g412(.A1(G95), .A2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n835), .B1(new_n841), .B2(new_n722), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G1991), .Z(new_n843));
  XOR2_X1   g418(.A(new_n842), .B(new_n843), .Z(new_n844));
  NOR3_X1   g419(.A1(new_n832), .A2(new_n833), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n828), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n826), .A2(new_n827), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT36), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OR3_X1    g423(.A1(new_n846), .A2(KEYINPUT36), .A3(new_n847), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n815), .B1(new_n848), .B2(new_n849), .ZN(G311));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n814), .ZN(G150));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n538), .B2(new_n539), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n530), .A2(G93), .A3(new_n517), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT72), .B1(new_n517), .B2(G543), .ZN(new_n858));
  INV_X1    g433(.A(new_n539), .ZN(new_n859));
  OAI21_X1  g434(.A(G55), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n530), .A2(G93), .A3(new_n517), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(KEYINPUT98), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G67), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n525), .A2(new_n527), .A3(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(G80), .A2(G543), .ZN(new_n866));
  OAI21_X1  g441(.A(G651), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(KEYINPUT100), .B(G860), .Z(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n640), .A2(G559), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT99), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n874), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n868), .A2(new_n566), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n564), .A2(new_n863), .A3(new_n867), .A4(new_n565), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n877), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT39), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n883), .A2(KEYINPUT101), .A3(new_n870), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT101), .B1(new_n883), .B2(new_n870), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n873), .B1(new_n884), .B2(new_n885), .ZN(G145));
  XOR2_X1   g461(.A(new_n840), .B(KEYINPUT105), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n657), .ZN(new_n888));
  INV_X1    g463(.A(new_n782), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n765), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n888), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n752), .B(G164), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n479), .A2(G130), .B1(new_n481), .B2(G142), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n894), .A2(KEYINPUT104), .ZN(new_n895));
  OR3_X1    g470(.A1(new_n464), .A2(KEYINPUT103), .A3(G118), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT103), .B1(new_n464), .B2(G118), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n896), .B(new_n897), .C1(KEYINPUT104), .C2(new_n894), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n893), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n892), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n891), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n666), .B(G160), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n487), .ZN(new_n903));
  AOI21_X1  g478(.A(G37), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(new_n903), .B2(new_n901), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g481(.A(new_n607), .B(G305), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n627), .A2(G303), .A3(new_n628), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G303), .B1(new_n627), .B2(new_n628), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n907), .A3(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT42), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n652), .A2(new_n881), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n651), .A2(new_n880), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n640), .A2(new_n591), .A3(new_n598), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n646), .A2(new_n640), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n920), .B(KEYINPUT41), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT41), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  NAND2_X1  g499(.A1(G299), .A2(new_n641), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n646), .A2(new_n640), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n928), .A3(KEYINPUT107), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n919), .A2(new_n923), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n921), .A2(new_n922), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n917), .A2(new_n918), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT106), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n916), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n916), .B1(new_n933), .B2(new_n930), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G868), .B2(new_n869), .ZN(G295));
  OAI21_X1  g512(.A(new_n936), .B1(G868), .B2(new_n869), .ZN(G331));
  AOI22_X1  g513(.A1(new_n867), .A2(new_n863), .B1(new_n564), .B2(new_n565), .ZN(new_n939));
  AND4_X1   g514(.A1(new_n564), .A2(new_n863), .A3(new_n867), .A4(new_n565), .ZN(new_n940));
  OAI21_X1  g515(.A(G301), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n878), .A2(G171), .A3(new_n879), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n941), .A2(G168), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G168), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n923), .B(new_n929), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n942), .ZN(new_n946));
  AOI21_X1  g521(.A(G171), .B1(new_n878), .B2(new_n879), .ZN(new_n947));
  OAI21_X1  g522(.A(G286), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n941), .A2(G168), .A3(new_n942), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n931), .A3(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n945), .A2(new_n915), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n943), .A2(new_n944), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n929), .A2(new_n923), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n915), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n915), .B1(new_n950), .B2(new_n945), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT108), .B1(new_n959), .B2(G37), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT43), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n951), .A2(G37), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n948), .A2(new_n949), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n924), .A2(new_n928), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(KEYINPUT109), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n950), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT109), .B1(new_n963), .B2(new_n964), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n955), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n962), .A2(new_n968), .A3(KEYINPUT43), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT44), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n958), .B2(new_n960), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n962), .A2(new_n968), .A3(new_n972), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(G164), .B2(G1384), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n471), .A2(new_n475), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n752), .B(new_n755), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n984), .B2(new_n889), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n986));
  INV_X1    g561(.A(G1996), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  NOR4_X1   g563(.A1(new_n978), .A2(KEYINPUT46), .A3(new_n981), .A4(G1996), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n990), .B(KEYINPUT47), .Z(new_n991));
  NOR2_X1   g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n992), .A2(KEYINPUT48), .A3(new_n982), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT48), .B1(new_n992), .B2(new_n982), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n841), .A2(new_n843), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n841), .A2(new_n843), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n978), .B(new_n981), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n982), .A2(G1996), .A3(new_n889), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(KEYINPUT110), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(KEYINPUT110), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n889), .A2(G1996), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n982), .B1(new_n984), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NOR4_X1   g578(.A1(new_n993), .A2(new_n994), .A3(new_n997), .A4(new_n1003), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n1003), .A2(new_n996), .B1(G2067), .B2(new_n752), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n991), .B(new_n1004), .C1(new_n982), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT126), .ZN(new_n1007));
  XNOR2_X1  g582(.A(G290), .B(G1986), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n997), .B(new_n1003), .C1(new_n1008), .C2(new_n982), .ZN(new_n1009));
  INV_X1    g584(.A(G1981), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n616), .A2(new_n619), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n611), .A2(new_n818), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n550), .B1(new_n613), .B2(new_n614), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n617), .A2(new_n618), .ZN(new_n1014));
  OAI21_X1  g589(.A(G1981), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1011), .A2(KEYINPUT49), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT49), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1011), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT113), .B(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n803), .B2(new_n804), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1021), .B2(new_n980), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n805), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n981), .B1(new_n1025), .B2(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g601(.A(G2090), .ZN(new_n1027));
  NOR4_X1   g602(.A1(G164), .A2(KEYINPUT111), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1026), .B(new_n1027), .C1(new_n1028), .C2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n805), .A2(KEYINPUT45), .A3(new_n1024), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n978), .A2(new_n1033), .A3(new_n980), .ZN(new_n1034));
  INV_X1    g609(.A(G1971), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT112), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  NAND4_X1  g615(.A1(G303), .A2(new_n1040), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G303), .A2(G8), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1037), .A2(new_n1045), .A3(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1021), .A2(new_n980), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1020), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1016), .A2(new_n1017), .A3(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n605), .B(G1976), .C1(new_n606), .C2(new_n550), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(KEYINPUT114), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1022), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1022), .B2(new_n1051), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n609), .A2(new_n1052), .A3(new_n818), .A4(new_n610), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1050), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1023), .B1(new_n1046), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT116), .B(KEYINPUT63), .ZN(new_n1061));
  INV_X1    g636(.A(G2084), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1026), .B(new_n1062), .C1(new_n1028), .C2(new_n1031), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1034), .A2(new_n729), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1020), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1065), .A2(KEYINPUT115), .A3(G168), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT115), .B1(new_n1065), .B2(G168), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1045), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n981), .B1(new_n1025), .B2(new_n977), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1971), .B1(new_n1070), .B2(new_n1033), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n980), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT50), .B(G1384), .C1(new_n803), .C2(new_n804), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1072), .A2(G2090), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1048), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(new_n1058), .A3(new_n1046), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1061), .B1(new_n1068), .B2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1058), .A2(new_n1046), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1037), .A2(G8), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1069), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1079), .B(new_n1082), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1060), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1034), .B2(G2078), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1070), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1033), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n805), .A2(new_n1030), .A3(new_n1024), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT111), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1021), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1072), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G1961), .ZN(new_n1093));
  OAI21_X1  g668(.A(G171), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT122), .B1(new_n1092), .B2(G1961), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1026), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  INV_X1    g672(.A(G1961), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n978), .A2(KEYINPUT123), .A3(new_n1033), .A4(new_n980), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT53), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1070), .A2(new_n443), .A3(new_n1033), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n978), .A2(new_n1033), .A3(new_n980), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1104), .A2(KEYINPUT53), .A3(new_n1100), .A4(new_n443), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1095), .A2(new_n1099), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1094), .B1(new_n1106), .B2(G171), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT124), .ZN(new_n1110));
  INV_X1    g685(.A(G8), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1112));
  NOR2_X1   g687(.A1(G168), .A2(new_n1020), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(G168), .B2(new_n1020), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT121), .B1(new_n1065), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1116), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1092), .A2(new_n1062), .B1(new_n729), .B2(new_n1034), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n1020), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1114), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1113), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1106), .A2(G171), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1108), .B1(new_n1127), .B2(G301), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1077), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1107), .A2(new_n1130), .A3(new_n1108), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1110), .A2(new_n1125), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(G1341), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1047), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT118), .B(G1996), .Z(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n1034), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n567), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1138), .B(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n580), .A2(new_n583), .A3(KEYINPUT76), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT57), .B(new_n598), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n587), .A2(new_n589), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(new_n597), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT117), .B(new_n1145), .C1(new_n1146), .C2(new_n597), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1144), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(G1956), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT56), .B(G2072), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n978), .A2(new_n1033), .A3(new_n980), .A4(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1158), .A2(new_n1144), .A3(new_n1150), .A4(new_n1149), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1141), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1159), .A3(new_n1141), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1140), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1047), .A2(G2067), .ZN(new_n1164));
  INV_X1    g739(.A(G1348), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1096), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(new_n1167), .A3(KEYINPUT60), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1164), .ZN(new_n1169));
  OAI211_X1 g744(.A(KEYINPUT60), .B(new_n1169), .C1(new_n1092), .C2(G1348), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT120), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1171), .A3(new_n640), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1170), .A2(KEYINPUT120), .A3(new_n641), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1166), .A2(KEYINPUT60), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1159), .B1(new_n641), .B2(new_n1166), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1163), .A2(new_n1175), .B1(new_n1176), .B2(new_n1157), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1084), .B1(new_n1132), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT125), .B1(new_n1125), .B2(KEYINPUT62), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n1181));
  AOI211_X1 g756(.A(new_n1180), .B(new_n1181), .C1(new_n1122), .C2(new_n1124), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1122), .A2(new_n1181), .A3(new_n1124), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1077), .A2(new_n1094), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1179), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1007), .B(new_n1009), .C1(new_n1178), .C2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1125), .A2(KEYINPUT62), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1180), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1125), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1107), .A2(new_n1130), .A3(new_n1108), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1130), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1129), .A2(new_n1125), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1176), .A2(new_n1157), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1138), .B(KEYINPUT59), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1157), .A2(new_n1159), .A3(new_n1141), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1200), .B1(new_n1201), .B2(new_n1160), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1198), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1196), .A2(new_n1197), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1193), .A2(new_n1204), .A3(new_n1084), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1007), .B1(new_n1205), .B2(new_n1009), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1006), .B1(new_n1188), .B2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g782(.A1(new_n702), .A2(G319), .A3(new_n685), .ZN(new_n1209));
  NOR2_X1   g783(.A1(G229), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g784(.A(new_n905), .B(new_n1210), .C1(new_n973), .C2(new_n974), .ZN(G225));
  INV_X1    g785(.A(G225), .ZN(G308));
endmodule


