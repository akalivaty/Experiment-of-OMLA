

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;

  XNOR2_X1 U322 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n436) );
  XNOR2_X1 U323 ( .A(n359), .B(n341), .ZN(n342) );
  INV_X1 U324 ( .A(n576), .ZN(n548) );
  XOR2_X1 U325 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n290) );
  XNOR2_X1 U326 ( .A(n343), .B(n342), .ZN(n366) );
  INV_X1 U327 ( .A(KEYINPUT22), .ZN(n424) );
  XNOR2_X1 U328 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U329 ( .A(KEYINPUT101), .B(KEYINPUT36), .ZN(n345) );
  XNOR2_X1 U330 ( .A(n427), .B(n426), .ZN(n430) );
  XNOR2_X1 U331 ( .A(n570), .B(n345), .ZN(n485) );
  XNOR2_X1 U332 ( .A(n461), .B(KEYINPUT26), .ZN(n576) );
  XNOR2_X1 U333 ( .A(n437), .B(n436), .ZN(n454) );
  XOR2_X1 U334 ( .A(KEYINPUT104), .B(n494), .Z(n503) );
  XNOR2_X1 U335 ( .A(n455), .B(KEYINPUT124), .ZN(n456) );
  XNOR2_X1 U336 ( .A(n457), .B(n456), .ZN(G1350GAT) );
  XNOR2_X1 U337 ( .A(G57GAT), .B(G64GAT), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n291), .B(KEYINPUT13), .ZN(n347) );
  XOR2_X1 U339 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n293) );
  XNOR2_X1 U340 ( .A(G211GAT), .B(G78GAT), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U342 ( .A(n347), .B(n294), .Z(n296) );
  XOR2_X1 U343 ( .A(G8GAT), .B(G1GAT), .Z(n310) );
  XOR2_X1 U344 ( .A(G22GAT), .B(G155GAT), .Z(n420) );
  XNOR2_X1 U345 ( .A(n310), .B(n420), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U347 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n298) );
  NAND2_X1 U348 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U350 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U351 ( .A(G71GAT), .B(G127GAT), .Z(n302) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n303), .B(KEYINPUT12), .ZN(n304) );
  XOR2_X1 U355 ( .A(n305), .B(n304), .Z(n557) );
  INV_X1 U356 ( .A(n557), .ZN(n587) );
  INV_X1 U357 ( .A(KEYINPUT54), .ZN(n392) );
  XOR2_X1 U358 ( .A(G141GAT), .B(G197GAT), .Z(n307) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(G36GAT), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n323) );
  XOR2_X1 U361 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n309) );
  XNOR2_X1 U362 ( .A(G22GAT), .B(KEYINPUT30), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n314) );
  XOR2_X1 U364 ( .A(G50GAT), .B(G43GAT), .Z(n312) );
  XOR2_X1 U365 ( .A(G113GAT), .B(G15GAT), .Z(n451) );
  XNOR2_X1 U366 ( .A(n451), .B(n310), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U368 ( .A(n314), .B(n313), .Z(n316) );
  NAND2_X1 U369 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U371 ( .A(n317), .B(KEYINPUT70), .Z(n321) );
  XOR2_X1 U372 ( .A(G29GAT), .B(KEYINPUT7), .Z(n319) );
  XNOR2_X1 U373 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n333) );
  XNOR2_X1 U375 ( .A(n333), .B(KEYINPUT29), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X2 U377 ( .A(n323), .B(n322), .Z(n562) );
  INV_X1 U378 ( .A(KEYINPUT79), .ZN(n344) );
  XOR2_X1 U379 ( .A(G36GAT), .B(G218GAT), .Z(n382) );
  XNOR2_X1 U380 ( .A(G43GAT), .B(G190GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n324), .B(G134GAT), .ZN(n440) );
  XNOR2_X1 U382 ( .A(n440), .B(KEYINPUT10), .ZN(n325) );
  AND2_X1 U383 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  NAND2_X1 U384 ( .A1(n325), .A2(n327), .ZN(n331) );
  INV_X1 U385 ( .A(KEYINPUT10), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n440), .B(n326), .ZN(n329) );
  INV_X1 U387 ( .A(n327), .ZN(n328) );
  NAND2_X1 U388 ( .A1(n329), .A2(n328), .ZN(n330) );
  NAND2_X1 U389 ( .A1(n331), .A2(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n382), .B(n332), .Z(n335) );
  XOR2_X1 U391 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U392 ( .A(n333), .B(n419), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n343) );
  XOR2_X1 U394 ( .A(KEYINPUT74), .B(G92GAT), .Z(n337) );
  XNOR2_X1 U395 ( .A(G99GAT), .B(G85GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U397 ( .A(G106GAT), .B(n338), .Z(n359) );
  XOR2_X1 U398 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n340) );
  XNOR2_X1 U399 ( .A(KEYINPUT77), .B(KEYINPUT9), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n344), .B(n366), .ZN(n570) );
  NOR2_X1 U402 ( .A1(n587), .A2(n485), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n346), .B(n290), .ZN(n362) );
  XOR2_X1 U404 ( .A(n347), .B(G204GAT), .Z(n349) );
  XOR2_X1 U405 ( .A(G120GAT), .B(G71GAT), .Z(n444) );
  XNOR2_X1 U406 ( .A(G176GAT), .B(n444), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n355) );
  XOR2_X1 U408 ( .A(G78GAT), .B(G148GAT), .Z(n351) );
  XNOR2_X1 U409 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n428) );
  XOR2_X1 U411 ( .A(n428), .B(KEYINPUT31), .Z(n353) );
  NAND2_X1 U412 ( .A1(G230GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U414 ( .A(n355), .B(n354), .Z(n361) );
  XOR2_X1 U415 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n357) );
  XNOR2_X1 U416 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n583) );
  NAND2_X1 U420 ( .A1(n362), .A2(n583), .ZN(n363) );
  NOR2_X1 U421 ( .A1(n562), .A2(n363), .ZN(n365) );
  INV_X1 U422 ( .A(KEYINPUT113), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n372) );
  XOR2_X1 U424 ( .A(KEYINPUT41), .B(n583), .Z(n565) );
  INV_X1 U425 ( .A(n565), .ZN(n553) );
  NAND2_X1 U426 ( .A1(n562), .A2(n553), .ZN(n367) );
  XNOR2_X1 U427 ( .A(KEYINPUT46), .B(n367), .ZN(n368) );
  NAND2_X1 U428 ( .A1(n368), .A2(n587), .ZN(n369) );
  NOR2_X1 U429 ( .A1(n366), .A2(n369), .ZN(n370) );
  XOR2_X1 U430 ( .A(KEYINPUT47), .B(n370), .Z(n371) );
  NOR2_X1 U431 ( .A1(n372), .A2(n371), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n373), .B(KEYINPUT48), .ZN(n531) );
  XOR2_X1 U433 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n375) );
  XNOR2_X1 U434 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U436 ( .A(n376), .B(G183GAT), .Z(n378) );
  XNOR2_X1 U437 ( .A(G169GAT), .B(G176GAT), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n450) );
  XOR2_X1 U439 ( .A(KEYINPUT97), .B(G92GAT), .Z(n380) );
  XNOR2_X1 U440 ( .A(G8GAT), .B(G190GAT), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U442 ( .A(n382), .B(n381), .Z(n384) );
  NAND2_X1 U443 ( .A1(G226GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U445 ( .A(n385), .B(KEYINPUT96), .Z(n389) );
  XOR2_X1 U446 ( .A(G204GAT), .B(G211GAT), .Z(n387) );
  XNOR2_X1 U447 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n432) );
  XNOR2_X1 U449 ( .A(n432), .B(G64GAT), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n450), .B(n390), .ZN(n497) );
  INV_X1 U452 ( .A(n497), .ZN(n521) );
  NOR2_X1 U453 ( .A1(n531), .A2(n521), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n574) );
  XOR2_X1 U455 ( .A(KEYINPUT94), .B(KEYINPUT1), .Z(n394) );
  XNOR2_X1 U456 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n415) );
  XOR2_X1 U458 ( .A(G57GAT), .B(G155GAT), .Z(n396) );
  XNOR2_X1 U459 ( .A(G120GAT), .B(G148GAT), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U461 ( .A(KEYINPUT92), .B(KEYINPUT95), .Z(n398) );
  XNOR2_X1 U462 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U464 ( .A(n400), .B(n399), .Z(n413) );
  XOR2_X1 U465 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n402) );
  XNOR2_X1 U466 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n431) );
  XOR2_X1 U468 ( .A(n431), .B(KEYINPUT93), .Z(n404) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n411) );
  XOR2_X1 U471 ( .A(KEYINPUT77), .B(G85GAT), .Z(n406) );
  XNOR2_X1 U472 ( .A(G113GAT), .B(G134GAT), .ZN(n405) );
  XNOR2_X1 U473 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U474 ( .A(n407), .B(G162GAT), .Z(n409) );
  XOR2_X1 U475 ( .A(KEYINPUT0), .B(G127GAT), .Z(n445) );
  XNOR2_X1 U476 ( .A(G29GAT), .B(n445), .ZN(n408) );
  XNOR2_X1 U477 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U480 ( .A(n415), .B(n414), .Z(n518) );
  XOR2_X1 U481 ( .A(KEYINPUT91), .B(KEYINPUT89), .Z(n417) );
  XNOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U484 ( .A(G106GAT), .B(G218GAT), .Z(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U487 ( .A(n423), .B(n422), .Z(n427) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n428), .B(KEYINPUT90), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U491 ( .A(n432), .B(n431), .Z(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n464) );
  NAND2_X1 U493 ( .A1(n518), .A2(n464), .ZN(n435) );
  OR2_X1 U494 ( .A1(n574), .A2(n435), .ZN(n437) );
  XOR2_X1 U495 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n439) );
  XNOR2_X1 U497 ( .A(G99GAT), .B(KEYINPUT64), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n449) );
  XOR2_X1 U501 ( .A(n445), .B(n444), .Z(n447) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U504 ( .A(n449), .B(n448), .Z(n453) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U506 ( .A(n453), .B(n452), .Z(n523) );
  INV_X1 U507 ( .A(n523), .ZN(n534) );
  NAND2_X1 U508 ( .A1(n454), .A2(n534), .ZN(n569) );
  NOR2_X1 U509 ( .A1(n587), .A2(n569), .ZN(n457) );
  INV_X1 U510 ( .A(G183GAT), .ZN(n455) );
  XNOR2_X1 U511 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U512 ( .A(n497), .B(KEYINPUT27), .ZN(n462) );
  INV_X1 U513 ( .A(n518), .ZN(n575) );
  NAND2_X1 U514 ( .A1(n462), .A2(n575), .ZN(n530) );
  XNOR2_X1 U515 ( .A(n523), .B(KEYINPUT87), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n530), .A2(n458), .ZN(n460) );
  XNOR2_X1 U517 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n459) );
  XOR2_X1 U518 ( .A(n459), .B(n464), .Z(n502) );
  INV_X1 U519 ( .A(n502), .ZN(n533) );
  NAND2_X1 U520 ( .A1(n460), .A2(n533), .ZN(n470) );
  NOR2_X1 U521 ( .A1(n464), .A2(n534), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n462), .A2(n576), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n534), .A2(n497), .ZN(n463) );
  NAND2_X1 U524 ( .A1(n464), .A2(n463), .ZN(n465) );
  XOR2_X1 U525 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  NAND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n468), .A2(n518), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT98), .ZN(n487) );
  XNOR2_X1 U530 ( .A(KEYINPUT82), .B(KEYINPUT16), .ZN(n473) );
  NOR2_X1 U531 ( .A1(n587), .A2(n570), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n474) );
  AND2_X1 U533 ( .A1(n487), .A2(n474), .ZN(n506) );
  NAND2_X1 U534 ( .A1(n583), .A2(n562), .ZN(n475) );
  XOR2_X1 U535 ( .A(KEYINPUT76), .B(n475), .Z(n491) );
  NAND2_X1 U536 ( .A1(n506), .A2(n491), .ZN(n476) );
  XNOR2_X1 U537 ( .A(KEYINPUT99), .B(n476), .ZN(n483) );
  NAND2_X1 U538 ( .A1(n483), .A2(n575), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U540 ( .A1(n497), .A2(n483), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n479), .B(KEYINPUT100), .ZN(n480) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(n480), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT35), .Z(n482) );
  NAND2_X1 U544 ( .A1(n483), .A2(n534), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(G1326GAT) );
  NAND2_X1 U546 ( .A1(n483), .A2(n502), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n484), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .Z(n496) );
  XOR2_X1 U549 ( .A(KEYINPUT105), .B(KEYINPUT38), .Z(n493) );
  NOR2_X1 U550 ( .A1(n557), .A2(n485), .ZN(n486) );
  NAND2_X1 U551 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U552 ( .A(KEYINPUT102), .B(n488), .ZN(n490) );
  XOR2_X1 U553 ( .A(KEYINPUT103), .B(KEYINPUT37), .Z(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(n516) );
  NAND2_X1 U555 ( .A1(n516), .A2(n491), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  NAND2_X1 U557 ( .A1(n503), .A2(n575), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n497), .A2(n503), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n500) );
  NAND2_X1 U562 ( .A1(n503), .A2(n534), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U564 ( .A(n501), .B(G43GAT), .Z(G1330GAT) );
  XOR2_X1 U565 ( .A(G50GAT), .B(KEYINPUT107), .Z(n505) );
  NAND2_X1 U566 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  NOR2_X1 U568 ( .A1(n562), .A2(n565), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n506), .A2(n517), .ZN(n512) );
  NOR2_X1 U570 ( .A1(n518), .A2(n512), .ZN(n507) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n507), .Z(n508) );
  XNOR2_X1 U572 ( .A(KEYINPUT42), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U573 ( .A1(n521), .A2(n512), .ZN(n509) );
  XOR2_X1 U574 ( .A(KEYINPUT108), .B(n509), .Z(n510) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(n510), .ZN(G1333GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n512), .ZN(n511) );
  XOR2_X1 U577 ( .A(G71GAT), .B(n511), .Z(G1334GAT) );
  NOR2_X1 U578 ( .A1(n533), .A2(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U581 ( .A(G78GAT), .B(n515), .Z(G1335GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n527) );
  NOR2_X1 U583 ( .A1(n518), .A2(n527), .ZN(n519) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n519), .Z(n520) );
  XNOR2_X1 U585 ( .A(KEYINPUT110), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n527), .ZN(n522) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n527), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n526), .ZN(G1338GAT) );
  NOR2_X1 U592 ( .A1(n533), .A2(n527), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n538) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT114), .B(n532), .Z(n549) );
  NAND2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n549), .A2(n535), .ZN(n536) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(n536), .Z(n544) );
  NAND2_X1 U601 ( .A1(n562), .A2(n544), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U604 ( .A1(n544), .A2(n553), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n542) );
  NAND2_X1 U607 ( .A1(n544), .A2(n557), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U611 ( .A1(n544), .A2(n570), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n547), .ZN(G1343GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n551) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n560), .A2(n562), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  NAND2_X1 U620 ( .A1(n560), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  XOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n366), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U628 ( .A(n562), .ZN(n578) );
  NOR2_X1 U629 ( .A1(n578), .A2(n569), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1348GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n569), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(n568), .ZN(G1349GAT) );
  INV_X1 U636 ( .A(n569), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT58), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n573), .ZN(G1351GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n589) );
  NOR2_X1 U642 ( .A1(n589), .A2(n578), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n589), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(n586), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n589), .ZN(n588) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n588), .Z(G1354GAT) );
  NOR2_X1 U653 ( .A1(n485), .A2(n589), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

