

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771;

  NOR2_X1 U379 ( .A1(n565), .A2(n564), .ZN(n678) );
  XOR2_X1 U380 ( .A(G119), .B(G110), .Z(n509) );
  INV_X1 U381 ( .A(n405), .ZN(n480) );
  XNOR2_X1 U382 ( .A(n551), .B(n356), .ZN(n380) );
  XOR2_X1 U383 ( .A(n550), .B(KEYINPUT40), .Z(n356) );
  XOR2_X1 U384 ( .A(G131), .B(KEYINPUT127), .Z(n357) );
  XOR2_X1 U385 ( .A(n522), .B(KEYINPUT68), .Z(n358) );
  NOR2_X1 U386 ( .A1(n608), .A2(n724), .ZN(n378) );
  NOR2_X1 U387 ( .A1(n725), .A2(n564), .ZN(n369) );
  NOR2_X1 U388 ( .A1(n594), .A2(n610), .ZN(n595) );
  XNOR2_X2 U389 ( .A(n358), .B(n487), .ZN(n758) );
  XNOR2_X2 U390 ( .A(n505), .B(n536), .ZN(n759) );
  INV_X1 U391 ( .A(n406), .ZN(n479) );
  INV_X1 U392 ( .A(KEYINPUT4), .ZN(n359) );
  XNOR2_X2 U393 ( .A(G134), .B(G131), .ZN(n522) );
  XNOR2_X1 U394 ( .A(n369), .B(KEYINPUT42), .ZN(n771) );
  NAND2_X1 U395 ( .A1(n385), .A2(n384), .ZN(n564) );
  XNOR2_X1 U396 ( .A(n549), .B(KEYINPUT39), .ZN(n584) );
  XNOR2_X1 U397 ( .A(n595), .B(KEYINPUT33), .ZN(n724) );
  AND2_X1 U398 ( .A1(n546), .A2(n547), .ZN(n548) );
  XNOR2_X1 U399 ( .A(n521), .B(n520), .ZN(n392) );
  NAND2_X2 U400 ( .A1(n449), .A2(n445), .ZN(n605) );
  XOR2_X1 U401 ( .A(KEYINPUT121), .B(n654), .Z(n655) );
  XNOR2_X1 U402 ( .A(KEYINPUT77), .B(n361), .ZN(n526) );
  NAND2_X1 U403 ( .A1(n458), .A2(KEYINPUT82), .ZN(n367) );
  XNOR2_X1 U404 ( .A(G902), .B(KEYINPUT15), .ZN(n629) );
  NOR2_X1 U405 ( .A1(n422), .A2(n367), .ZN(n419) );
  AND2_X2 U406 ( .A1(n628), .A2(n745), .ZN(n422) );
  XNOR2_X2 U407 ( .A(n486), .B(n359), .ZN(n487) );
  XNOR2_X1 U408 ( .A(n380), .B(n357), .ZN(G33) );
  XNOR2_X1 U409 ( .A(n411), .B(KEYINPUT45), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n411), .B(KEYINPUT45), .ZN(n745) );
  BUF_X1 U411 ( .A(n700), .Z(n426) );
  XNOR2_X2 U412 ( .A(G107), .B(G116), .ZN(n406) );
  XNOR2_X2 U413 ( .A(n400), .B(n539), .ZN(n368) );
  XNOR2_X2 U414 ( .A(n758), .B(G146), .ZN(n400) );
  XNOR2_X1 U415 ( .A(n605), .B(KEYINPUT1), .ZN(n693) );
  XNOR2_X1 U416 ( .A(n700), .B(n375), .ZN(n594) );
  AND2_X1 U417 ( .A1(n597), .A2(n697), .ZN(n598) );
  NAND2_X1 U418 ( .A1(n370), .A2(n697), .ZN(n540) );
  NAND2_X1 U419 ( .A1(n504), .A2(n590), .ZN(n370) );
  INV_X1 U420 ( .A(KEYINPUT78), .ZN(n454) );
  NAND2_X1 U421 ( .A1(n494), .A2(G214), .ZN(n709) );
  NAND2_X1 U422 ( .A1(n426), .A2(KEYINPUT28), .ZN(n387) );
  NAND2_X1 U423 ( .A1(n390), .A2(n389), .ZN(n388) );
  NOR2_X1 U424 ( .A1(n426), .A2(KEYINPUT28), .ZN(n389) );
  INV_X1 U425 ( .A(KEYINPUT0), .ZN(n418) );
  XNOR2_X1 U426 ( .A(n434), .B(n433), .ZN(n510) );
  INV_X1 U427 ( .A(KEYINPUT8), .ZN(n433) );
  NAND2_X1 U428 ( .A1(n761), .A2(G234), .ZN(n434) );
  XOR2_X1 U429 ( .A(KEYINPUT24), .B(KEYINPUT72), .Z(n507) );
  XNOR2_X1 U430 ( .A(n477), .B(n476), .ZN(n436) );
  XNOR2_X1 U431 ( .A(G134), .B(G122), .ZN(n476) );
  XOR2_X1 U432 ( .A(G137), .B(G140), .Z(n536) );
  XOR2_X1 U433 ( .A(G110), .B(G107), .Z(n535) );
  XNOR2_X1 U434 ( .A(G101), .B(G104), .ZN(n534) );
  INV_X1 U435 ( .A(KEYINPUT64), .ZN(n443) );
  INV_X1 U436 ( .A(KEYINPUT100), .ZN(n579) );
  XNOR2_X1 U437 ( .A(n471), .B(n427), .ZN(n569) );
  XNOR2_X1 U438 ( .A(n472), .B(n428), .ZN(n427) );
  INV_X1 U439 ( .A(G475), .ZN(n428) );
  AND2_X1 U440 ( .A1(n451), .A2(n450), .ZN(n449) );
  NAND2_X1 U441 ( .A1(n448), .A2(n447), .ZN(n446) );
  INV_X1 U442 ( .A(n594), .ZN(n374) );
  INV_X2 U443 ( .A(G953), .ZN(n761) );
  AND2_X1 U444 ( .A1(n396), .A2(n401), .ZN(n395) );
  INV_X1 U445 ( .A(KEYINPUT47), .ZN(n431) );
  NAND2_X1 U446 ( .A1(n394), .A2(KEYINPUT47), .ZN(n393) );
  INV_X1 U447 ( .A(KEYINPUT2), .ZN(n458) );
  INV_X1 U448 ( .A(G237), .ZN(n490) );
  XNOR2_X1 U449 ( .A(n371), .B(KEYINPUT90), .ZN(n590) );
  NAND2_X1 U450 ( .A1(n372), .A2(n761), .ZN(n371) );
  XNOR2_X1 U451 ( .A(KEYINPUT5), .B(G137), .ZN(n527) );
  XNOR2_X1 U452 ( .A(G119), .B(G116), .ZN(n523) );
  XOR2_X1 U453 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n467) );
  XNOR2_X1 U454 ( .A(G131), .B(G113), .ZN(n466) );
  XNOR2_X1 U455 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n463) );
  XNOR2_X1 U456 ( .A(G143), .B(G140), .ZN(n461) );
  XNOR2_X1 U457 ( .A(n437), .B(n481), .ZN(n752) );
  XNOR2_X1 U458 ( .A(n438), .B(n525), .ZN(n437) );
  NAND2_X1 U459 ( .A1(G234), .A2(G237), .ZN(n499) );
  XNOR2_X1 U460 ( .A(n373), .B(KEYINPUT89), .ZN(n500) );
  INV_X1 U461 ( .A(KEYINPUT14), .ZN(n373) );
  INV_X1 U462 ( .A(G469), .ZN(n448) );
  NAND2_X1 U463 ( .A1(G902), .A2(G469), .ZN(n450) );
  XOR2_X1 U464 ( .A(G146), .B(G125), .Z(n485) );
  NAND2_X1 U465 ( .A1(n363), .A2(n452), .ZN(n691) );
  XNOR2_X1 U466 ( .A(n496), .B(n495), .ZN(n725) );
  NOR2_X1 U467 ( .A1(n391), .A2(n712), .ZN(n496) );
  AND2_X1 U468 ( .A1(n680), .A2(n555), .ZN(n576) );
  AND2_X1 U469 ( .A1(n388), .A2(n386), .ZN(n385) );
  AND2_X1 U470 ( .A1(n387), .A2(n605), .ZN(n386) );
  XNOR2_X1 U471 ( .A(n383), .B(n513), .ZN(n654) );
  XNOR2_X1 U472 ( .A(n759), .B(n508), .ZN(n383) );
  XNOR2_X1 U473 ( .A(n475), .B(n435), .ZN(n740) );
  XNOR2_X1 U474 ( .A(n436), .B(n406), .ZN(n435) );
  XNOR2_X1 U475 ( .A(n642), .B(n641), .ZN(n643) );
  AND2_X1 U476 ( .A1(n634), .A2(G953), .ZN(n744) );
  NOR2_X1 U477 ( .A1(n582), .A2(n570), .ZN(n583) );
  XNOR2_X1 U478 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U479 ( .A(n579), .B(KEYINPUT43), .ZN(n580) );
  NAND2_X1 U480 ( .A1(n377), .A2(n596), .ZN(n376) );
  XNOR2_X1 U481 ( .A(n378), .B(KEYINPUT34), .ZN(n377) );
  INV_X1 U482 ( .A(KEYINPUT65), .ZN(n429) );
  NAND2_X1 U483 ( .A1(n601), .A2(n600), .ZN(n659) );
  OR2_X1 U484 ( .A1(G953), .A2(G237), .ZN(n361) );
  INV_X1 U485 ( .A(n401), .ZN(n677) );
  AND2_X1 U486 ( .A1(n399), .A2(n659), .ZN(n362) );
  AND2_X1 U487 ( .A1(n456), .A2(n424), .ZN(n363) );
  AND2_X1 U488 ( .A1(n596), .A2(n570), .ZN(n364) );
  NOR2_X1 U489 ( .A1(n740), .A2(G902), .ZN(n365) );
  INV_X1 U490 ( .A(G902), .ZN(n447) );
  BUF_X1 U491 ( .A(n693), .Z(n425) );
  INV_X1 U492 ( .A(n425), .ZN(n442) );
  AND2_X1 U493 ( .A1(n630), .A2(n458), .ZN(n366) );
  NAND2_X1 U494 ( .A1(n761), .A2(G224), .ZN(n483) );
  NAND2_X1 U495 ( .A1(n368), .A2(G469), .ZN(n451) );
  OR2_X1 U496 ( .A1(n368), .A2(n446), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n368), .B(n735), .ZN(n736) );
  INV_X1 U498 ( .A(n771), .ZN(n379) );
  INV_X1 U499 ( .A(n723), .ZN(n372) );
  NOR2_X2 U500 ( .A1(n618), .A2(n374), .ZN(n616) );
  INV_X1 U501 ( .A(KEYINPUT6), .ZN(n375) );
  XNOR2_X2 U502 ( .A(G122), .B(G104), .ZN(n405) );
  XNOR2_X2 U503 ( .A(n376), .B(KEYINPUT35), .ZN(n416) );
  NAND2_X1 U504 ( .A1(n380), .A2(n379), .ZN(n553) );
  XNOR2_X1 U505 ( .A(n381), .B(n398), .ZN(n414) );
  NAND2_X1 U506 ( .A1(n382), .A2(n362), .ZN(n381) );
  NAND2_X1 U507 ( .A1(n416), .A2(KEYINPUT44), .ZN(n382) );
  XNOR2_X2 U508 ( .A(n462), .B(KEYINPUT10), .ZN(n505) );
  NAND2_X1 U509 ( .A1(n392), .A2(KEYINPUT28), .ZN(n384) );
  INV_X1 U510 ( .A(n392), .ZN(n390) );
  NOR2_X1 U511 ( .A1(n602), .A2(n391), .ZN(n714) );
  NAND2_X1 U512 ( .A1(n710), .A2(n709), .ZN(n391) );
  NOR2_X1 U513 ( .A1(n594), .A2(n392), .ZN(n555) );
  NAND2_X1 U514 ( .A1(n395), .A2(n393), .ZN(n571) );
  NAND2_X1 U515 ( .A1(n678), .A2(n567), .ZN(n394) );
  NAND2_X1 U516 ( .A1(n678), .A2(n397), .ZN(n396) );
  AND2_X1 U517 ( .A1(n432), .A2(n431), .ZN(n397) );
  INV_X1 U518 ( .A(KEYINPUT84), .ZN(n398) );
  OR2_X2 U519 ( .A1(n614), .A2(n602), .ZN(n399) );
  XNOR2_X1 U520 ( .A(n531), .B(n400), .ZN(n631) );
  NAND2_X1 U521 ( .A1(n548), .A2(n364), .ZN(n401) );
  BUF_X1 U522 ( .A(n752), .Z(n402) );
  INV_X1 U523 ( .A(n455), .ZN(n403) );
  XNOR2_X1 U524 ( .A(n631), .B(KEYINPUT62), .ZN(n632) );
  OR2_X2 U525 ( .A1(n700), .A2(n543), .ZN(n545) );
  XNOR2_X2 U526 ( .A(G146), .B(G125), .ZN(n462) );
  XNOR2_X1 U527 ( .A(n575), .B(n574), .ZN(n586) );
  XNOR2_X1 U528 ( .A(n402), .B(n489), .ZN(n404) );
  NAND2_X1 U529 ( .A1(n480), .A2(n479), .ZN(n407) );
  NAND2_X1 U530 ( .A1(n405), .A2(n406), .ZN(n408) );
  NAND2_X1 U531 ( .A1(n407), .A2(n408), .ZN(n438) );
  XNOR2_X1 U532 ( .A(n752), .B(n489), .ZN(n649) );
  XNOR2_X1 U533 ( .A(n622), .B(n621), .ZN(n413) );
  XNOR2_X1 U534 ( .A(n430), .B(n429), .ZN(n620) );
  XNOR2_X2 U535 ( .A(n617), .B(KEYINPUT32), .ZN(n770) );
  NOR2_X2 U536 ( .A1(n618), .A2(n441), .ZN(n430) );
  BUF_X1 U537 ( .A(n684), .Z(n409) );
  XNOR2_X1 U538 ( .A(n562), .B(KEYINPUT19), .ZN(n593) );
  XNOR2_X2 U539 ( .A(n410), .B(KEYINPUT86), .ZN(n562) );
  NAND2_X2 U540 ( .A1(n554), .A2(n709), .ZN(n410) );
  XNOR2_X2 U541 ( .A(n492), .B(n491), .ZN(n554) );
  NAND2_X1 U542 ( .A1(n593), .A2(n592), .ZN(n415) );
  NAND2_X1 U543 ( .A1(n414), .A2(n412), .ZN(n411) );
  NAND2_X1 U544 ( .A1(n413), .A2(n624), .ZN(n412) );
  XNOR2_X2 U545 ( .A(n415), .B(n418), .ZN(n609) );
  INV_X1 U546 ( .A(n416), .ZN(n417) );
  NAND2_X1 U547 ( .A1(n416), .A2(n623), .ZN(n624) );
  XNOR2_X1 U548 ( .A(n417), .B(G122), .ZN(G24) );
  INV_X1 U549 ( .A(n609), .ZN(n608) );
  NOR2_X1 U550 ( .A1(n420), .A2(n419), .ZN(n423) );
  NAND2_X1 U551 ( .A1(n421), .A2(n626), .ZN(n420) );
  NAND2_X1 U552 ( .A1(n422), .A2(n366), .ZN(n421) );
  NAND2_X1 U553 ( .A1(n423), .A2(n691), .ZN(n444) );
  NAND2_X1 U554 ( .A1(n455), .A2(KEYINPUT78), .ZN(n424) );
  NAND2_X1 U555 ( .A1(n586), .A2(n585), .ZN(n760) );
  XNOR2_X1 U556 ( .A(n505), .B(n463), .ZN(n464) );
  XNOR2_X1 U557 ( .A(n470), .B(n469), .ZN(n642) );
  XNOR2_X1 U558 ( .A(n602), .B(n566), .ZN(n432) );
  NAND2_X1 U559 ( .A1(n510), .A2(G217), .ZN(n474) );
  OR2_X2 U560 ( .A1(n631), .A2(G902), .ZN(n533) );
  INV_X1 U561 ( .A(n760), .ZN(n688) );
  NAND2_X1 U562 ( .A1(n457), .A2(KEYINPUT78), .ZN(n456) );
  XNOR2_X2 U563 ( .A(n440), .B(n439), .ZN(n525) );
  XNOR2_X2 U564 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n439) );
  XNOR2_X2 U565 ( .A(G113), .B(G101), .ZN(n440) );
  NAND2_X1 U566 ( .A1(n442), .A2(n426), .ZN(n441) );
  XNOR2_X2 U567 ( .A(n599), .B(KEYINPUT22), .ZN(n618) );
  XNOR2_X2 U568 ( .A(n444), .B(n443), .ZN(n734) );
  XNOR2_X2 U569 ( .A(G143), .B(G128), .ZN(n486) );
  INV_X1 U570 ( .A(n625), .ZN(n457) );
  NAND2_X1 U571 ( .A1(n625), .A2(n453), .ZN(n452) );
  AND2_X1 U572 ( .A1(n360), .A2(n454), .ZN(n453) );
  INV_X1 U573 ( .A(n360), .ZN(n455) );
  XNOR2_X1 U574 ( .A(n742), .B(n741), .ZN(n743) );
  BUF_X1 U575 ( .A(n734), .Z(n739) );
  XNOR2_X1 U576 ( .A(n740), .B(KEYINPUT120), .ZN(n741) );
  XOR2_X1 U577 ( .A(n467), .B(n466), .Z(n459) );
  AND2_X1 U578 ( .A1(G227), .A2(n761), .ZN(n460) );
  INV_X1 U579 ( .A(n696), .ZN(n697) );
  INV_X1 U580 ( .A(KEYINPUT69), .ZN(n520) );
  XNOR2_X1 U581 ( .A(n468), .B(n459), .ZN(n469) );
  XNOR2_X1 U582 ( .A(n538), .B(n537), .ZN(n539) );
  AND2_X1 U583 ( .A1(n569), .A2(n559), .ZN(n680) );
  XNOR2_X1 U584 ( .A(n480), .B(n461), .ZN(n465) );
  XOR2_X1 U585 ( .A(n465), .B(n464), .Z(n470) );
  NAND2_X1 U586 ( .A1(G214), .A2(n526), .ZN(n468) );
  NOR2_X1 U587 ( .A1(G902), .A2(n642), .ZN(n471) );
  INV_X1 U588 ( .A(KEYINPUT13), .ZN(n472) );
  XNOR2_X1 U589 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n477) );
  XNOR2_X1 U590 ( .A(n486), .B(KEYINPUT96), .ZN(n473) );
  XNOR2_X1 U591 ( .A(n474), .B(n473), .ZN(n475) );
  INV_X1 U592 ( .A(G478), .ZN(n478) );
  XNOR2_X1 U593 ( .A(n365), .B(n478), .ZN(n568) );
  NOR2_X1 U594 ( .A1(n569), .A2(n568), .ZN(n597) );
  INV_X1 U595 ( .A(n597), .ZN(n712) );
  XOR2_X1 U596 ( .A(KEYINPUT16), .B(n509), .Z(n481) );
  XNOR2_X2 U597 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n482) );
  XNOR2_X1 U598 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U599 ( .A(n485), .B(n484), .ZN(n488) );
  XNOR2_X1 U600 ( .A(n488), .B(n487), .ZN(n489) );
  NAND2_X1 U601 ( .A1(n649), .A2(n629), .ZN(n492) );
  NAND2_X1 U602 ( .A1(n447), .A2(n490), .ZN(n494) );
  AND2_X1 U603 ( .A1(n494), .A2(G210), .ZN(n491) );
  BUF_X1 U604 ( .A(n554), .Z(n570) );
  XNOR2_X1 U605 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n493) );
  XNOR2_X1 U606 ( .A(n570), .B(n493), .ZN(n710) );
  XOR2_X1 U607 ( .A(KEYINPUT103), .B(KEYINPUT41), .Z(n495) );
  NAND2_X1 U608 ( .A1(n629), .A2(G234), .ZN(n497) );
  XNOR2_X1 U609 ( .A(n497), .B(KEYINPUT20), .ZN(n514) );
  NAND2_X1 U610 ( .A1(n514), .A2(G221), .ZN(n498) );
  XNOR2_X1 U611 ( .A(KEYINPUT21), .B(n498), .ZN(n696) );
  XNOR2_X1 U612 ( .A(n500), .B(n499), .ZN(n503) );
  NAND2_X1 U613 ( .A1(G902), .A2(n503), .ZN(n587) );
  NOR2_X1 U614 ( .A1(G900), .A2(n587), .ZN(n501) );
  NAND2_X1 U615 ( .A1(G953), .A2(n501), .ZN(n502) );
  XNOR2_X1 U616 ( .A(KEYINPUT98), .B(n502), .ZN(n504) );
  NAND2_X1 U617 ( .A1(G952), .A2(n503), .ZN(n723) );
  XOR2_X1 U618 ( .A(KEYINPUT70), .B(n540), .Z(n519) );
  XNOR2_X1 U619 ( .A(G128), .B(KEYINPUT92), .ZN(n506) );
  XNOR2_X1 U620 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U621 ( .A(n509), .B(KEYINPUT23), .Z(n512) );
  NAND2_X1 U622 ( .A1(G221), .A2(n510), .ZN(n511) );
  XNOR2_X1 U623 ( .A(n512), .B(n511), .ZN(n513) );
  NOR2_X1 U624 ( .A1(n654), .A2(G902), .ZN(n518) );
  XOR2_X1 U625 ( .A(KEYINPUT80), .B(KEYINPUT25), .Z(n516) );
  NAND2_X1 U626 ( .A1(n514), .A2(G217), .ZN(n515) );
  XNOR2_X1 U627 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X2 U628 ( .A(n518), .B(n517), .ZN(n619) );
  NAND2_X1 U629 ( .A1(n519), .A2(n619), .ZN(n521) );
  XNOR2_X1 U630 ( .A(n523), .B(KEYINPUT93), .ZN(n524) );
  XNOR2_X1 U631 ( .A(n525), .B(n524), .ZN(n530) );
  NAND2_X1 U632 ( .A1(n526), .A2(G210), .ZN(n528) );
  XNOR2_X1 U633 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U634 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U635 ( .A(KEYINPUT73), .B(G472), .ZN(n532) );
  XNOR2_X2 U636 ( .A(n533), .B(n532), .ZN(n700) );
  XNOR2_X1 U637 ( .A(n535), .B(n534), .ZN(n538) );
  XNOR2_X1 U638 ( .A(n536), .B(n460), .ZN(n537) );
  NOR2_X1 U639 ( .A1(n619), .A2(n540), .ZN(n541) );
  NAND2_X1 U640 ( .A1(n605), .A2(n541), .ZN(n542) );
  XNOR2_X1 U641 ( .A(n542), .B(KEYINPUT79), .ZN(n547) );
  INV_X1 U642 ( .A(n709), .ZN(n543) );
  INV_X1 U643 ( .A(KEYINPUT30), .ZN(n544) );
  XNOR2_X1 U644 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U645 ( .A1(n548), .A2(n710), .ZN(n549) );
  INV_X1 U646 ( .A(n568), .ZN(n559) );
  NAND2_X1 U647 ( .A1(n584), .A2(n680), .ZN(n551) );
  INV_X1 U648 ( .A(KEYINPUT102), .ZN(n550) );
  INV_X1 U649 ( .A(KEYINPUT46), .ZN(n552) );
  XNOR2_X1 U650 ( .A(n553), .B(n552), .ZN(n573) );
  INV_X1 U651 ( .A(n576), .ZN(n556) );
  NOR2_X1 U652 ( .A1(n562), .A2(n556), .ZN(n557) );
  XOR2_X1 U653 ( .A(KEYINPUT36), .B(n557), .Z(n558) );
  NOR2_X1 U654 ( .A1(n558), .A2(n442), .ZN(n686) );
  INV_X1 U655 ( .A(KEYINPUT74), .ZN(n566) );
  NOR2_X1 U656 ( .A1(n569), .A2(n559), .ZN(n561) );
  INV_X1 U657 ( .A(KEYINPUT97), .ZN(n560) );
  XNOR2_X1 U658 ( .A(n561), .B(n560), .ZN(n683) );
  NOR2_X1 U659 ( .A1(n680), .A2(n683), .ZN(n602) );
  BUF_X1 U660 ( .A(n593), .Z(n563) );
  INV_X1 U661 ( .A(n563), .ZN(n565) );
  NOR2_X1 U662 ( .A1(n602), .A2(n566), .ZN(n567) );
  AND2_X1 U663 ( .A1(n569), .A2(n568), .ZN(n596) );
  NOR2_X1 U664 ( .A1(n686), .A2(n571), .ZN(n572) );
  NAND2_X1 U665 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U666 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n574) );
  NAND2_X1 U667 ( .A1(n576), .A2(n709), .ZN(n577) );
  XNOR2_X1 U668 ( .A(KEYINPUT99), .B(n577), .ZN(n578) );
  NAND2_X1 U669 ( .A1(n578), .A2(n442), .ZN(n581) );
  XNOR2_X1 U670 ( .A(n583), .B(KEYINPUT101), .ZN(n769) );
  NAND2_X1 U671 ( .A1(n683), .A2(n584), .ZN(n638) );
  AND2_X1 U672 ( .A1(n769), .A2(n638), .ZN(n585) );
  AND2_X2 U673 ( .A1(KEYINPUT2), .A2(n688), .ZN(n625) );
  NOR2_X1 U674 ( .A1(G898), .A2(n761), .ZN(n754) );
  INV_X1 U675 ( .A(n587), .ZN(n588) );
  NAND2_X1 U676 ( .A1(n754), .A2(n588), .ZN(n589) );
  XOR2_X1 U677 ( .A(KEYINPUT91), .B(n589), .Z(n591) );
  NAND2_X1 U678 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U679 ( .A1(n696), .A2(n619), .ZN(n694) );
  NAND2_X1 U680 ( .A1(n694), .A2(n693), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n609), .A2(n598), .ZN(n599) );
  BUF_X1 U682 ( .A(n616), .Z(n601) );
  NOR2_X1 U683 ( .A1(n425), .A2(n619), .ZN(n600) );
  INV_X1 U684 ( .A(n694), .ZN(n604) );
  INV_X1 U685 ( .A(n426), .ZN(n603) );
  NOR2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n668) );
  BUF_X1 U689 ( .A(n609), .Z(n612) );
  OR2_X1 U690 ( .A1(n426), .A2(n610), .ZN(n705) );
  INV_X1 U691 ( .A(n705), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U693 ( .A(KEYINPUT31), .B(n613), .ZN(n684) );
  NOR2_X1 U694 ( .A1(n684), .A2(n668), .ZN(n614) );
  INV_X1 U695 ( .A(n619), .ZN(n698) );
  NOR2_X1 U696 ( .A1(n442), .A2(n698), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n671) );
  NAND2_X1 U699 ( .A1(n770), .A2(n671), .ZN(n622) );
  OR2_X1 U700 ( .A1(KEYINPUT85), .A2(KEYINPUT44), .ZN(n621) );
  INV_X1 U701 ( .A(KEYINPUT44), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n629), .A2(KEYINPUT82), .ZN(n626) );
  INV_X1 U703 ( .A(KEYINPUT76), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n760), .B(n627), .ZN(n628) );
  NOR2_X1 U705 ( .A1(n629), .A2(KEYINPUT82), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n734), .A2(G472), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(n632), .ZN(n635) );
  INV_X1 U708 ( .A(G952), .ZN(n634) );
  NOR2_X2 U709 ( .A1(n635), .A2(n744), .ZN(n637) );
  XNOR2_X1 U710 ( .A(KEYINPUT63), .B(KEYINPUT87), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n637), .B(n636), .ZN(G57) );
  XNOR2_X1 U712 ( .A(n638), .B(G134), .ZN(G36) );
  NAND2_X1 U713 ( .A1(n734), .A2(G475), .ZN(n644) );
  XOR2_X1 U714 ( .A(KEYINPUT88), .B(KEYINPUT66), .Z(n640) );
  XNOR2_X1 U715 ( .A(KEYINPUT59), .B(KEYINPUT119), .ZN(n639) );
  XOR2_X1 U716 ( .A(n640), .B(n639), .Z(n641) );
  XNOR2_X1 U717 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X2 U718 ( .A1(n645), .A2(n744), .ZN(n647) );
  XOR2_X1 U719 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(G60) );
  NAND2_X1 U721 ( .A1(n734), .A2(G210), .ZN(n651) );
  XNOR2_X1 U722 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n404), .B(n648), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X2 U725 ( .A1(n652), .A2(n744), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n653), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U727 ( .A1(n734), .A2(G217), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n656), .B(n655), .ZN(n657) );
  NOR2_X2 U729 ( .A1(n657), .A2(n744), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n658), .B(KEYINPUT122), .ZN(G66) );
  XNOR2_X1 U731 ( .A(G101), .B(KEYINPUT104), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(G3) );
  XOR2_X1 U733 ( .A(G104), .B(KEYINPUT105), .Z(n662) );
  NAND2_X1 U734 ( .A1(n668), .A2(n680), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n662), .B(n661), .ZN(G6) );
  XOR2_X1 U736 ( .A(KEYINPUT106), .B(KEYINPUT108), .Z(n664) );
  XNOR2_X1 U737 ( .A(KEYINPUT26), .B(KEYINPUT27), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U739 ( .A(n665), .B(KEYINPUT109), .Z(n667) );
  XNOR2_X1 U740 ( .A(G107), .B(KEYINPUT107), .ZN(n666) );
  XNOR2_X1 U741 ( .A(n667), .B(n666), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n668), .A2(n683), .ZN(n669) );
  XOR2_X1 U743 ( .A(n670), .B(n669), .Z(G9) );
  XNOR2_X1 U744 ( .A(G110), .B(KEYINPUT110), .ZN(n673) );
  BUF_X1 U745 ( .A(n671), .Z(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(G12) );
  XOR2_X1 U747 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n675) );
  NAND2_X1 U748 ( .A1(n678), .A2(n683), .ZN(n674) );
  XNOR2_X1 U749 ( .A(n675), .B(n674), .ZN(n676) );
  XOR2_X1 U750 ( .A(G128), .B(n676), .Z(G30) );
  XOR2_X1 U751 ( .A(G143), .B(n677), .Z(G45) );
  NAND2_X1 U752 ( .A1(n678), .A2(n680), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n679), .B(G146), .ZN(G48) );
  NAND2_X1 U754 ( .A1(n409), .A2(n680), .ZN(n681) );
  XNOR2_X1 U755 ( .A(n681), .B(KEYINPUT112), .ZN(n682) );
  XNOR2_X1 U756 ( .A(G113), .B(n682), .ZN(G15) );
  NAND2_X1 U757 ( .A1(n409), .A2(n683), .ZN(n685) );
  XNOR2_X1 U758 ( .A(n685), .B(G116), .ZN(G18) );
  XNOR2_X1 U759 ( .A(G125), .B(n686), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n687), .B(KEYINPUT37), .ZN(G27) );
  AND2_X1 U761 ( .A1(n403), .A2(n688), .ZN(n689) );
  NOR2_X1 U762 ( .A1(n689), .A2(KEYINPUT2), .ZN(n690) );
  XNOR2_X1 U763 ( .A(KEYINPUT81), .B(n690), .ZN(n692) );
  NAND2_X1 U764 ( .A1(n692), .A2(n691), .ZN(n730) );
  NOR2_X1 U765 ( .A1(n694), .A2(n425), .ZN(n695) );
  XNOR2_X1 U766 ( .A(n695), .B(KEYINPUT50), .ZN(n703) );
  NOR2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U768 ( .A(n699), .B(KEYINPUT49), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n701), .A2(n426), .ZN(n702) );
  NOR2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U771 ( .A(n704), .B(KEYINPUT113), .ZN(n706) );
  AND2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U773 ( .A(KEYINPUT51), .B(n707), .Z(n708) );
  NOR2_X1 U774 ( .A1(n725), .A2(n708), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U777 ( .A(n713), .B(KEYINPUT114), .ZN(n715) );
  NOR2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U779 ( .A1(n716), .A2(n724), .ZN(n717) );
  NOR2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n721) );
  XNOR2_X1 U781 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n719) );
  XNOR2_X1 U782 ( .A(n719), .B(KEYINPUT52), .ZN(n720) );
  XOR2_X1 U783 ( .A(n721), .B(n720), .Z(n722) );
  NOR2_X1 U784 ( .A1(n723), .A2(n722), .ZN(n727) );
  NOR2_X1 U785 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U786 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U787 ( .A(KEYINPUT117), .B(n728), .Z(n729) );
  NAND2_X1 U788 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U789 ( .A(KEYINPUT118), .B(n731), .ZN(n732) );
  NOR2_X1 U790 ( .A1(n732), .A2(G953), .ZN(n733) );
  XNOR2_X1 U791 ( .A(n733), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U792 ( .A1(n739), .A2(G469), .ZN(n737) );
  XOR2_X1 U793 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n735) );
  XNOR2_X1 U794 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U795 ( .A1(n744), .A2(n738), .ZN(G54) );
  NAND2_X1 U796 ( .A1(n739), .A2(G478), .ZN(n742) );
  NOR2_X1 U797 ( .A1(n744), .A2(n743), .ZN(G63) );
  INV_X1 U798 ( .A(n403), .ZN(n746) );
  NOR2_X1 U799 ( .A1(G953), .A2(n746), .ZN(n747) );
  XNOR2_X1 U800 ( .A(KEYINPUT123), .B(n747), .ZN(n751) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n748) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n748), .ZN(n749) );
  NAND2_X1 U803 ( .A1(n749), .A2(G898), .ZN(n750) );
  NAND2_X1 U804 ( .A1(n751), .A2(n750), .ZN(n756) );
  XNOR2_X1 U805 ( .A(KEYINPUT125), .B(n402), .ZN(n753) );
  NOR2_X1 U806 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U807 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U808 ( .A(KEYINPUT124), .B(n757), .ZN(G69) );
  XNOR2_X1 U809 ( .A(n758), .B(n759), .ZN(n763) );
  XNOR2_X1 U810 ( .A(n760), .B(n763), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n762), .A2(n761), .ZN(n768) );
  XNOR2_X1 U812 ( .A(n763), .B(G227), .ZN(n764) );
  NAND2_X1 U813 ( .A1(n764), .A2(G900), .ZN(n765) );
  XNOR2_X1 U814 ( .A(KEYINPUT126), .B(n765), .ZN(n766) );
  NAND2_X1 U815 ( .A1(n766), .A2(G953), .ZN(n767) );
  NAND2_X1 U816 ( .A1(n768), .A2(n767), .ZN(G72) );
  XNOR2_X1 U817 ( .A(n769), .B(G140), .ZN(G42) );
  XNOR2_X1 U818 ( .A(n770), .B(G119), .ZN(G21) );
  XOR2_X1 U819 ( .A(G137), .B(n771), .Z(G39) );
endmodule

