//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1191,
    new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  OR4_X1    g028(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n463), .A2(new_n465), .A3(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n473));
  INV_X1    g048(.A(G100), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(new_n461), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(new_n465), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n461), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n476), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND2_X1  g058(.A1(G102), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT4), .A2(G138), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n477), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n461), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n463), .A2(new_n465), .A3(G126), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G114), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT69), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n488), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n477), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n497), .A2(G138), .A3(new_n461), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n487), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n506), .A2(G62), .A3(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n515), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n510), .A2(KEYINPUT71), .A3(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n508), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n507), .B1(new_n520), .B2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT72), .B1(new_n518), .B2(new_n505), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n516), .A2(new_n517), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n523), .A2(new_n506), .A3(new_n524), .A4(new_n514), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n522), .A2(G88), .A3(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n521), .A2(KEYINPUT73), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT73), .B1(new_n521), .B2(new_n526), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n522), .A2(new_n525), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n518), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n523), .A2(KEYINPUT75), .A3(new_n514), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n534), .A2(G543), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT74), .Z(new_n542));
  NAND4_X1  g117(.A1(new_n532), .A2(new_n538), .A3(new_n540), .A4(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n531), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n505), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT76), .Z(new_n550));
  XOR2_X1   g125(.A(KEYINPUT77), .B(G52), .Z(new_n551));
  NAND2_X1  g126(.A1(new_n537), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n545), .A2(new_n550), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n505), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n537), .A2(G43), .B1(G651), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n531), .A2(G81), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(G860), .A3(new_n559), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  AND2_X1   g140(.A1(new_n534), .A2(new_n535), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n506), .A2(G65), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT78), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n534), .A2(G53), .A3(G543), .A4(new_n535), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n522), .A2(G91), .A3(new_n525), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n567), .A2(new_n571), .A3(new_n574), .A4(new_n575), .ZN(G299));
  NOR2_X1   g151(.A1(new_n527), .A2(new_n528), .ZN(G303));
  NAND3_X1  g152(.A1(new_n522), .A2(G87), .A3(new_n525), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n534), .A2(G49), .A3(G543), .A4(new_n535), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AND3_X1   g156(.A1(new_n506), .A2(G61), .A3(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G651), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n518), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n582), .B1(new_n585), .B2(G543), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n522), .A2(G86), .A3(new_n525), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n537), .A2(G47), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n522), .A2(G85), .A3(new_n525), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n512), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n530), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n505), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n595), .A2(new_n598), .B1(G651), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n537), .A2(G54), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n594), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n594), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G168), .B2(new_n607), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(G168), .B2(new_n607), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n557), .A2(G651), .ZN(new_n613));
  INV_X1    g188(.A(G43), .ZN(new_n614));
  INV_X1    g189(.A(G81), .ZN(new_n615));
  OAI221_X1 g190(.A(new_n613), .B1(new_n536), .B2(new_n614), .C1(new_n615), .C2(new_n530), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n604), .A2(new_n611), .ZN(new_n617));
  MUX2_X1   g192(.A(new_n616), .B(new_n617), .S(G868), .Z(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n478), .A2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n480), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT79), .B(G2100), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n625), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n637), .B(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(G14), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT18), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(KEYINPUT80), .ZN(new_n650));
  OAI21_X1  g225(.A(KEYINPUT17), .B1(new_n650), .B2(new_n645), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(new_n647), .Z(new_n652));
  AND2_X1   g227(.A1(new_n650), .A2(new_n645), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT81), .ZN(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n657), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n663), .A3(new_n661), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n661), .A2(new_n657), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n665), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n664), .B(new_n667), .C1(new_n669), .C2(new_n663), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1991), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1986), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(G229));
  NAND2_X1  g251(.A1(new_n480), .A2(G139), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT25), .Z(new_n679));
  AOI22_X1  g254(.A1(new_n497), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n679), .C1(new_n680), .C2(new_n461), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT88), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT89), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G29), .ZN(new_n684));
  INV_X1    g259(.A(G33), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(G29), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G2072), .ZN(new_n687));
  INV_X1    g262(.A(G2072), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n684), .B(new_n688), .C1(G29), .C2(new_n685), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G35), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G162), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  INV_X1    g269(.A(G2090), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n687), .A2(new_n689), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n478), .A2(G129), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n480), .A2(G141), .ZN(new_n699));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT26), .Z(new_n701));
  NAND3_X1  g276(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT90), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G32), .B(new_n704), .S(G29), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT27), .B(G1996), .Z(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT91), .ZN(new_n708));
  NAND2_X1  g283(.A1(G171), .A2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G5), .B2(G16), .ZN(new_n710));
  INV_X1    g285(.A(G1961), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n695), .A2(new_n694), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n690), .A2(G26), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n478), .A2(G128), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n480), .A2(G140), .ZN(new_n715));
  NOR2_X1   g290(.A1(G104), .A2(G2105), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n714), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n713), .B1(new_n718), .B2(G29), .ZN(new_n719));
  MUX2_X1   g294(.A(new_n713), .B(new_n719), .S(KEYINPUT28), .Z(new_n720));
  INV_X1    g295(.A(G2067), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  NOR2_X1   g298(.A1(G164), .A2(new_n690), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G27), .B2(new_n690), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n722), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  NAND2_X1  g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n727), .A2(new_n690), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G160), .B2(new_n690), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n705), .A2(new_n706), .B1(G2084), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n624), .A2(new_n690), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n690), .B1(new_n733), .B2(G28), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(KEYINPUT93), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n734), .A2(KEYINPUT93), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n735), .B(new_n736), .C1(new_n733), .C2(G28), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n731), .B(new_n738), .C1(G2084), .C2(new_n730), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n725), .A2(new_n723), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  NOR3_X1   g316(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n712), .A2(new_n726), .A3(new_n742), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n697), .A2(new_n708), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n710), .A2(new_n711), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT94), .ZN(new_n746));
  INV_X1    g321(.A(G16), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n604), .B2(new_n747), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1348), .ZN(new_n750));
  MUX2_X1   g325(.A(G19), .B(new_n616), .S(G16), .Z(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT87), .B(G1341), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n747), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n747), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT92), .B(G1966), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n750), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n747), .A2(G20), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT96), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  INV_X1    g336(.A(G299), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n747), .ZN(new_n763));
  INV_X1    g338(.A(G1956), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n744), .A2(new_n746), .A3(new_n758), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT97), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT98), .ZN(new_n768));
  NOR2_X1   g343(.A1(G16), .A2(G22), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G166), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1971), .ZN(new_n771));
  MUX2_X1   g346(.A(G6), .B(G305), .S(G16), .Z(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT32), .B(G1981), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(KEYINPUT84), .B1(G16), .B2(G23), .ZN(new_n776));
  OR3_X1    g351(.A1(KEYINPUT84), .A2(G16), .A3(G23), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT85), .ZN(new_n778));
  NAND2_X1  g353(.A1(G288), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT85), .A4(new_n580), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n776), .B(new_n777), .C1(new_n782), .C2(new_n747), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT33), .B(G1976), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n775), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n478), .A2(G119), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT82), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(G95), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n480), .A2(G131), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT83), .ZN(new_n795));
  MUX2_X1   g370(.A(G25), .B(new_n795), .S(G29), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT35), .B(G1991), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n747), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n747), .B2(G24), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n798), .B1(G1986), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n787), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT86), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT34), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n775), .A2(new_n810), .A3(new_n785), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n804), .A2(new_n807), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n787), .A2(new_n803), .A3(new_n809), .A4(new_n811), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n813), .A2(new_n805), .A3(new_n806), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n805), .A2(new_n806), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n767), .B(new_n768), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n766), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n816), .B1(new_n812), .B2(new_n814), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT98), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n817), .A2(new_n821), .ZN(G311));
  OAI21_X1  g397(.A(new_n767), .B1(new_n815), .B2(new_n816), .ZN(G150));
  NAND3_X1  g398(.A1(new_n522), .A2(G93), .A3(new_n525), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n505), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT99), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n824), .B1(new_n536), .B2(new_n825), .C1(new_n829), .C2(new_n512), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n602), .A2(new_n603), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n611), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n830), .A2(new_n559), .A3(new_n558), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n829), .A2(new_n512), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n536), .A2(new_n825), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n616), .A2(new_n839), .A3(new_n824), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT39), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n835), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n832), .B1(new_n843), .B2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT100), .Z(G145));
  INV_X1    g420(.A(G160), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n624), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n478), .A2(G130), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n480), .A2(G142), .ZN(new_n850));
  NOR2_X1   g425(.A1(G106), .A2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n627), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n795), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n482), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n482), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n848), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n847), .A3(new_n856), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n718), .B(KEYINPUT101), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G164), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(new_n704), .Z(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n683), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n682), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n859), .A2(new_n861), .A3(new_n867), .A4(new_n868), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g449(.A(new_n799), .B1(new_n527), .B2(new_n528), .ZN(new_n875));
  NAND2_X1  g450(.A1(G303), .A2(G290), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n781), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(G305), .B(KEYINPUT102), .Z(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n781), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n799), .A2(new_n527), .A3(new_n528), .ZN(new_n883));
  NOR2_X1   g458(.A1(G303), .A2(G290), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n782), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n879), .B1(new_n885), .B2(new_n877), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n833), .A2(G299), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n833), .A2(G299), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n617), .B(new_n841), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n891), .A2(new_n892), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n897), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n888), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n888), .A2(new_n900), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n607), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n830), .A2(new_n607), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n903), .A2(KEYINPUT103), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT103), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(G295));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n901), .A2(new_n902), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G868), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n911), .B2(new_n904), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n903), .A2(KEYINPUT104), .A3(new_n905), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(G331));
  NAND3_X1  g489(.A1(new_n836), .A2(new_n840), .A3(G286), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(G286), .B1(new_n836), .B2(new_n840), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n916), .A2(new_n917), .A3(G301), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n841), .A2(G168), .ZN(new_n919));
  AOI21_X1  g494(.A(G171), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n893), .B(new_n895), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(G301), .B1(new_n916), .B2(new_n917), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(G171), .A3(new_n915), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n899), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n887), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n887), .B1(new_n921), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .A4(new_n871), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n921), .A2(new_n924), .ZN(new_n931));
  INV_X1    g506(.A(new_n887), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n887), .A2(new_n921), .A3(new_n924), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n871), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n933), .A2(new_n929), .A3(new_n871), .A4(new_n934), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT105), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n930), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(KEYINPUT44), .A3(new_n937), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(G397));
  INV_X1    g518(.A(KEYINPUT55), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(G303), .B2(G8), .ZN(new_n945));
  INV_X1    g520(.A(G8), .ZN(new_n946));
  NOR4_X1   g521(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT55), .A4(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n499), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT112), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n497), .A2(G138), .A3(new_n461), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n461), .B1(new_n489), .B2(new_n494), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(new_n488), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n955), .B2(new_n487), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n952), .A2(KEYINPUT50), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT106), .B1(G160), .B2(G40), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  INV_X1    g536(.A(G40), .ZN(new_n962));
  NOR4_X1   g537(.A1(new_n468), .A2(new_n471), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n956), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n959), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  AOI21_X1  g543(.A(G2090), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n964), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n957), .B1(new_n499), .B2(new_n950), .ZN(new_n971));
  AOI211_X1 g546(.A(KEYINPUT112), .B(G1384), .C1(new_n955), .C2(new_n487), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n970), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT115), .A3(new_n966), .ZN(new_n975));
  INV_X1    g550(.A(G1971), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n951), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n956), .A2(KEYINPUT45), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n956), .B2(KEYINPUT45), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n977), .B(G1384), .C1(new_n955), .C2(new_n487), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n964), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n969), .A2(new_n975), .B1(new_n976), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n949), .B1(new_n987), .B2(new_n946), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n964), .B1(new_n971), .B2(new_n972), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G8), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n779), .B2(new_n780), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n993));
  INV_X1    g568(.A(G288), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(G1976), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n990), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n997));
  INV_X1    g572(.A(G1981), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n586), .A2(new_n998), .A3(new_n587), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n586), .B2(new_n587), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G305), .A2(G1981), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n586), .A2(new_n998), .A3(new_n587), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(KEYINPUT49), .A3(new_n1003), .ZN(new_n1004));
  AND4_X1   g579(.A1(G8), .A2(new_n1001), .A3(new_n1004), .A4(new_n989), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT52), .B1(new_n990), .B2(new_n992), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n990), .C2(new_n992), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n996), .B(new_n1005), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n970), .B1(new_n981), .B2(new_n984), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n951), .A2(KEYINPUT50), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n964), .A3(new_n1013), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n1011), .A2(G1971), .B1(new_n1014), .B2(G2090), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(G8), .A3(new_n948), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n970), .B1(new_n973), .B2(new_n977), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1966), .B1(new_n1017), .B2(new_n980), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1014), .A2(G2084), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1020), .A2(new_n946), .A3(G286), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n988), .A2(new_n1010), .A3(new_n1016), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT63), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n996), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1005), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n781), .A2(G1976), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(G8), .A3(new_n989), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT113), .B1(new_n1028), .B2(KEYINPUT52), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1009), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1025), .B(new_n1026), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n948), .B1(new_n1015), .B2(G8), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT116), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1016), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n952), .A2(new_n977), .A3(new_n958), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(new_n964), .A3(new_n980), .ZN(new_n1036));
  INV_X1    g611(.A(G1966), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(G2084), .B2(new_n1014), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1015), .A2(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n949), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1025), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1033), .A2(new_n1041), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1024), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n990), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1005), .A2(G1976), .A3(G288), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1050), .B2(new_n999), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n1031), .B2(new_n1016), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT114), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1051), .B(new_n1054), .C1(new_n1031), .C2(new_n1016), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n967), .A2(new_n764), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n531), .A2(G91), .B1(new_n573), .B2(new_n572), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n571), .A4(new_n567), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n982), .A2(new_n983), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n951), .A2(new_n979), .A3(new_n977), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n964), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1057), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1348), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1014), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n989), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT117), .B(new_n964), .C1(new_n971), .C2(new_n972), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n721), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1067), .A2(new_n604), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1062), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1956), .B1(new_n974), .B2(new_n966), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1063), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n970), .B(new_n1078), .C1(new_n981), .C2(new_n984), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(G1341), .ZN(new_n1084));
  INV_X1    g659(.A(G1996), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1082), .A2(new_n1084), .B1(new_n1011), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n1087));
  OR3_X1    g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n616), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1057), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1062), .B1(new_n1057), .B2(new_n1066), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1080), .A2(new_n1067), .A3(KEYINPUT61), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1087), .B1(new_n1086), .B2(new_n616), .ZN(new_n1094));
  AND4_X1   g669(.A1(new_n1088), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n1074), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1069), .A2(new_n1073), .A3(KEYINPUT119), .A4(KEYINPUT60), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n604), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1074), .A2(new_n1097), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1096), .B(new_n833), .C1(new_n1074), .C2(new_n1097), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1081), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n969), .A2(new_n975), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n986), .A2(new_n976), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n948), .B1(new_n1107), .B2(G8), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1044), .A2(new_n1016), .A3(new_n1025), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G286), .A2(G8), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT120), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1039), .B2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1039), .B(G8), .C1(KEYINPUT121), .C2(new_n1113), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1113), .A2(KEYINPUT121), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1020), .B2(new_n946), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1114), .B(new_n1115), .C1(new_n1117), .C2(new_n1112), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT123), .B1(new_n1036), .B2(G2078), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1017), .A2(new_n1120), .A3(new_n723), .A4(new_n980), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(KEYINPUT53), .A3(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n723), .B(new_n964), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1123), .A2(new_n1124), .B1(new_n1014), .B2(new_n711), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(G301), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1014), .A2(new_n711), .ZN(new_n1128));
  NAND2_X1  g703(.A1(G160), .A2(G40), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n985), .A2(KEYINPUT53), .A3(new_n723), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(G171), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1126), .A2(new_n1133), .A3(KEYINPUT54), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1135));
  AOI21_X1  g710(.A(G301), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1132), .A2(G171), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1110), .A2(new_n1118), .A3(new_n1134), .A4(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1048), .B(new_n1056), .C1(new_n1104), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1118), .A2(KEYINPUT62), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1118), .A2(KEYINPUT62), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n1110), .A4(new_n1136), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1024), .A2(new_n1047), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1146), .B(KEYINPUT125), .C1(new_n1104), .C2(new_n1139), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n970), .A2(new_n978), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(G1996), .A3(new_n704), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1150), .A2(KEYINPUT109), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n718), .B(new_n721), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(G1996), .B2(new_n704), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1149), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(KEYINPUT109), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1156), .B(KEYINPUT110), .Z(new_n1157));
  AND2_X1   g732(.A1(new_n795), .A2(new_n797), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n795), .A2(new_n797), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1149), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n799), .A2(new_n808), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT107), .ZN(new_n1163));
  NAND2_X1  g738(.A1(G290), .A2(G1986), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT108), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1161), .B1(new_n1149), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1148), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1163), .A2(new_n1149), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT126), .Z(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT48), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1171), .A2(new_n1161), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT46), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1149), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1174), .B2(G1996), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1152), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1149), .B1(new_n704), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1149), .A2(KEYINPUT46), .A3(new_n1085), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT47), .Z(new_n1180));
  NAND2_X1  g755(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n718), .A2(G2067), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1174), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1172), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1168), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g760(.A1(G401), .A2(G227), .ZN(new_n1187));
  AND2_X1   g761(.A1(new_n873), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g762(.A1(G229), .A2(new_n459), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n939), .A2(new_n1188), .A3(new_n1189), .ZN(G225));
  NAND2_X1  g764(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1191));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n1192));
  NAND4_X1  g766(.A1(new_n939), .A2(new_n1188), .A3(new_n1192), .A4(new_n1189), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1193), .ZN(G308));
endmodule


