//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n538, new_n540, new_n541, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT68), .Z(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  NAND3_X1  g032(.A1(new_n457), .A2(G101), .A3(G2104), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(new_n459));
  INV_X1    g034(.A(G137), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(new_n457), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(new_n457), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(G160));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n471), .A2(new_n457), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n457), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  NAND4_X1  g054(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n457), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n461), .A2(KEYINPUT4), .A3(G138), .A4(new_n457), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT70), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n485), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n484), .B1(new_n491), .B2(new_n493), .ZN(G164));
  AND2_X1   g069(.A1(KEYINPUT6), .A2(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT6), .A2(G651), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G50), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n496), .B2(new_n495), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n498), .A2(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  XOR2_X1   g084(.A(new_n509), .B(KEYINPUT71), .Z(new_n510));
  NAND2_X1  g085(.A1(new_n504), .A2(G62), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(new_n512), .ZN(G166));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  INV_X1    g090(.A(G51), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n498), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n504), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n497), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(G168));
  AOI22_X1  g097(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n508), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT72), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n495), .A2(new_n496), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n501), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(G90), .B1(G52), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  AOI22_X1  g106(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n508), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT73), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n527), .A2(G81), .B1(G43), .B2(new_n528), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G860), .ZN(G153));
  AND3_X1   g112(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G36), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(G188));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n505), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n497), .A2(KEYINPUT75), .A3(new_n504), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G91), .ZN(new_n547));
  NAND2_X1  g122(.A1(KEYINPUT74), .A2(G53), .ZN(new_n548));
  OR3_X1    g123(.A1(new_n498), .A2(KEYINPUT9), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT9), .B1(new_n498), .B2(new_n548), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n508), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n547), .A2(new_n551), .A3(new_n553), .ZN(G299));
  INV_X1    g129(.A(G168), .ZN(G286));
  INV_X1    g130(.A(G166), .ZN(G303));
  NAND3_X1  g131(.A1(new_n544), .A2(new_n545), .A3(G87), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT76), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n544), .A2(new_n545), .A3(new_n559), .A4(G87), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n504), .A2(G74), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(new_n528), .B2(G49), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G288));
  OAI211_X1 g139(.A(G48), .B(G543), .C1(new_n495), .C2(new_n496), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n544), .A2(new_n545), .A3(G86), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n504), .A2(G61), .ZN(new_n571));
  AND2_X1   g146(.A1(G73), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n569), .A2(new_n570), .A3(new_n573), .ZN(G305));
  INV_X1    g149(.A(G47), .ZN(new_n575));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n498), .A2(new_n575), .B1(new_n505), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n508), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n577), .A2(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n546), .A2(G92), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT10), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n518), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n528), .B2(G54), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n581), .A2(KEYINPUT78), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n582), .B1(new_n592), .B2(new_n593), .ZN(G284));
  AOI21_X1  g169(.A(new_n582), .B1(new_n592), .B2(new_n593), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  AND2_X1   g174(.A1(new_n585), .A2(new_n589), .ZN(new_n600));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G860), .ZN(G148));
  NOR2_X1   g177(.A1(new_n590), .A2(G559), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n536), .ZN(G323));
  XOR2_X1   g181(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n607));
  XNOR2_X1  g182(.A(G323), .B(new_n607), .ZN(G282));
  NAND2_X1  g183(.A1(new_n472), .A2(G2104), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n472), .A2(G135), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n474), .A2(G123), .ZN(new_n616));
  NOR3_X1   g191(.A1(new_n457), .A2(KEYINPUT80), .A3(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT80), .B1(new_n457), .B2(G111), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n618), .A2(G2104), .A3(new_n619), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n613), .A2(new_n614), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n633), .A2(new_n636), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(G401));
  XNOR2_X1  g215(.A(G2084), .B(G2090), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT82), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT17), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n642), .A2(new_n644), .ZN(new_n650));
  NOR2_X1   g225(.A1(G2072), .A2(G2078), .ZN(new_n651));
  OAI22_X1  g226(.A1(new_n650), .A2(new_n648), .B1(new_n442), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2096), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n661), .A2(KEYINPUT84), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT83), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n661), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT20), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n680), .A3(new_n678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G16), .A2(G23), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(G288), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT90), .Z(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT33), .B(G1976), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  MUX2_X1   g267(.A(G6), .B(G305), .S(G16), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT32), .B(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n687), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n687), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1971), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n691), .A2(new_n692), .A3(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  AOI22_X1  g279(.A1(G119), .A2(new_n474), .B1(new_n472), .B2(G131), .ZN(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n706));
  INV_X1    g281(.A(G107), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G2105), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT86), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n710), .B2(new_n703), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  MUX2_X1   g288(.A(G24), .B(G290), .S(G16), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT87), .B(G1986), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT88), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n713), .B(new_n717), .C1(KEYINPUT91), .C2(KEYINPUT36), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n701), .A2(new_n702), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n703), .A2(G35), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G162), .B2(new_n703), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT29), .Z(new_n724));
  INV_X1    g299(.A(G2090), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT97), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n687), .A2(G19), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n536), .B2(new_n687), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1341), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G5), .A2(G16), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT96), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G301), .B2(new_n687), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n703), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n703), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2078), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n703), .A2(G32), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT26), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G129), .B2(new_n474), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n467), .A2(G2105), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n472), .A2(G141), .B1(G105), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT95), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n724), .B2(new_n725), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n457), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n472), .A2(G139), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n754), .B(new_n755), .C1(new_n457), .C2(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G33), .B(new_n757), .S(G29), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G2072), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT24), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n703), .B1(new_n760), .B2(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n760), .B2(G34), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G160), .B2(G29), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n687), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n687), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n759), .B1(G2084), .B2(new_n763), .C1(G1966), .C2(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT31), .B(G11), .Z(new_n767));
  NOR2_X1   g342(.A1(new_n621), .A2(new_n703), .ZN(new_n768));
  INV_X1    g343(.A(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT30), .ZN(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n769), .B2(KEYINPUT30), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n767), .B(new_n768), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n765), .A2(G1966), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n748), .A2(new_n749), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n763), .A2(G2084), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n772), .A2(new_n773), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n752), .A2(new_n766), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n687), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n597), .B2(new_n687), .ZN(new_n780));
  INV_X1    g355(.A(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT94), .B1(new_n758), .B2(G2072), .ZN(new_n783));
  OR3_X1    g358(.A1(new_n758), .A2(KEYINPUT94), .A3(G2072), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n703), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n472), .A2(G140), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n474), .A2(G128), .ZN(new_n788));
  OR2_X1    g363(.A1(G104), .A2(G2105), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n789), .B(G2104), .C1(G116), .C2(new_n457), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n786), .B1(new_n792), .B2(new_n703), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT93), .B(G2067), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AND4_X1   g370(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n731), .A2(new_n740), .A3(new_n777), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G4), .A2(G16), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n600), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT92), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1348), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n719), .B2(new_n720), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n721), .A2(new_n803), .ZN(G311));
  OR2_X1    g379(.A1(new_n721), .A2(new_n803), .ZN(G150));
  AOI22_X1  g380(.A1(new_n527), .A2(G93), .B1(G55), .B2(new_n528), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(new_n508), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n536), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n812), .B2(new_n811), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n536), .A2(KEYINPUT99), .A3(new_n810), .A4(new_n808), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT38), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n590), .A2(new_n601), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT100), .B(G860), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n808), .B2(new_n810), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT37), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(G145));
  XNOR2_X1  g401(.A(new_n710), .B(new_n610), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n474), .A2(G130), .ZN(new_n828));
  OR2_X1    g403(.A1(G106), .A2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(G2104), .C1(G118), .C2(new_n457), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G142), .B2(new_n472), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n827), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT102), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n485), .A2(KEYINPUT101), .A3(new_n489), .ZN(new_n835));
  AOI21_X1  g410(.A(KEYINPUT101), .B1(new_n485), .B2(new_n489), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n482), .B(new_n483), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n791), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n757), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(new_n747), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n834), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n621), .B(new_n478), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(G160), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G37), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n843), .B1(new_n834), .B2(new_n840), .ZN(new_n846));
  INV_X1    g421(.A(new_n833), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g425(.A1(new_n816), .A2(new_n604), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n814), .A2(new_n603), .A3(new_n815), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n585), .A2(new_n597), .A3(new_n589), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n597), .B1(new_n585), .B2(new_n589), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n859));
  INV_X1    g434(.A(new_n856), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n860), .B2(new_n854), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n855), .A2(KEYINPUT41), .A3(new_n856), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n858), .B1(new_n863), .B2(new_n853), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT42), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(KEYINPUT104), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI221_X1 g442(.A(new_n858), .B1(KEYINPUT104), .B2(new_n865), .C1(new_n863), .C2(new_n853), .ZN(new_n868));
  XNOR2_X1  g443(.A(G305), .B(G166), .ZN(new_n869));
  INV_X1    g444(.A(new_n563), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n558), .B2(new_n560), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G290), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(KEYINPUT104), .B2(new_n865), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n867), .A2(new_n868), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n867), .B2(new_n868), .ZN(new_n880));
  OAI21_X1  g455(.A(G868), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n811), .A2(new_n591), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(G295));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n882), .ZN(G331));
  XNOR2_X1  g459(.A(G301), .B(G168), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n816), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n814), .A2(new_n815), .A3(new_n885), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(new_n857), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n860), .A2(new_n859), .A3(new_n854), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT41), .B1(new_n855), .B2(new_n856), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n887), .A2(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n877), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n857), .A3(new_n888), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n814), .A2(new_n815), .A3(new_n885), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n885), .B1(new_n814), .B2(new_n815), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n894), .B(new_n876), .C1(new_n897), .C2(new_n863), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n845), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n891), .A2(new_n890), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n862), .A2(KEYINPUT106), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n905), .B(new_n906), .C1(new_n895), .C2(new_n896), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n894), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n877), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(new_n845), .A3(new_n898), .A4(new_n900), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n902), .A2(new_n903), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n898), .A2(new_n845), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n876), .B1(new_n907), .B2(new_n894), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n893), .A2(new_n898), .A3(new_n845), .A4(new_n900), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n903), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n911), .A2(new_n916), .ZN(G397));
  INV_X1    g492(.A(G1384), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n837), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(G160), .A2(G40), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G1996), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n747), .B(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G2067), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n791), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n710), .B(new_n712), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n923), .ZN(new_n931));
  XOR2_X1   g506(.A(G290), .B(G1986), .Z(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT107), .ZN(new_n934));
  NAND2_X1  g509(.A1(G303), .A2(G8), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT55), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(KEYINPUT110), .B(G1971), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G40), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n463), .A2(new_n465), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n485), .A2(new_n492), .A3(new_n489), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n492), .B1(new_n485), .B2(new_n489), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n482), .B(new_n483), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n918), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n942), .B1(new_n946), .B2(new_n920), .ZN(new_n947));
  AOI211_X1 g522(.A(KEYINPUT108), .B(KEYINPUT45), .C1(new_n945), .C2(new_n918), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n835), .A2(new_n836), .ZN(new_n950));
  OAI211_X1 g525(.A(KEYINPUT45), .B(new_n918), .C1(new_n950), .C2(new_n484), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT109), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n837), .A2(new_n953), .A3(KEYINPUT45), .A4(new_n918), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(KEYINPUT111), .B(new_n939), .C1(new_n949), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n837), .A2(new_n958), .A3(new_n918), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT112), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n837), .A2(new_n961), .A3(new_n958), .A4(new_n918), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n960), .A2(new_n941), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n957), .B1(new_n964), .B2(G2090), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n960), .A2(new_n941), .A3(new_n963), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n966), .A2(KEYINPUT113), .A3(new_n725), .A4(new_n962), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n956), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n491), .A2(new_n493), .ZN(new_n969));
  INV_X1    g544(.A(new_n484), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT108), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n946), .A2(new_n942), .A3(new_n920), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n922), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n952), .A2(new_n954), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n938), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(KEYINPUT111), .ZN(new_n977));
  OAI211_X1 g552(.A(G8), .B(new_n937), .C1(new_n968), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n871), .A2(G1976), .ZN(new_n979));
  INV_X1    g554(.A(new_n836), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n485), .A2(KEYINPUT101), .A3(new_n489), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n982), .B2(new_n970), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n941), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(G8), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT52), .ZN(new_n986));
  INV_X1    g561(.A(G1976), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT52), .B1(G288), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n922), .A2(new_n919), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n991), .A3(new_n979), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n527), .A2(G86), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n573), .A2(new_n993), .A3(new_n568), .A4(new_n567), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G1981), .ZN(new_n995));
  INV_X1    g570(.A(G1981), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n569), .A2(new_n570), .A3(new_n996), .A4(new_n573), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(KEYINPUT114), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(KEYINPUT114), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n997), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n991), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n986), .A2(new_n992), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n941), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n983), .A2(new_n958), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1005), .A2(new_n1006), .A3(G2090), .ZN(new_n1007));
  OAI21_X1  g582(.A(G8), .B1(new_n976), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n1008), .B2(new_n936), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n978), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n945), .A2(KEYINPUT45), .A3(new_n918), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT116), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n971), .A2(new_n1014), .A3(KEYINPUT45), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1013), .A2(new_n1015), .A3(new_n941), .A4(new_n921), .ZN(new_n1016));
  INV_X1    g591(.A(G1966), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n922), .B1(KEYINPUT50), .B2(new_n946), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT117), .B(G2084), .Z(new_n1020));
  NAND4_X1  g595(.A1(new_n1019), .A2(new_n962), .A3(new_n960), .A4(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(G168), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  AOI21_X1  g598(.A(G168), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT51), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT62), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n972), .A2(new_n973), .ZN(new_n1031));
  INV_X1    g606(.A(G2078), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1031), .A2(new_n975), .A3(new_n1032), .A4(new_n941), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1034), .A2(G2078), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n921), .A2(new_n941), .A3(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1036), .A2(new_n1038), .B1(new_n964), .B2(new_n735), .ZN(new_n1039));
  AOI21_X1  g614(.A(G301), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1011), .A2(new_n1029), .A3(new_n1030), .A4(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n978), .A2(new_n1009), .A3(new_n1040), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT124), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1022), .A2(new_n1027), .A3(G8), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1021), .ZN(new_n1047));
  OAI21_X1  g622(.A(G286), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(G8), .A3(new_n1022), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1045), .B1(new_n1049), .B2(KEYINPUT51), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT125), .B1(new_n1050), .B2(new_n1026), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1050), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT125), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(KEYINPUT62), .ZN(new_n1054));
  AND4_X1   g629(.A1(new_n1041), .A2(new_n1044), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1003), .A2(new_n987), .A3(new_n871), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n997), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n991), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1004), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n986), .A2(new_n992), .A3(new_n1003), .A4(KEYINPUT115), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1058), .B1(new_n1062), .B2(new_n978), .ZN(new_n1063));
  AOI211_X1 g638(.A(new_n990), .B(G286), .C1(new_n1018), .C2(new_n1021), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n978), .A2(new_n1009), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT63), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(G8), .B1(new_n968), .B2(new_n977), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n936), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G286), .A2(new_n990), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT63), .B(new_n1070), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1069), .A2(new_n978), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1063), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1010), .A2(new_n1050), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n1076));
  XNOR2_X1  g651(.A(G299), .B(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1031), .A2(new_n975), .A3(new_n941), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n781), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n984), .A2(G2067), .ZN(new_n1082));
  INV_X1    g657(.A(G1348), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n964), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n590), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1079), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1081), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1031), .A2(new_n975), .A3(new_n924), .A4(new_n941), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT58), .B(G1341), .Z(new_n1089));
  NAND2_X1  g664(.A1(new_n984), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n536), .A2(KEYINPUT118), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n964), .A2(new_n1083), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n590), .B1(new_n1097), .B2(new_n1082), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1084), .B2(new_n600), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1084), .A2(new_n1099), .A3(new_n600), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1096), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1079), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n1081), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1077), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(KEYINPUT61), .A3(new_n1086), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1087), .B1(new_n1104), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1038), .A2(new_n975), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1035), .A2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n964), .A2(KEYINPUT120), .A3(new_n735), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT120), .B1(new_n964), .B2(new_n735), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT123), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n964), .A2(new_n735), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n964), .A2(KEYINPUT120), .A3(new_n735), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1035), .A4(new_n1114), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1119), .A2(G171), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1035), .A2(new_n1039), .A3(G301), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1035), .A2(new_n1039), .A3(KEYINPUT122), .A4(G301), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1127), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1075), .A2(new_n1113), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1124), .A2(G301), .A3(new_n1035), .A4(new_n1114), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1040), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1136), .B1(new_n1139), .B2(new_n1128), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT121), .B(KEYINPUT54), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1074), .B1(new_n1135), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n934), .B1(new_n1055), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT48), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G290), .A2(G1986), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1145), .B1(new_n931), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n923), .A2(KEYINPUT48), .A3(new_n1146), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1148), .A2(new_n930), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT46), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n931), .B2(G1996), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n923), .A2(KEYINPUT46), .A3(new_n924), .ZN(new_n1153));
  INV_X1    g728(.A(new_n927), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n923), .B1(new_n1154), .B2(new_n747), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1156), .B(KEYINPUT47), .Z(new_n1157));
  NAND2_X1  g732(.A1(new_n710), .A2(new_n712), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n928), .A2(new_n1158), .B1(G2067), .B2(new_n791), .ZN(new_n1159));
  AOI211_X1 g734(.A(new_n1150), .B(new_n1157), .C1(new_n923), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1144), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g736(.A(G229), .ZN(new_n1163));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1164));
  OAI21_X1  g738(.A(G319), .B1(new_n638), .B2(new_n639), .ZN(new_n1165));
  OR3_X1    g739(.A1(G227), .A2(new_n1165), .A3(KEYINPUT126), .ZN(new_n1166));
  OAI21_X1  g740(.A(KEYINPUT126), .B1(G227), .B2(new_n1165), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AND3_X1   g742(.A1(new_n1163), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1170));
  OAI21_X1  g744(.A(new_n849), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1171), .B1(new_n902), .B2(new_n910), .ZN(G308));
  NAND2_X1  g746(.A1(new_n902), .A2(new_n910), .ZN(new_n1173));
  OAI211_X1 g747(.A(new_n1173), .B(new_n849), .C1(new_n1170), .C2(new_n1169), .ZN(G225));
endmodule


