//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT64), .Z(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  AND2_X1   g0046(.A1(G1), .A2(G13), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n249), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G222), .A2(G1698), .ZN(new_n257));
  XOR2_X1   g0057(.A(KEYINPUT67), .B(G223), .Z(new_n258));
  AOI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G1698), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n259), .B2(new_n254), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT66), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n263), .B(new_n205), .C1(G41), .C2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n266), .B1(new_n247), .B2(new_n248), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G226), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n205), .A2(new_n272), .B1(new_n247), .B2(new_n248), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n260), .B(new_n268), .C1(new_n269), .C2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n214), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n206), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n280), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G50), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n206), .B1(new_n201), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n279), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n286), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n205), .A2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G50), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT69), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n279), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n289), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT68), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n290), .A2(new_n279), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n297), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n293), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n277), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT70), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(KEYINPUT70), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n307), .B(new_n308), .C1(G179), .C2(new_n275), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT74), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n293), .A2(KEYINPUT73), .A3(new_n304), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT73), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n299), .A2(new_n300), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n296), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n312), .B1(new_n315), .B2(new_n292), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT9), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n311), .A2(new_n316), .A3(KEYINPUT74), .A4(KEYINPUT9), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n275), .A2(G200), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n275), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n318), .B2(new_n317), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n322), .B1(new_n321), .B2(new_n326), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n309), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n251), .A2(new_n253), .A3(G232), .A4(G1698), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT3), .B(G33), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT75), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(G232), .A4(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G1698), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n251), .A2(new_n253), .A3(G226), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n249), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n265), .A2(new_n267), .B1(new_n273), .B2(G238), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT13), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n339), .B1(new_n334), .B2(new_n331), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n345), .B(new_n342), .C1(new_n346), .C2(new_n249), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT78), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(G169), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n276), .B1(new_n344), .B2(new_n347), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT78), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n349), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n344), .A2(G179), .A3(new_n347), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n351), .A2(new_n353), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n283), .A2(G50), .ZN(new_n359));
  XOR2_X1   g0159(.A(new_n359), .B(KEYINPUT76), .Z(new_n360));
  OAI22_X1  g0160(.A1(new_n281), .A2(new_n255), .B1(new_n206), .B2(G68), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n279), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT11), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT11), .B(new_n279), .C1(new_n360), .C2(new_n361), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n364), .A2(KEYINPUT77), .A3(new_n365), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT12), .B1(new_n289), .B2(G68), .ZN(new_n370));
  OR3_X1    g0170(.A1(new_n289), .A2(KEYINPUT12), .A3(G68), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n218), .B1(new_n205), .B2(G20), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n370), .A2(new_n371), .B1(new_n302), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n358), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n348), .A2(new_n324), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n344), .B2(new_n347), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n374), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G244), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n268), .B1(new_n382), .B2(new_n274), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n332), .A2(G232), .A3(new_n336), .ZN(new_n384));
  INV_X1    g0184(.A(G107), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n332), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n254), .A2(new_n219), .A3(new_n336), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n249), .B1(new_n388), .B2(KEYINPUT71), .ZN(new_n389));
  OR3_X1    g0189(.A1(new_n386), .A2(KEYINPUT71), .A3(new_n387), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n383), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G179), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n280), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT15), .B(G87), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  OR3_X1    g0198(.A1(new_n397), .A2(new_n398), .A3(new_n281), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n397), .B2(new_n281), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n279), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n294), .A2(G77), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n302), .A2(new_n404), .B1(new_n255), .B2(new_n290), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n391), .B2(G169), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n394), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n391), .B2(G190), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n377), .B2(new_n391), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n269), .A2(G1698), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G223), .B2(G1698), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n414), .A2(new_n254), .B1(new_n250), .B2(new_n220), .ZN(new_n415));
  INV_X1    g0215(.A(new_n249), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n265), .A2(new_n267), .B1(new_n273), .B2(G232), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n417), .A2(new_n418), .A3(G190), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n377), .B1(new_n417), .B2(new_n418), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G58), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n218), .ZN(new_n423));
  OAI21_X1  g0223(.A(G20), .B1(new_n423), .B2(new_n201), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n283), .A2(G159), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n251), .B2(new_n253), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n252), .A2(G33), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n206), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT7), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(KEYINPUT16), .B(new_n426), .C1(new_n433), .C2(new_n218), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n424), .A2(new_n425), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT79), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n252), .B2(G33), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n250), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n253), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n427), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n432), .B1(new_n332), .B2(G20), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n435), .B1(new_n443), .B2(G68), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n279), .B(new_n434), .C1(new_n444), .C2(KEYINPUT16), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n280), .B1(new_n205), .B2(G20), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n301), .B2(new_n303), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n280), .A2(new_n290), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n421), .A2(new_n445), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n447), .A2(new_n448), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n254), .A2(new_n440), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n442), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n435), .B1(new_n456), .B2(G68), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n298), .B1(new_n457), .B2(KEYINPUT16), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT16), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n218), .B1(new_n441), .B2(new_n442), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(new_n435), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n454), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n452), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n462), .A2(new_n450), .A3(new_n421), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n453), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(KEYINPUT80), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n445), .A2(new_n449), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n417), .A2(new_n418), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n392), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(G169), .B2(new_n471), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n467), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT18), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT18), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n467), .A2(new_n470), .A3(new_n474), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n466), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NOR4_X1   g0279(.A1(new_n329), .A2(new_n381), .A3(new_n412), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n271), .A2(G1), .ZN(new_n481));
  AND2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n484), .A2(G264), .A3(new_n249), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n251), .A2(new_n253), .A3(G257), .A4(G1698), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n251), .A2(new_n253), .A3(G250), .A4(new_n336), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G294), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n249), .B1(new_n489), .B2(KEYINPUT92), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT92), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n486), .A2(new_n487), .A3(new_n491), .A4(new_n488), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n485), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n267), .A2(new_n481), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n276), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n495), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n497), .B(new_n485), .C1(new_n490), .C2(new_n492), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n496), .A2(KEYINPUT93), .B1(G179), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n489), .A2(KEYINPUT92), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(new_n416), .A3(new_n492), .ZN(new_n501));
  INV_X1    g0301(.A(new_n485), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n495), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT93), .B1(new_n503), .B2(G169), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n251), .A2(new_n253), .A3(new_n206), .A4(G87), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT88), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n332), .A2(KEYINPUT88), .A3(new_n206), .A4(G87), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(new_n506), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT22), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT89), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT89), .A4(KEYINPUT22), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT23), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n385), .A3(G20), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT90), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n516), .B2(new_n385), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n517), .A2(new_n518), .B1(new_n521), .B2(G20), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n514), .A2(new_n515), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT24), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n298), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n514), .A2(KEYINPUT24), .A3(new_n515), .A4(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR3_X1    g0328(.A1(new_n289), .A2(KEYINPUT25), .A3(G107), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT25), .B1(new_n289), .B2(G107), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n205), .A2(G33), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n214), .A2(new_n289), .A3(new_n278), .A4(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n529), .B(new_n530), .C1(new_n533), .C2(new_n385), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n534), .A2(KEYINPUT91), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(KEYINPUT91), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n499), .A2(new_n505), .B1(new_n528), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n493), .A2(new_n324), .A3(new_n495), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(G200), .B2(new_n498), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n528), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n484), .A2(G270), .A3(new_n249), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT86), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT86), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n484), .A2(new_n545), .A3(G270), .A4(new_n249), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n497), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G283), .ZN(new_n548));
  INV_X1    g0348(.A(G97), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n206), .C1(G33), .C2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G116), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G20), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n279), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT20), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n550), .A2(KEYINPUT20), .A3(new_n279), .A4(new_n552), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n289), .A2(G116), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n532), .B2(G116), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n251), .A2(new_n253), .A3(G264), .A4(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n251), .A2(new_n253), .A3(G257), .A4(new_n336), .ZN(new_n562));
  INV_X1    g0362(.A(G303), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n332), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n416), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n547), .A2(new_n560), .A3(G179), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n544), .A2(new_n546), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n495), .A3(new_n565), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n276), .B1(new_n557), .B2(new_n559), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI211_X1 g0373(.A(new_n567), .B(KEYINPUT21), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n560), .B1(new_n569), .B2(G200), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n324), .B2(new_n569), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n251), .A2(new_n253), .A3(G244), .A4(new_n336), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n332), .A2(KEYINPUT4), .A3(G244), .A4(new_n336), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n332), .A2(G250), .A3(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n548), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n416), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n484), .A2(G257), .A3(new_n249), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n495), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n588), .A3(new_n392), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n284), .A2(new_n255), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n549), .A2(new_n385), .A3(KEYINPUT6), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT6), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G97), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n385), .A2(KEYINPUT82), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G107), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n591), .A2(new_n593), .A3(new_n595), .A4(new_n597), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n590), .B1(new_n601), .B2(G20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n443), .A2(G107), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n298), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n532), .A2(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n290), .A2(new_n549), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n589), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n587), .B1(new_n584), .B2(new_n416), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(G169), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT84), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT19), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n206), .B1(new_n338), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n220), .A2(new_n549), .A3(new_n385), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n251), .A2(new_n253), .A3(new_n206), .A4(G68), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n612), .B1(new_n281), .B2(new_n549), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n279), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n397), .A2(new_n290), .ZN(new_n620));
  INV_X1    g0420(.A(new_n397), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n532), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n249), .B(G250), .C1(G1), .C2(new_n271), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n267), .A2(new_n481), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n251), .A2(new_n253), .A3(G238), .A4(new_n336), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT85), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT85), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n332), .A2(new_n629), .A3(G238), .A4(new_n336), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n251), .A2(new_n253), .A3(G244), .A4(G1698), .ZN(new_n632));
  NAND2_X1  g0432(.A1(G33), .A2(G116), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n626), .B1(new_n636), .B2(new_n416), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n623), .B1(new_n637), .B2(new_n392), .ZN(new_n638));
  INV_X1    g0438(.A(new_n626), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n634), .B1(new_n630), .B2(new_n628), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(new_n249), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n276), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n619), .B(new_n620), .C1(new_n220), .C2(new_n533), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n641), .B2(G200), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n637), .A2(G190), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n638), .A2(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND4_X1   g0446(.A1(new_n591), .A2(new_n593), .A3(new_n595), .A4(new_n597), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n591), .A2(new_n593), .B1(new_n595), .B2(new_n597), .ZN(new_n648));
  OAI21_X1  g0448(.A(G20), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n590), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n385), .B1(new_n441), .B2(new_n442), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n279), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(new_n605), .A3(new_n606), .ZN(new_n654));
  INV_X1    g0454(.A(new_n610), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT84), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n654), .A2(new_n655), .A3(new_n656), .A4(new_n589), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n604), .A2(new_n607), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n585), .A2(new_n588), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G200), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT83), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n609), .A2(new_n661), .A3(G190), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(new_n609), .B2(G190), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n658), .B(new_n660), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n611), .A2(new_n646), .A3(new_n657), .A4(new_n664), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n480), .A2(new_n542), .A3(new_n578), .A4(new_n665), .ZN(G372));
  NAND2_X1  g0466(.A1(new_n638), .A2(new_n642), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n611), .A2(new_n657), .ZN(new_n669));
  XOR2_X1   g0469(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(new_n646), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n644), .A2(new_n645), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n654), .A2(new_n655), .A3(new_n589), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n668), .B1(new_n672), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n503), .A2(KEYINPUT93), .A3(G169), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n493), .A2(G179), .A3(new_n495), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n504), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n526), .A2(new_n527), .B1(new_n535), .B2(new_n536), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n575), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n541), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n665), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n480), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n309), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n473), .A2(new_n462), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT18), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n380), .A2(new_n408), .B1(new_n358), .B2(new_n374), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n465), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n327), .A2(new_n328), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n689), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n688), .A2(new_n695), .ZN(G369));
  NAND3_X1  g0496(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n542), .B1(new_n683), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n538), .A2(new_n702), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT96), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(KEYINPUT96), .A3(new_n705), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n560), .A2(new_n702), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT95), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n578), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n575), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n575), .A2(new_n702), .ZN(new_n717));
  INV_X1    g0517(.A(new_n708), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n706), .ZN(new_n719));
  INV_X1    g0519(.A(new_n538), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n702), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n716), .A2(new_n719), .A3(new_n722), .ZN(G399));
  INV_X1    g0523(.A(new_n209), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G41), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n614), .A2(G116), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(G1), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n212), .B2(new_n726), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n687), .A2(new_n703), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT100), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n702), .B1(new_n678), .B2(new_n686), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT100), .B1(new_n735), .B2(KEYINPUT29), .ZN(new_n736));
  INV_X1    g0536(.A(new_n686), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n671), .B1(new_n669), .B2(new_n646), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n675), .A2(new_n673), .A3(new_n676), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n667), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(KEYINPUT29), .B(new_n703), .C1(new_n737), .C2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n734), .A2(new_n736), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n542), .A2(new_n578), .A3(new_n665), .A4(new_n703), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n659), .A2(new_n641), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n568), .A2(G179), .A3(new_n495), .A4(new_n565), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT97), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n547), .A2(KEYINPUT97), .A3(G179), .A4(new_n565), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n744), .A2(new_n747), .A3(new_n493), .A4(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n569), .A2(new_n641), .A3(new_n392), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT98), .B1(new_n498), .B2(new_n609), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT98), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n503), .A2(new_n754), .A3(new_n659), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n749), .A2(new_n750), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT31), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n703), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n749), .A2(KEYINPUT99), .A3(new_n750), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT99), .B1(new_n749), .B2(new_n750), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n703), .B1(new_n765), .B2(new_n757), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n743), .B(new_n762), .C1(new_n766), .C2(KEYINPUT31), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G330), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n742), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n730), .B1(new_n770), .B2(G1), .ZN(G364));
  AND2_X1   g0571(.A1(new_n206), .A2(G13), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n205), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n725), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n715), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G330), .B2(new_n713), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n775), .B(KEYINPUT101), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n209), .A2(new_n332), .ZN(new_n779));
  INV_X1    g0579(.A(G355), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n780), .B1(G116), .B2(new_n209), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n724), .A2(new_n332), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n271), .B2(new_n213), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n245), .A2(G45), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(G20), .B1(KEYINPUT102), .B2(G169), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(KEYINPUT102), .A2(G169), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n214), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n778), .B1(new_n786), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n324), .A2(new_n377), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n206), .A2(G179), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n563), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  NOR2_X1   g0601(.A1(new_n206), .A2(new_n392), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n377), .A2(G190), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n798), .A2(new_n803), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n801), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n802), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n808), .A2(new_n324), .A3(G200), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n800), .B(new_n807), .C1(G322), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G179), .A2(G200), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G190), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G294), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n797), .A2(new_n802), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n332), .B1(new_n816), .B2(G326), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n808), .A2(G190), .A3(G200), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n811), .A2(G20), .A3(new_n324), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n818), .A2(G311), .B1(G329), .B2(new_n820), .ZN(new_n821));
  AND4_X1   g0621(.A1(new_n810), .A2(new_n814), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT104), .ZN(new_n824));
  INV_X1    g0624(.A(new_n818), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n825), .A2(new_n255), .B1(new_n286), .B2(new_n815), .ZN(new_n826));
  INV_X1    g0626(.A(new_n804), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n254), .B(new_n826), .C1(G68), .C2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT103), .B(KEYINPUT32), .Z(new_n829));
  INV_X1    g0629(.A(G159), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n830), .B2(new_n819), .ZN(new_n831));
  INV_X1    g0631(.A(new_n813), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n549), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n829), .A2(new_n830), .A3(new_n819), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n805), .A2(new_n385), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n799), .A2(new_n220), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(G58), .C2(new_n809), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n828), .A2(new_n831), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n823), .A2(KEYINPUT104), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n824), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n796), .B1(new_n841), .B2(new_n790), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n793), .B(KEYINPUT105), .Z(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n713), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n777), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G396));
  NAND2_X1  g0646(.A1(new_n406), .A2(new_n702), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n411), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n409), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n394), .A2(new_n407), .A3(new_n702), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n735), .B(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n775), .B1(new_n854), .B2(new_n768), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n768), .B2(new_n854), .ZN(new_n856));
  INV_X1    g0656(.A(new_n778), .ZN(new_n857));
  INV_X1    g0657(.A(new_n790), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n792), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT106), .Z(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n857), .B1(new_n255), .B2(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n816), .A2(G303), .B1(G311), .B2(new_n820), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n863), .B1(new_n385), .B2(new_n799), .C1(new_n825), .C2(new_n551), .ZN(new_n864));
  INV_X1    g0664(.A(new_n809), .ZN(new_n865));
  INV_X1    g0665(.A(G294), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n865), .A2(new_n866), .B1(new_n804), .B2(new_n806), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n254), .B1(new_n805), .B2(new_n220), .ZN(new_n868));
  NOR4_X1   g0668(.A1(new_n864), .A2(new_n833), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(G137), .A2(new_n816), .B1(new_n827), .B2(G150), .ZN(new_n870));
  INV_X1    g0670(.A(G143), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n870), .B1(new_n865), .B2(new_n871), .C1(new_n830), .C2(new_n825), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT34), .ZN(new_n873));
  INV_X1    g0673(.A(new_n805), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(G68), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n875), .B1(new_n286), .B2(new_n799), .C1(new_n422), .C2(new_n832), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n254), .B1(new_n820), .B2(G132), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n877), .A2(KEYINPUT107), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(KEYINPUT107), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n869), .B1(new_n873), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n850), .B1(new_n848), .B2(new_n409), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n862), .B1(new_n858), .B2(new_n881), .C1(new_n882), .C2(new_n792), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n856), .A2(new_n883), .ZN(G384));
  NAND2_X1  g0684(.A1(new_n215), .A2(G116), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n601), .B2(KEYINPUT35), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(KEYINPUT35), .B2(new_n601), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT36), .Z(new_n888));
  OR3_X1    g0688(.A1(new_n212), .A2(new_n255), .A3(new_n423), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n286), .A2(G68), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n205), .B(G13), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n457), .A2(KEYINPUT16), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n454), .B1(new_n895), .B2(new_n458), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n700), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n465), .B1(KEYINPUT18), .B2(new_n475), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(new_n478), .ZN(new_n900));
  INV_X1    g0700(.A(new_n700), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n467), .A2(new_n470), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n462), .A2(new_n421), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n475), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n473), .B2(new_n896), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n906), .B2(new_n897), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n893), .B1(new_n900), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n479), .A2(new_n897), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n907), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(KEYINPUT108), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n687), .A2(new_n703), .A3(new_n882), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n851), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT108), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n916), .B(new_n893), .C1(new_n900), .C2(new_n908), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n374), .A2(new_n702), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n375), .A2(new_n380), .A3(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n374), .B(new_n702), .C1(new_n358), .C2(new_n379), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n913), .A2(new_n915), .A3(new_n917), .A4(new_n921), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n691), .A2(new_n901), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT109), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n917), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n690), .B1(new_n462), .B2(new_n421), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n903), .B1(new_n927), .B2(new_n902), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n475), .A2(new_n903), .A3(new_n904), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n902), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n902), .B1(new_n691), .B2(new_n466), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n893), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n933), .A3(new_n912), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n375), .A2(new_n702), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT110), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT109), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n922), .A2(new_n941), .A3(new_n923), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n925), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n734), .A2(new_n736), .A3(new_n480), .A4(new_n741), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n944), .A2(new_n695), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n943), .B(new_n945), .Z(new_n946));
  INV_X1    g0746(.A(G330), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n852), .B1(new_n919), .B2(new_n920), .ZN(new_n948));
  INV_X1    g0748(.A(new_n764), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n749), .A2(KEYINPUT99), .A3(new_n750), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n757), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n702), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n760), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n766), .A2(KEYINPUT31), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n954), .A3(new_n743), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n913), .A2(new_n917), .A3(new_n948), .A4(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT40), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n743), .B1(new_n766), .B2(KEYINPUT31), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n952), .A2(new_n760), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n921), .A2(new_n882), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n957), .B1(new_n932), .B2(new_n912), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n956), .A2(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n480), .A2(new_n955), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n947), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n946), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n205), .B2(new_n772), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n946), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n892), .B1(new_n969), .B2(new_n970), .ZN(G367));
  INV_X1    g0771(.A(new_n717), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n707), .B2(new_n708), .ZN(new_n973));
  INV_X1    g0773(.A(new_n669), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n974), .B(new_n664), .C1(new_n658), .C2(new_n703), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n676), .A2(new_n703), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n538), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n702), .B1(new_n980), .B2(new_n974), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n978), .B2(KEYINPUT42), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n643), .A2(new_n702), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n646), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n667), .A2(new_n984), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n983), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n979), .A2(new_n982), .A3(new_n989), .A4(new_n988), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n716), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n977), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n994), .B(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n725), .B(KEYINPUT41), .Z(new_n999));
  INV_X1    g0799(.A(KEYINPUT44), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n977), .B1(KEYINPUT111), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n973), .B2(new_n721), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1000), .A2(KEYINPUT111), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT112), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1001), .B(new_n1004), .C1(new_n973), .C2(new_n721), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n719), .A2(new_n722), .A3(new_n977), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n719), .A2(KEYINPUT45), .A3(new_n722), .A4(new_n977), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1009), .A2(new_n716), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1014), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n995), .B1(new_n1016), .B2(new_n1008), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n707), .A2(new_n708), .A3(new_n972), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n719), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n714), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n719), .A2(new_n1018), .A3(new_n715), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1015), .A2(new_n1017), .A3(new_n770), .A4(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n999), .B1(new_n1024), .B2(new_n770), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n998), .B1(new_n1025), .B2(new_n774), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n794), .B1(new_n209), .B2(new_n397), .C1(new_n783), .C2(new_n237), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n805), .A2(new_n255), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n865), .A2(new_n282), .B1(new_n815), .B2(new_n871), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n799), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1028), .B(new_n1029), .C1(G58), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(G137), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n825), .A2(new_n286), .B1(new_n819), .B2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n254), .B(new_n1033), .C1(G159), .C2(new_n827), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n813), .A2(G68), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1031), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n820), .A2(G317), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n809), .A2(G303), .B1(new_n816), .B2(G311), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n332), .B1(new_n818), .B2(G283), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G294), .A2(new_n827), .B1(new_n874), .B2(G97), .ZN(new_n1041));
  AND4_X1   g0841(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n799), .A2(new_n551), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1043), .A2(KEYINPUT46), .B1(G107), .B2(new_n813), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(KEYINPUT46), .C2(new_n1043), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1037), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT47), .Z(new_n1048));
  OAI211_X1 g0848(.A(new_n778), .B(new_n1027), .C1(new_n1048), .C2(new_n858), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT114), .Z(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n843), .B2(new_n987), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1026), .A2(new_n1051), .ZN(G387));
  OR2_X1    g0852(.A1(new_n709), .A2(new_n843), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G303), .A2(new_n818), .B1(new_n809), .B2(G317), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G322), .A2(new_n816), .B1(new_n827), .B2(G311), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT48), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(KEYINPUT48), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1030), .A2(G294), .B1(new_n813), .B2(G283), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n254), .B1(new_n805), .B2(new_n551), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G326), .B2(new_n820), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n815), .A2(new_n830), .B1(new_n799), .B2(new_n255), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n254), .B(new_n1067), .C1(G97), .C2(new_n874), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n827), .A2(new_n395), .B1(new_n820), .B2(G150), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G50), .A2(new_n809), .B1(new_n818), .B2(G68), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n832), .A2(new_n397), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n858), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n727), .B(new_n271), .C1(new_n218), .C2(new_n255), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(KEYINPUT115), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT50), .B1(new_n280), .B2(G50), .ZN(new_n1077));
  OR3_X1    g0877(.A1(new_n280), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1075), .A2(KEYINPUT115), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n782), .B1(new_n1079), .B2(new_n1080), .C1(new_n234), .C2(new_n271), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(G107), .B2(new_n209), .C1(new_n727), .C2(new_n779), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n857), .B(new_n1074), .C1(new_n794), .C2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1023), .A2(new_n774), .B1(new_n1053), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1022), .A2(new_n769), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n770), .A2(new_n1021), .A3(new_n1020), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n725), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(new_n1087), .ZN(G393));
  AOI21_X1  g0888(.A(new_n716), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1016), .A2(new_n1008), .A3(new_n995), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n725), .A3(new_n1024), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n975), .A2(new_n793), .A3(new_n976), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT116), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n809), .A2(G311), .B1(new_n816), .B2(G317), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT52), .Z(new_n1096));
  AOI22_X1  g0896(.A1(new_n818), .A2(G294), .B1(G303), .B2(new_n827), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1030), .A2(G283), .B1(new_n820), .B2(G322), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n332), .B(new_n836), .C1(G116), .C2(new_n813), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n809), .A2(G159), .B1(new_n816), .B2(G150), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT51), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n286), .A2(new_n804), .B1(new_n799), .B2(new_n218), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n825), .A2(new_n280), .B1(new_n819), .B2(new_n871), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n332), .B1(new_n805), .B2(new_n220), .C1(new_n832), .C2(new_n255), .ZN(new_n1105));
  OR4_X1    g0905(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1100), .B1(new_n1107), .B2(KEYINPUT117), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT117), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n790), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n242), .A2(new_n782), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n795), .B1(G97), .B2(new_n724), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n857), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1094), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n774), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1092), .A2(new_n1117), .ZN(G390));
  AOI21_X1  g0918(.A(new_n850), .B1(new_n735), .B2(new_n882), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n921), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n938), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n926), .A2(new_n934), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n932), .A2(new_n912), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n740), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n702), .B1(new_n1124), .B2(new_n686), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n850), .B1(new_n1125), .B2(new_n849), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n938), .B(new_n1123), .C1(new_n1126), .C2(new_n1120), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n948), .A2(new_n955), .A3(G330), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n767), .A2(G330), .A3(new_n882), .A4(new_n921), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1122), .A2(new_n1127), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(new_n773), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n926), .A2(new_n791), .A3(new_n934), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n825), .A2(new_n549), .B1(new_n819), .B2(new_n866), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n837), .A2(new_n332), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n875), .C1(new_n385), .C2(new_n804), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1137), .B(new_n1139), .C1(G283), .C2(new_n816), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n809), .A2(G116), .B1(G77), .B2(new_n813), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT118), .Z(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT54), .B(G143), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n332), .B1(new_n825), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(G132), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n865), .A2(new_n1145), .B1(new_n804), .B2(new_n1032), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G159), .C2(new_n813), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n816), .A2(G128), .B1(G125), .B2(new_n820), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n286), .B2(new_n805), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT53), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n799), .B2(new_n282), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1030), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1149), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1140), .A2(new_n1142), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n778), .B1(new_n395), .B2(new_n860), .C1(new_n1154), .C2(new_n858), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT119), .Z(new_n1156));
  AOI21_X1  g0956(.A(new_n1135), .B1(new_n1136), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n480), .A2(new_n955), .A3(G330), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n944), .A2(new_n695), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n767), .A2(G330), .A3(new_n882), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1120), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1129), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n915), .ZN(new_n1163));
  OAI211_X1 g0963(.A(G330), .B(new_n882), .C1(new_n958), .C2(new_n959), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1120), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n1126), .A3(new_n1132), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1159), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1134), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1131), .A2(new_n1167), .A3(new_n1133), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n725), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1157), .A2(new_n1171), .ZN(G378));
  NAND2_X1  g0972(.A1(new_n317), .A2(new_n901), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n694), .A2(new_n309), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n329), .A2(new_n317), .A3(new_n901), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1174), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n791), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1145), .A2(new_n804), .B1(new_n799), .B2(new_n1143), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n809), .A2(G128), .B1(new_n816), .B2(G125), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n1032), .B2(new_n825), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G150), .C2(new_n813), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n250), .B(new_n270), .C1(new_n805), .C2(new_n830), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G124), .B2(new_n820), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n254), .A2(new_n270), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G77), .B2(new_n1030), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT120), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G116), .A2(new_n816), .B1(new_n827), .B2(G97), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n806), .B2(new_n819), .C1(new_n397), .C2(new_n825), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1035), .B1(new_n422), .B2(new_n805), .C1(new_n865), .C2(new_n385), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1194), .B(new_n286), .C1(G33), .C2(G41), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1193), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n790), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n775), .B1(new_n860), .B2(G50), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT121), .Z(new_n1207));
  NAND3_X1  g1007(.A1(new_n1183), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n940), .A2(new_n942), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n956), .A2(new_n957), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n947), .B1(new_n962), .B2(new_n963), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1182), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1181), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1210), .A2(new_n1214), .A3(new_n925), .A4(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1211), .A2(new_n1212), .A3(new_n1181), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1181), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n943), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1209), .B1(new_n1220), .B2(new_n774), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1159), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1170), .A2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1210), .A2(new_n925), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n943), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1223), .B(KEYINPUT57), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n725), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1221), .B1(new_n1227), .B2(new_n1228), .ZN(G375));
  NAND2_X1  g1029(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(new_n1222), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n999), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1168), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1230), .A2(new_n774), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n778), .B1(G68), .B2(new_n860), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n815), .A2(new_n866), .B1(new_n804), .B2(new_n551), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G107), .B2(new_n818), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT122), .Z(new_n1239));
  NOR3_X1   g1039(.A1(new_n1071), .A2(new_n332), .A3(new_n1028), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1030), .A2(G97), .B1(new_n820), .B2(G303), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n806), .C2(new_n865), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n865), .A2(new_n1032), .B1(new_n799), .B2(new_n830), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G132), .B2(new_n816), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n804), .A2(new_n1143), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G128), .B2(new_n820), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n332), .B1(new_n805), .B2(new_n422), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT124), .Z(new_n1248));
  NAND3_X1  g1048(.A1(new_n1244), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n818), .A2(G150), .B1(G50), .B2(new_n813), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT123), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1239), .A2(new_n1242), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1236), .B1(new_n1252), .B2(new_n790), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n921), .B2(new_n792), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1234), .A2(new_n1235), .A3(new_n1254), .ZN(G381));
  NAND3_X1  g1055(.A1(new_n1084), .A2(new_n1087), .A3(new_n845), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1256), .ZN(new_n1257));
  OR4_X1    g1057(.A1(G387), .A2(new_n1257), .A3(G375), .A4(G378), .ZN(G407));
  INV_X1    g1058(.A(G213), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(G343), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(G375), .A2(G378), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(KEYINPUT125), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(KEYINPUT125), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(G407), .A2(G213), .A3(new_n1264), .A4(new_n1265), .ZN(G409));
  NAND2_X1  g1066(.A1(G393), .A2(G396), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1256), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1092), .B2(new_n1117), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1092), .A2(new_n1117), .A3(new_n1268), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(new_n1026), .A3(new_n1051), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1271), .ZN(new_n1273));
  OAI21_X1  g1073(.A(G387), .B1(new_n1273), .B2(new_n1269), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1157), .A2(new_n1171), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1216), .A2(KEYINPUT126), .A3(new_n1219), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT126), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n773), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1220), .A2(new_n1233), .A3(new_n1223), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1208), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1276), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1221), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1260), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1235), .A2(new_n1254), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1232), .B1(new_n1167), .B2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1167), .A2(new_n1286), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n726), .B1(new_n1288), .B2(new_n1231), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1285), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(G384), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1290), .A2(G384), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT62), .B1(new_n1284), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1261), .ZN(new_n1298));
  AOI211_X1 g1098(.A(KEYINPUT127), .B(new_n1260), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1294), .A2(KEYINPUT62), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1295), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(G2897), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1261), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1293), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1305), .B2(new_n1291), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1294), .A2(new_n1304), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1275), .B1(new_n1302), .B2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1284), .B1(new_n1308), .B2(new_n1307), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT63), .B1(new_n1284), .B2(new_n1294), .ZN(new_n1315));
  NOR4_X1   g1115(.A1(new_n1314), .A2(new_n1315), .A3(KEYINPUT61), .A4(new_n1275), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1294), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1313), .A2(new_n1318), .ZN(G405));
  AND2_X1   g1119(.A1(G375), .A2(new_n1276), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1283), .ZN(new_n1321));
  OR3_X1    g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1294), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1294), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(new_n1275), .ZN(G402));
endmodule


