

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n659), .A2(G651), .ZN(n663) );
  NAND2_X1 U550 ( .A1(n524), .A2(n521), .ZN(n908) );
  NAND2_X2 U551 ( .A1(n793), .A2(n795), .ZN(n747) );
  XNOR2_X1 U552 ( .A(n706), .B(n539), .ZN(n538) );
  OR2_X1 U553 ( .A1(G2105), .A2(n698), .ZN(n699) );
  INV_X1 U554 ( .A(KEYINPUT27), .ZN(n539) );
  NAND2_X1 U555 ( .A1(n533), .A2(n532), .ZN(n531) );
  NOR2_X1 U556 ( .A1(n763), .A2(n520), .ZN(n532) );
  INV_X1 U557 ( .A(KEYINPUT103), .ZN(n530) );
  NAND2_X1 U558 ( .A1(G2105), .A2(KEYINPUT17), .ZN(n522) );
  NAND2_X1 U559 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n523) );
  NOR2_X1 U560 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n526) );
  NOR2_X1 U561 ( .A1(n771), .A2(n787), .ZN(n541) );
  NOR2_X2 U562 ( .A1(n704), .A2(n527), .ZN(n793) );
  NAND2_X1 U563 ( .A1(n528), .A2(G40), .ZN(n527) );
  INV_X1 U564 ( .A(n703), .ZN(n528) );
  OR2_X1 U565 ( .A1(n704), .A2(n703), .ZN(n529) );
  NOR2_X1 U566 ( .A1(n536), .A2(n534), .ZN(n726) );
  NAND2_X1 U567 ( .A1(n537), .A2(n518), .ZN(n536) );
  AND2_X1 U568 ( .A1(n535), .A2(n707), .ZN(n534) );
  NOR2_X1 U569 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U570 ( .A(n531), .B(n530), .ZN(n764) );
  NAND2_X1 U571 ( .A1(n526), .A2(n525), .ZN(n524) );
  AND2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n521) );
  INV_X1 U573 ( .A(G2105), .ZN(n525) );
  XNOR2_X1 U574 ( .A(n699), .B(KEYINPUT23), .ZN(n700) );
  INV_X1 U575 ( .A(KEYINPUT110), .ZN(n791) );
  AND2_X1 U576 ( .A1(n517), .A2(n540), .ZN(n792) );
  XNOR2_X1 U577 ( .A(n541), .B(KEYINPUT109), .ZN(n540) );
  XNOR2_X1 U578 ( .A(n953), .B(G160), .ZN(n921) );
  AND2_X1 U579 ( .A1(n788), .A2(n519), .ZN(n517) );
  NAND2_X1 U580 ( .A1(n747), .A2(G1956), .ZN(n518) );
  OR2_X1 U581 ( .A1(n790), .A2(n789), .ZN(n519) );
  AND2_X1 U582 ( .A1(G8), .A2(n762), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n529), .B(G2084), .ZN(n943) );
  INV_X1 U584 ( .A(n529), .ZN(G160) );
  NAND2_X1 U585 ( .A1(n760), .A2(n761), .ZN(n533) );
  INV_X1 U586 ( .A(n538), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n538), .A2(KEYINPUT99), .ZN(n537) );
  NAND2_X1 U588 ( .A1(n705), .A2(G2072), .ZN(n706) );
  INV_X1 U589 ( .A(KEYINPUT28), .ZN(n708) );
  XNOR2_X1 U590 ( .A(KEYINPUT102), .B(KEYINPUT30), .ZN(n741) );
  XNOR2_X1 U591 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U592 ( .A1(n745), .A2(n744), .ZN(n746) );
  INV_X1 U593 ( .A(KEYINPUT104), .ZN(n756) );
  XOR2_X1 U594 ( .A(KEYINPUT15), .B(n600), .Z(n996) );
  NOR2_X1 U595 ( .A1(G2105), .A2(n544), .ZN(n909) );
  NAND2_X1 U596 ( .A1(G138), .A2(n908), .ZN(n543) );
  INV_X1 U597 ( .A(G2104), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G102), .A2(n909), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n548) );
  AND2_X1 U600 ( .A1(n544), .A2(G2105), .ZN(n903) );
  NAND2_X1 U601 ( .A1(G126), .A2(n903), .ZN(n546) );
  AND2_X1 U602 ( .A1(G2105), .A2(G2104), .ZN(n904) );
  NAND2_X1 U603 ( .A1(G114), .A2(n904), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U605 ( .A1(n548), .A2(n547), .ZN(G164) );
  NOR2_X1 U606 ( .A1(G543), .A2(G651), .ZN(n649) );
  NAND2_X1 U607 ( .A1(n649), .A2(G85), .ZN(n550) );
  XOR2_X1 U608 ( .A(KEYINPUT0), .B(G543), .Z(n659) );
  XNOR2_X1 U609 ( .A(KEYINPUT67), .B(G651), .ZN(n551) );
  NOR2_X1 U610 ( .A1(n659), .A2(n551), .ZN(n652) );
  NAND2_X1 U611 ( .A1(G72), .A2(n652), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n663), .A2(G47), .ZN(n554) );
  NOR2_X1 U614 ( .A1(G543), .A2(n551), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT1), .B(n552), .Z(n594) );
  BUF_X1 U616 ( .A(n594), .Z(n662) );
  NAND2_X1 U617 ( .A1(G60), .A2(n662), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U619 ( .A1(n556), .A2(n555), .ZN(G290) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  NAND2_X1 U624 ( .A1(G89), .A2(n649), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT4), .B(n557), .Z(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(KEYINPUT75), .ZN(n560) );
  NAND2_X1 U627 ( .A1(G76), .A2(n652), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(KEYINPUT5), .B(n561), .ZN(n569) );
  XNOR2_X1 U630 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n663), .A2(G51), .ZN(n562) );
  XNOR2_X1 U632 ( .A(n562), .B(KEYINPUT76), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G63), .A2(n662), .ZN(n563) );
  NAND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U635 ( .A(n565), .B(KEYINPUT6), .ZN(n566) );
  XNOR2_X1 U636 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(KEYINPUT7), .B(n570), .ZN(G168) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U642 ( .A(G223), .ZN(n857) );
  NAND2_X1 U643 ( .A1(n857), .A2(G567), .ZN(n572) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  XOR2_X1 U645 ( .A(G860), .B(KEYINPUT72), .Z(n614) );
  NAND2_X1 U646 ( .A1(n649), .A2(G81), .ZN(n573) );
  XNOR2_X1 U647 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U648 ( .A1(G68), .A2(n652), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U650 ( .A(KEYINPUT13), .B(n576), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n662), .A2(G56), .ZN(n577) );
  XOR2_X1 U652 ( .A(KEYINPUT14), .B(n577), .Z(n580) );
  NAND2_X1 U653 ( .A1(G43), .A2(n663), .ZN(n578) );
  XNOR2_X1 U654 ( .A(KEYINPUT71), .B(n578), .ZN(n579) );
  NOR2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n992) );
  OR2_X1 U657 ( .A1(n614), .A2(n992), .ZN(G153) );
  NAND2_X1 U658 ( .A1(n663), .A2(G52), .ZN(n584) );
  NAND2_X1 U659 ( .A1(G64), .A2(n662), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n649), .A2(G90), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT68), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G77), .A2(n652), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U665 ( .A(KEYINPUT9), .B(n588), .Z(n589) );
  NOR2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U667 ( .A(KEYINPUT69), .B(n591), .Z(G171) );
  INV_X1 U668 ( .A(G171), .ZN(G301) );
  NAND2_X1 U669 ( .A1(n663), .A2(G54), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n649), .A2(G92), .ZN(n593) );
  NAND2_X1 U671 ( .A1(G79), .A2(n652), .ZN(n592) );
  NAND2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U673 ( .A1(G66), .A2(n594), .ZN(n595) );
  XNOR2_X1 U674 ( .A(KEYINPUT73), .B(n595), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U677 ( .A1(G868), .A2(n996), .ZN(n602) );
  INV_X1 U678 ( .A(G868), .ZN(n611) );
  NOR2_X1 U679 ( .A1(n611), .A2(G301), .ZN(n601) );
  NOR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U681 ( .A(KEYINPUT74), .B(n603), .ZN(G284) );
  NAND2_X1 U682 ( .A1(n649), .A2(G91), .ZN(n605) );
  NAND2_X1 U683 ( .A1(G65), .A2(n662), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n652), .A2(G78), .ZN(n606) );
  XOR2_X1 U686 ( .A(KEYINPUT70), .B(n606), .Z(n607) );
  NOR2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n663), .A2(G53), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(G299) );
  NOR2_X1 U690 ( .A1(G286), .A2(n611), .ZN(n613) );
  NOR2_X1 U691 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n614), .A2(G559), .ZN(n615) );
  INV_X1 U694 ( .A(n996), .ZN(n926) );
  NAND2_X1 U695 ( .A1(n615), .A2(n926), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n616), .B(KEYINPUT16), .ZN(n617) );
  XOR2_X1 U697 ( .A(KEYINPUT79), .B(n617), .Z(G148) );
  NOR2_X1 U698 ( .A1(G868), .A2(n992), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G868), .A2(n926), .ZN(n618) );
  NOR2_X1 U700 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U701 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U702 ( .A1(G123), .A2(n903), .ZN(n621) );
  XNOR2_X1 U703 ( .A(n621), .B(KEYINPUT80), .ZN(n622) );
  XNOR2_X1 U704 ( .A(n622), .B(KEYINPUT18), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G111), .A2(n904), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G135), .A2(n908), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G99), .A2(n909), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U711 ( .A(KEYINPUT81), .B(n629), .Z(n945) );
  XNOR2_X1 U712 ( .A(G2096), .B(n945), .ZN(n631) );
  INV_X1 U713 ( .A(G2100), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(G156) );
  NAND2_X1 U715 ( .A1(G559), .A2(n926), .ZN(n632) );
  XNOR2_X1 U716 ( .A(n632), .B(KEYINPUT82), .ZN(n676) );
  XNOR2_X1 U717 ( .A(n676), .B(n992), .ZN(n633) );
  NOR2_X1 U718 ( .A1(n633), .A2(G860), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n649), .A2(G93), .ZN(n635) );
  NAND2_X1 U720 ( .A1(G80), .A2(n652), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n663), .A2(G55), .ZN(n637) );
  NAND2_X1 U723 ( .A1(G67), .A2(n662), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n678) );
  XNOR2_X1 U726 ( .A(n640), .B(n678), .ZN(G145) );
  NAND2_X1 U727 ( .A1(G86), .A2(n649), .ZN(n641) );
  XNOR2_X1 U728 ( .A(n641), .B(KEYINPUT86), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n663), .A2(G48), .ZN(n643) );
  NAND2_X1 U730 ( .A1(G61), .A2(n662), .ZN(n642) );
  NAND2_X1 U731 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n652), .A2(G73), .ZN(n644) );
  XOR2_X1 U733 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U734 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U735 ( .A1(n648), .A2(n647), .ZN(G305) );
  NAND2_X1 U736 ( .A1(n663), .A2(G50), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n649), .A2(G88), .ZN(n651) );
  NAND2_X1 U738 ( .A1(G62), .A2(n662), .ZN(n650) );
  NAND2_X1 U739 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U740 ( .A1(G75), .A2(n652), .ZN(n653) );
  XNOR2_X1 U741 ( .A(KEYINPUT87), .B(n653), .ZN(n654) );
  NOR2_X1 U742 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U743 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U744 ( .A(KEYINPUT88), .B(n658), .Z(G166) );
  NAND2_X1 U745 ( .A1(n659), .A2(G87), .ZN(n660) );
  XOR2_X1 U746 ( .A(KEYINPUT84), .B(n660), .Z(n661) );
  NOR2_X1 U747 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n663), .A2(G49), .ZN(n664) );
  NAND2_X1 U749 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U750 ( .A1(G74), .A2(G651), .ZN(n666) );
  XNOR2_X1 U751 ( .A(KEYINPUT83), .B(n666), .ZN(n667) );
  NOR2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U753 ( .A(KEYINPUT85), .B(n669), .ZN(G288) );
  XOR2_X1 U754 ( .A(G166), .B(G288), .Z(n670) );
  XNOR2_X1 U755 ( .A(G305), .B(n670), .ZN(n673) );
  XNOR2_X1 U756 ( .A(KEYINPUT19), .B(G290), .ZN(n671) );
  XNOR2_X1 U757 ( .A(n671), .B(n992), .ZN(n672) );
  XOR2_X1 U758 ( .A(n673), .B(n672), .Z(n675) );
  INV_X1 U759 ( .A(G299), .ZN(n725) );
  XNOR2_X1 U760 ( .A(n725), .B(n678), .ZN(n674) );
  XNOR2_X1 U761 ( .A(n675), .B(n674), .ZN(n925) );
  XNOR2_X1 U762 ( .A(n676), .B(n925), .ZN(n677) );
  NAND2_X1 U763 ( .A1(n677), .A2(G868), .ZN(n680) );
  OR2_X1 U764 ( .A1(G868), .A2(n678), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n680), .A2(n679), .ZN(G295) );
  XNOR2_X1 U766 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n683) );
  NAND2_X1 U767 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XNOR2_X1 U768 ( .A(n681), .B(KEYINPUT89), .ZN(n682) );
  XNOR2_X1 U769 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U770 ( .A1(G2090), .A2(n684), .ZN(n685) );
  XNOR2_X1 U771 ( .A(KEYINPUT21), .B(n685), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n686), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U773 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U774 ( .A1(G220), .A2(G219), .ZN(n687) );
  XOR2_X1 U775 ( .A(KEYINPUT22), .B(n687), .Z(n688) );
  NOR2_X1 U776 ( .A1(G218), .A2(n688), .ZN(n689) );
  NAND2_X1 U777 ( .A1(G96), .A2(n689), .ZN(n862) );
  NAND2_X1 U778 ( .A1(n862), .A2(G2106), .ZN(n693) );
  NAND2_X1 U779 ( .A1(G69), .A2(G120), .ZN(n690) );
  NOR2_X1 U780 ( .A1(G237), .A2(n690), .ZN(n691) );
  NAND2_X1 U781 ( .A1(G108), .A2(n691), .ZN(n863) );
  NAND2_X1 U782 ( .A1(n863), .A2(G567), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n864) );
  NAND2_X1 U784 ( .A1(G661), .A2(G483), .ZN(n694) );
  NOR2_X1 U785 ( .A1(n864), .A2(n694), .ZN(n861) );
  NAND2_X1 U786 ( .A1(n861), .A2(G36), .ZN(G176) );
  XNOR2_X1 U787 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  NAND2_X1 U788 ( .A1(n908), .A2(G137), .ZN(n696) );
  NAND2_X1 U789 ( .A1(G113), .A2(n904), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U791 ( .A(n697), .B(KEYINPUT66), .ZN(n704) );
  NAND2_X1 U792 ( .A1(G2104), .A2(G101), .ZN(n698) );
  XNOR2_X1 U793 ( .A(n700), .B(KEYINPUT65), .ZN(n702) );
  NAND2_X1 U794 ( .A1(G125), .A2(n903), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X2 U796 ( .A1(G164), .A2(G1384), .ZN(n795) );
  INV_X1 U797 ( .A(n747), .ZN(n705) );
  INV_X1 U798 ( .A(KEYINPUT99), .ZN(n707) );
  NOR2_X1 U799 ( .A1(n726), .A2(n725), .ZN(n709) );
  XNOR2_X1 U800 ( .A(n709), .B(n708), .ZN(n730) );
  XNOR2_X1 U801 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n716) );
  NOR2_X1 U802 ( .A1(G1996), .A2(n716), .ZN(n710) );
  NOR2_X1 U803 ( .A1(n992), .A2(n710), .ZN(n714) );
  NAND2_X1 U804 ( .A1(G1348), .A2(n747), .ZN(n712) );
  INV_X1 U805 ( .A(n747), .ZN(n733) );
  NAND2_X1 U806 ( .A1(G2067), .A2(n733), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n722) );
  NAND2_X1 U808 ( .A1(n996), .A2(n722), .ZN(n713) );
  NAND2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n721) );
  INV_X1 U810 ( .A(G1341), .ZN(n1011) );
  NAND2_X1 U811 ( .A1(n1011), .A2(n716), .ZN(n715) );
  NAND2_X1 U812 ( .A1(n715), .A2(n747), .ZN(n719) );
  INV_X1 U813 ( .A(G1996), .ZN(n966) );
  NOR2_X1 U814 ( .A1(n966), .A2(n747), .ZN(n717) );
  NAND2_X1 U815 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U816 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U817 ( .A1(n721), .A2(n720), .ZN(n724) );
  NOR2_X1 U818 ( .A1(n722), .A2(n996), .ZN(n723) );
  NOR2_X1 U819 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n732) );
  XNOR2_X1 U823 ( .A(KEYINPUT100), .B(KEYINPUT29), .ZN(n731) );
  XNOR2_X1 U824 ( .A(n732), .B(n731), .ZN(n737) );
  XNOR2_X1 U825 ( .A(G2078), .B(KEYINPUT25), .ZN(n965) );
  NOR2_X1 U826 ( .A1(n747), .A2(n965), .ZN(n735) );
  INV_X1 U827 ( .A(G1961), .ZN(n993) );
  NOR2_X1 U828 ( .A1(n733), .A2(n993), .ZN(n734) );
  NOR2_X1 U829 ( .A1(n735), .A2(n734), .ZN(n739) );
  AND2_X1 U830 ( .A1(G171), .A2(n739), .ZN(n736) );
  XNOR2_X1 U831 ( .A(n738), .B(KEYINPUT101), .ZN(n760) );
  NOR2_X1 U832 ( .A1(G171), .A2(n739), .ZN(n745) );
  NAND2_X1 U833 ( .A1(G8), .A2(n747), .ZN(n770) );
  NOR2_X1 U834 ( .A1(G1966), .A2(n770), .ZN(n763) );
  NOR2_X1 U835 ( .A1(G2084), .A2(n747), .ZN(n762) );
  NOR2_X1 U836 ( .A1(n763), .A2(n762), .ZN(n740) );
  NAND2_X1 U837 ( .A1(G8), .A2(n740), .ZN(n742) );
  NOR2_X1 U838 ( .A1(G168), .A2(n743), .ZN(n744) );
  XOR2_X1 U839 ( .A(KEYINPUT31), .B(n746), .Z(n761) );
  NOR2_X1 U840 ( .A1(G1971), .A2(n770), .ZN(n749) );
  NOR2_X1 U841 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n750), .A2(G303), .ZN(n752) );
  AND2_X1 U844 ( .A1(n761), .A2(n752), .ZN(n751) );
  NAND2_X1 U845 ( .A1(n760), .A2(n751), .ZN(n755) );
  INV_X1 U846 ( .A(n752), .ZN(n753) );
  OR2_X1 U847 ( .A1(n753), .A2(G286), .ZN(n754) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n757) );
  XNOR2_X1 U849 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n758), .A2(G8), .ZN(n759) );
  XNOR2_X1 U851 ( .A(n759), .B(KEYINPUT32), .ZN(n765) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U853 ( .A(n766), .B(KEYINPUT105), .ZN(n772) );
  NOR2_X1 U854 ( .A1(G303), .A2(G2090), .ZN(n767) );
  NAND2_X1 U855 ( .A1(G8), .A2(n767), .ZN(n768) );
  XOR2_X1 U856 ( .A(KEYINPUT108), .B(n768), .Z(n769) );
  NOR2_X1 U857 ( .A1(n772), .A2(n769), .ZN(n771) );
  INV_X1 U858 ( .A(n770), .ZN(n787) );
  INV_X1 U859 ( .A(n772), .ZN(n774) );
  NOR2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n777) );
  NOR2_X1 U861 ( .A1(G303), .A2(G1971), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n777), .A2(n773), .ZN(n1008) );
  NAND2_X1 U863 ( .A1(n774), .A2(n1008), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G288), .A2(G1976), .ZN(n775) );
  XOR2_X1 U865 ( .A(KEYINPUT106), .B(n775), .Z(n991) );
  XNOR2_X1 U866 ( .A(KEYINPUT107), .B(G1981), .ZN(n776) );
  XNOR2_X1 U867 ( .A(n776), .B(G305), .ZN(n1001) );
  AND2_X1 U868 ( .A1(n787), .A2(n777), .ZN(n778) );
  NAND2_X1 U869 ( .A1(KEYINPUT33), .A2(n778), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n1001), .A2(n779), .ZN(n789) );
  NOR2_X1 U871 ( .A1(n991), .A2(n789), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n785) );
  NOR2_X1 U873 ( .A1(G1981), .A2(G305), .ZN(n782) );
  XOR2_X1 U874 ( .A(n782), .B(KEYINPUT24), .Z(n783) );
  XNOR2_X1 U875 ( .A(KEYINPUT98), .B(n783), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  INV_X1 U878 ( .A(KEYINPUT33), .ZN(n790) );
  XNOR2_X1 U879 ( .A(n792), .B(n791), .ZN(n830) );
  XNOR2_X1 U880 ( .A(G1986), .B(G290), .ZN(n987) );
  INV_X1 U881 ( .A(n793), .ZN(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n841) );
  NAND2_X1 U883 ( .A1(n987), .A2(n841), .ZN(n796) );
  XNOR2_X1 U884 ( .A(n796), .B(KEYINPUT92), .ZN(n809) );
  XNOR2_X1 U885 ( .A(KEYINPUT37), .B(G2067), .ZN(n839) );
  NAND2_X1 U886 ( .A1(G140), .A2(n908), .ZN(n799) );
  NAND2_X1 U887 ( .A1(n909), .A2(G104), .ZN(n797) );
  XOR2_X1 U888 ( .A(KEYINPUT93), .B(n797), .Z(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n802) );
  XOR2_X1 U890 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n800) );
  XNOR2_X1 U891 ( .A(KEYINPUT34), .B(n800), .ZN(n801) );
  XNOR2_X1 U892 ( .A(n802), .B(n801), .ZN(n807) );
  NAND2_X1 U893 ( .A1(G128), .A2(n903), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G116), .A2(n904), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U896 ( .A(KEYINPUT35), .B(n805), .Z(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U898 ( .A(KEYINPUT36), .B(n808), .ZN(n922) );
  NOR2_X1 U899 ( .A1(n839), .A2(n922), .ZN(n942) );
  NAND2_X1 U900 ( .A1(n841), .A2(n942), .ZN(n837) );
  NAND2_X1 U901 ( .A1(n809), .A2(n837), .ZN(n828) );
  NAND2_X1 U902 ( .A1(G119), .A2(n903), .ZN(n811) );
  NAND2_X1 U903 ( .A1(G107), .A2(n904), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n815) );
  NAND2_X1 U905 ( .A1(G131), .A2(n908), .ZN(n813) );
  NAND2_X1 U906 ( .A1(G95), .A2(n909), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n899) );
  INV_X1 U909 ( .A(G1991), .ZN(n963) );
  NOR2_X1 U910 ( .A1(n899), .A2(n963), .ZN(n825) );
  NAND2_X1 U911 ( .A1(G141), .A2(n908), .ZN(n816) );
  XNOR2_X1 U912 ( .A(n816), .B(KEYINPUT96), .ZN(n823) );
  NAND2_X1 U913 ( .A1(G129), .A2(n903), .ZN(n818) );
  NAND2_X1 U914 ( .A1(G117), .A2(n904), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n909), .A2(G105), .ZN(n819) );
  XOR2_X1 U917 ( .A(KEYINPUT38), .B(n819), .Z(n820) );
  NOR2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n900) );
  AND2_X1 U920 ( .A1(n900), .A2(G1996), .ZN(n824) );
  NOR2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n940) );
  INV_X1 U922 ( .A(n841), .ZN(n826) );
  NOR2_X1 U923 ( .A1(n940), .A2(n826), .ZN(n833) );
  XOR2_X1 U924 ( .A(KEYINPUT97), .B(n833), .Z(n827) );
  NOR2_X1 U925 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n844) );
  NOR2_X1 U927 ( .A1(G1996), .A2(n900), .ZN(n937) );
  NOR2_X1 U928 ( .A1(G1986), .A2(G290), .ZN(n831) );
  AND2_X1 U929 ( .A1(n963), .A2(n899), .ZN(n941) );
  NOR2_X1 U930 ( .A1(n831), .A2(n941), .ZN(n832) );
  NOR2_X1 U931 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U932 ( .A(KEYINPUT111), .B(n834), .Z(n835) );
  NOR2_X1 U933 ( .A1(n937), .A2(n835), .ZN(n836) );
  XNOR2_X1 U934 ( .A(KEYINPUT39), .B(n836), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n838), .A2(n837), .ZN(n840) );
  NAND2_X1 U936 ( .A1(n839), .A2(n922), .ZN(n951) );
  NAND2_X1 U937 ( .A1(n840), .A2(n951), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U939 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U940 ( .A(n845), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U941 ( .A(G2446), .B(G2451), .ZN(n855) );
  XOR2_X1 U942 ( .A(G2430), .B(KEYINPUT113), .Z(n847) );
  XNOR2_X1 U943 ( .A(G2454), .B(G2435), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U945 ( .A(G2438), .B(KEYINPUT112), .Z(n849) );
  XNOR2_X1 U946 ( .A(G1341), .B(G1348), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U948 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U949 ( .A(G2427), .B(G2443), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(n856) );
  NAND2_X1 U952 ( .A1(n856), .A2(G14), .ZN(n930) );
  XOR2_X1 U953 ( .A(KEYINPUT114), .B(n930), .Z(G401) );
  NAND2_X1 U954 ( .A1(G2106), .A2(n857), .ZN(G217) );
  AND2_X1 U955 ( .A1(G15), .A2(G2), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G661), .A2(n858), .ZN(G259) );
  NAND2_X1 U957 ( .A1(G3), .A2(G1), .ZN(n859) );
  XOR2_X1 U958 ( .A(KEYINPUT115), .B(n859), .Z(n860) );
  NAND2_X1 U959 ( .A1(n861), .A2(n860), .ZN(G188) );
  INV_X1 U961 ( .A(G120), .ZN(G236) );
  INV_X1 U962 ( .A(G96), .ZN(G221) );
  INV_X1 U963 ( .A(G69), .ZN(G235) );
  NOR2_X1 U964 ( .A1(n863), .A2(n862), .ZN(G325) );
  INV_X1 U965 ( .A(G325), .ZN(G261) );
  INV_X1 U966 ( .A(n864), .ZN(G319) );
  XOR2_X1 U967 ( .A(G2096), .B(KEYINPUT43), .Z(n866) );
  XNOR2_X1 U968 ( .A(G2072), .B(G2678), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U970 ( .A(n867), .B(KEYINPUT116), .Z(n869) );
  XNOR2_X1 U971 ( .A(G2067), .B(G2090), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U973 ( .A(KEYINPUT42), .B(G2100), .Z(n871) );
  XNOR2_X1 U974 ( .A(G2078), .B(G2084), .ZN(n870) );
  XNOR2_X1 U975 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U976 ( .A(n873), .B(n872), .ZN(G227) );
  XOR2_X1 U977 ( .A(G1976), .B(G1961), .Z(n875) );
  XNOR2_X1 U978 ( .A(G1986), .B(G1966), .ZN(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U980 ( .A(n876), .B(G2474), .Z(n878) );
  XNOR2_X1 U981 ( .A(G1956), .B(G1971), .ZN(n877) );
  XNOR2_X1 U982 ( .A(n878), .B(n877), .ZN(n882) );
  XOR2_X1 U983 ( .A(KEYINPUT41), .B(G1981), .Z(n880) );
  XNOR2_X1 U984 ( .A(G1996), .B(G1991), .ZN(n879) );
  XNOR2_X1 U985 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U986 ( .A(n882), .B(n881), .ZN(G229) );
  NAND2_X1 U987 ( .A1(G124), .A2(n903), .ZN(n883) );
  XNOR2_X1 U988 ( .A(n883), .B(KEYINPUT44), .ZN(n886) );
  NAND2_X1 U989 ( .A1(G100), .A2(n909), .ZN(n884) );
  XOR2_X1 U990 ( .A(KEYINPUT117), .B(n884), .Z(n885) );
  NAND2_X1 U991 ( .A1(n886), .A2(n885), .ZN(n890) );
  NAND2_X1 U992 ( .A1(G136), .A2(n908), .ZN(n888) );
  NAND2_X1 U993 ( .A1(G112), .A2(n904), .ZN(n887) );
  NAND2_X1 U994 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U995 ( .A1(n890), .A2(n889), .ZN(G162) );
  NAND2_X1 U996 ( .A1(G139), .A2(n908), .ZN(n892) );
  NAND2_X1 U997 ( .A1(G103), .A2(n909), .ZN(n891) );
  NAND2_X1 U998 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U999 ( .A(KEYINPUT119), .B(n893), .Z(n898) );
  NAND2_X1 U1000 ( .A1(G127), .A2(n903), .ZN(n895) );
  NAND2_X1 U1001 ( .A1(G115), .A2(n904), .ZN(n894) );
  NAND2_X1 U1002 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U1003 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U1004 ( .A1(n898), .A2(n897), .ZN(n953) );
  XOR2_X1 U1005 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n902) );
  XOR2_X1 U1006 ( .A(n900), .B(n899), .Z(n901) );
  XNOR2_X1 U1007 ( .A(n902), .B(n901), .ZN(n916) );
  NAND2_X1 U1008 ( .A1(G130), .A2(n903), .ZN(n906) );
  NAND2_X1 U1009 ( .A1(G118), .A2(n904), .ZN(n905) );
  NAND2_X1 U1010 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1011 ( .A(KEYINPUT118), .B(n907), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(G142), .A2(n908), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(G106), .A2(n909), .ZN(n910) );
  NAND2_X1 U1014 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1015 ( .A(n912), .B(KEYINPUT45), .Z(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1017 ( .A(n916), .B(n915), .Z(n917) );
  XOR2_X1 U1018 ( .A(n917), .B(G162), .Z(n919) );
  XNOR2_X1 U1019 ( .A(G164), .B(n945), .ZN(n918) );
  XNOR2_X1 U1020 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(n921), .B(n920), .ZN(n923) );
  XOR2_X1 U1022 ( .A(n923), .B(n922), .Z(n924) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n924), .ZN(G395) );
  XOR2_X1 U1024 ( .A(n925), .B(G286), .Z(n928) );
  XNOR2_X1 U1025 ( .A(G171), .B(n926), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(n928), .B(n927), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(G37), .A2(n929), .ZN(G397) );
  NAND2_X1 U1028 ( .A1(G319), .A2(n930), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(G227), .A2(G229), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(KEYINPUT49), .B(n931), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(G395), .A2(G397), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(G225) );
  INV_X1 U1034 ( .A(G225), .ZN(G308) );
  INV_X1 U1035 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1038 ( .A(KEYINPUT51), .B(n938), .Z(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n950) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT120), .B(n943), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1044 ( .A(KEYINPUT121), .B(n948), .Z(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n958) );
  XOR2_X1 U1047 ( .A(G2072), .B(n953), .Z(n955) );
  XOR2_X1 U1048 ( .A(G164), .B(G2078), .Z(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1050 ( .A(KEYINPUT50), .B(n956), .Z(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(KEYINPUT52), .B(n959), .ZN(n961) );
  INV_X1 U1053 ( .A(KEYINPUT55), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n962), .A2(G29), .ZN(n1042) );
  XNOR2_X1 U1056 ( .A(G29), .B(KEYINPUT123), .ZN(n984) );
  XNOR2_X1 U1057 ( .A(G25), .B(n963), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(G28), .ZN(n971) );
  XOR2_X1 U1059 ( .A(n965), .B(G27), .Z(n968) );
  XOR2_X1 U1060 ( .A(n966), .B(G32), .Z(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1062 ( .A(KEYINPUT122), .B(n969), .Z(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(G2067), .B(G26), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(G33), .B(G2072), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT53), .ZN(n979) );
  XOR2_X1 U1069 ( .A(G2084), .B(G34), .Z(n977) );
  XNOR2_X1 U1070 ( .A(KEYINPUT54), .B(n977), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G35), .B(G2090), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(KEYINPUT55), .B(n982), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(G11), .A2(n985), .ZN(n1040) );
  XNOR2_X1 U1077 ( .A(G16), .B(KEYINPUT56), .ZN(n1010) );
  XNOR2_X1 U1078 ( .A(G1956), .B(G299), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(G303), .A2(G1971), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n1000) );
  XNOR2_X1 U1083 ( .A(n1011), .B(n992), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G301), .B(n993), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G1348), .B(n996), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G168), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(n1003), .B(KEYINPUT57), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(KEYINPUT124), .B(n1004), .Z(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1038) );
  INV_X1 U1096 ( .A(G16), .ZN(n1036) );
  XNOR2_X1 U1097 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n1034) );
  XNOR2_X1 U1098 ( .A(G1961), .B(G5), .ZN(n1024) );
  XNOR2_X1 U1099 ( .A(G19), .B(n1011), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(G1956), .B(G20), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G6), .B(G1981), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT59), .B(G1348), .Z(n1016) );
  XNOR2_X1 U1105 ( .A(G4), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT60), .B(n1019), .Z(n1021) );
  XNOR2_X1 U1108 ( .A(G1966), .B(G21), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(KEYINPUT125), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(KEYINPUT126), .B(n1025), .ZN(n1032) );
  XOR2_X1 U1113 ( .A(G1986), .B(G24), .Z(n1027) );
  XOR2_X1 U1114 ( .A(G1971), .B(G22), .Z(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(G23), .B(G1976), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1118 ( .A(KEYINPUT58), .B(n1030), .ZN(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1120 ( .A(n1034), .B(n1033), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1122 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1123 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NAND2_X1 U1124 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1043), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

