//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G137), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT65), .B1(new_n196), .B2(G134), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(new_n198), .C1(new_n194), .C2(G137), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(G131), .B1(new_n199), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n194), .B2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n201), .A4(new_n195), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT64), .A2(G143), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT64), .A2(G143), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n211), .B1(new_n214), .B2(G146), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n209), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n215), .A2(new_n216), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n224));
  INV_X1    g038(.A(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT2), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G113), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n224), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n233));
  INV_X1    g047(.A(G116), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G119), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT68), .A3(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(G119), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT67), .A4(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n226), .A2(new_n228), .A3(new_n224), .ZN(new_n243));
  OAI22_X1  g057(.A1(new_n241), .A2(new_n242), .B1(new_n243), .B2(new_n229), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n208), .A2(new_n223), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  OR2_X1    g059(.A1(KEYINPUT64), .A2(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT64), .A2(G143), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(G146), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n248), .A2(new_n210), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT1), .B1(new_n252), .B2(G146), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n217), .A2(new_n219), .B1(G128), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT70), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n195), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n194), .A2(G137), .ZN(new_n257));
  OAI21_X1  g071(.A(G131), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n207), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n248), .A2(new_n210), .A3(new_n250), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT64), .B(G143), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n218), .B1(new_n262), .B2(new_n209), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n249), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n260), .B(new_n261), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n255), .A2(new_n259), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n245), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT72), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n208), .A2(new_n223), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n207), .A3(new_n258), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n244), .A2(new_n240), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n245), .A2(new_n266), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n268), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT28), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n267), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n193), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n277), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n276), .B1(new_n245), .B2(new_n266), .ZN(new_n284));
  INV_X1    g098(.A(new_n193), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT66), .B1(new_n272), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n289));
  AOI211_X1 g103(.A(new_n289), .B(KEYINPUT30), .C1(new_n269), .C2(new_n271), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n208), .B2(new_n223), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n291), .A2(new_n266), .A3(KEYINPUT71), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT71), .B1(new_n291), .B2(new_n266), .ZN(new_n293));
  OAI22_X1  g107(.A1(new_n288), .A2(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n286), .B1(new_n294), .B2(new_n273), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n291), .A2(new_n266), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n291), .A2(new_n266), .A3(KEYINPUT71), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n223), .A2(new_n208), .B1(new_n259), .B2(new_n270), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n289), .B1(new_n303), .B2(KEYINPUT30), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n272), .A2(KEYINPUT66), .A3(new_n287), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n306), .A3(new_n274), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT31), .A3(new_n286), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n282), .B1(new_n297), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G472), .A2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n187), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT32), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n279), .A2(new_n281), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n285), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n307), .A2(KEYINPUT31), .A3(new_n286), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT31), .B1(new_n307), .B2(new_n286), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT73), .A3(new_n310), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n312), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n312), .A2(new_n319), .A3(KEYINPUT74), .A4(new_n313), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n283), .A2(new_n284), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n266), .A2(new_n269), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n273), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT28), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n281), .B(KEYINPUT77), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n285), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G902), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n307), .A2(new_n325), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT76), .B1(new_n335), .B2(new_n285), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n337), .B(new_n193), .C1(new_n307), .C2(new_n325), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n281), .A2(new_n193), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(new_n278), .B2(KEYINPUT28), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n330), .B1(new_n341), .B2(new_n342), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n334), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G472), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT78), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n268), .A2(new_n277), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n300), .A2(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(new_n274), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n337), .B1(new_n352), .B2(new_n193), .ZN(new_n353));
  INV_X1    g167(.A(new_n340), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n279), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT29), .B1(new_n355), .B2(KEYINPUT75), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n335), .A2(KEYINPUT76), .A3(new_n285), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n353), .A2(new_n356), .A3(new_n357), .A4(new_n343), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n332), .A2(new_n333), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n348), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n309), .A2(new_n311), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n360), .A2(new_n361), .B1(new_n362), .B2(KEYINPUT32), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n324), .A2(new_n349), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n189), .A2(G227), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n365), .B(new_n366), .Z(new_n367));
  AND2_X1   g181(.A1(new_n255), .A2(new_n265), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n369));
  INV_X1    g183(.A(G101), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G104), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G107), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n371), .A3(G104), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n377), .A2(new_n374), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(new_n373), .B2(G107), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n370), .A4(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n377), .A3(new_n374), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT85), .B1(new_n382), .B2(G101), .ZN(new_n383));
  AOI211_X1 g197(.A(new_n369), .B(new_n375), .C1(new_n381), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n383), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT84), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n388), .A3(G101), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n385), .A2(KEYINPUT4), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n215), .A2(new_n216), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n220), .A2(new_n222), .ZN(new_n392));
  XOR2_X1   g206(.A(KEYINPUT86), .B(KEYINPUT4), .Z(new_n393));
  NAND3_X1  g207(.A1(new_n382), .A2(G101), .A3(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n368), .A2(new_n384), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n208), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT88), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n375), .B1(new_n381), .B2(new_n383), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n249), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n260), .B1(new_n400), .B2(new_n215), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XOR2_X1   g216(.A(KEYINPUT87), .B(KEYINPUT10), .Z(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n398), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AOI211_X1 g219(.A(KEYINPUT88), .B(new_n403), .C1(new_n399), .C2(new_n401), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n396), .B(new_n397), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT89), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n399), .A2(new_n401), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT88), .B1(new_n409), .B2(new_n403), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n402), .A2(new_n398), .A3(new_n404), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT89), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n397), .A4(new_n396), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n367), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT90), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n399), .A2(new_n270), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n416), .B(new_n208), .C1(new_n409), .C2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT91), .A3(KEYINPUT12), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n420));
  INV_X1    g234(.A(new_n399), .ZN(new_n421));
  INV_X1    g235(.A(new_n270), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n397), .B1(new_n423), .B2(new_n402), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n420), .B1(new_n424), .B2(new_n416), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n208), .B1(new_n409), .B2(new_n417), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(KEYINPUT91), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n419), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n415), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n367), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n408), .A2(new_n414), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n387), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n381), .A2(new_n383), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n395), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n399), .A2(new_n255), .A3(KEYINPUT10), .A4(new_n265), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n410), .B2(new_n411), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n439), .A2(new_n397), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n432), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n431), .B1(new_n441), .B2(KEYINPUT93), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT93), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n415), .A2(new_n430), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(new_n333), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n432), .B1(new_n430), .B2(new_n433), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n439), .A2(new_n397), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n415), .B2(KEYINPUT92), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n433), .A2(new_n432), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n448), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G469), .B1(new_n454), .B2(G902), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n447), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G214), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(G952), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n458), .A2(KEYINPUT101), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(KEYINPUT101), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n189), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(G234), .B2(G237), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(G898), .ZN(new_n463));
  AOI211_X1 g277(.A(new_n333), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G125), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n223), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n422), .A2(new_n467), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G224), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G953), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n470), .B(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n244), .A2(new_n240), .A3(new_n394), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n390), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n239), .A2(new_n231), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(KEYINPUT94), .A2(KEYINPUT5), .ZN(new_n478));
  NOR2_X1   g292(.A1(KEYINPUT94), .A2(KEYINPUT5), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n480), .A2(new_n235), .A3(new_n237), .A4(new_n238), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT95), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n478), .A2(new_n479), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n234), .A2(G119), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n225), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n481), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n482), .B1(new_n481), .B2(new_n485), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n399), .B(new_n477), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n475), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n490));
  XNOR2_X1  g304(.A(G110), .B(G122), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT97), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT97), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n489), .A2(new_n495), .A3(new_n490), .A4(new_n492), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n489), .A2(new_n492), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n475), .A2(new_n491), .A3(new_n488), .ZN(new_n499));
  AND4_X1   g313(.A1(KEYINPUT96), .A2(new_n498), .A3(KEYINPUT6), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n490), .B1(new_n489), .B2(new_n492), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT96), .B1(new_n501), .B2(new_n499), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n473), .B(new_n497), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n472), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT7), .A4(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n505), .A2(KEYINPUT99), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(KEYINPUT99), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n468), .A2(new_n469), .B1(KEYINPUT7), .B2(new_n504), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n499), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n486), .A2(new_n487), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n421), .B1(new_n511), .B2(new_n476), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n241), .A2(KEYINPUT98), .A3(KEYINPUT5), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT98), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n239), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n513), .A2(new_n485), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n399), .A2(new_n517), .A3(new_n477), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n491), .B(KEYINPUT8), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n510), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n509), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G210), .B1(G237), .B2(G902), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n503), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n523), .B1(new_n503), .B2(new_n522), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n457), .B(new_n466), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT81), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT82), .B1(new_n528), .B2(G125), .ZN(new_n529));
  NAND2_X1  g343(.A1(KEYINPUT82), .A2(G125), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(G140), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT82), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n467), .B2(KEYINPUT81), .ZN(new_n534));
  INV_X1    g348(.A(G140), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n527), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT16), .B1(new_n535), .B2(G125), .ZN(new_n538));
  OAI21_X1  g352(.A(G146), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n538), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n535), .B1(new_n534), .B2(new_n530), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n529), .A2(G140), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n209), .B(new_n540), .C1(new_n543), .C2(new_n527), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n188), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n545));
  INV_X1    g359(.A(G214), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n546), .A2(G237), .A3(G953), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n262), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(KEYINPUT17), .A3(G131), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(G131), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n214), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n206), .A3(new_n545), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n539), .A2(new_n544), .A3(new_n549), .A4(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n548), .A2(new_n557), .A3(new_n206), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n552), .A2(new_n545), .B1(KEYINPUT18), .B2(G131), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n535), .A2(G125), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n467), .A2(G140), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G146), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n209), .B1(new_n532), .B2(new_n536), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n558), .A2(new_n559), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G113), .B(G122), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(new_n373), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n556), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n556), .B2(new_n565), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n333), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G475), .ZN(new_n572));
  INV_X1    g386(.A(new_n562), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT19), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n575), .B(new_n209), .C1(new_n543), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n550), .A2(new_n553), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n539), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n579), .A2(new_n565), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n568), .B1(new_n580), .B2(new_n567), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT20), .ZN(new_n582));
  NOR2_X1   g396(.A1(G475), .A2(G902), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n582), .B1(new_n581), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n572), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n214), .A2(G128), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n249), .A2(G143), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n194), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(G116), .B(G122), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n371), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n589), .A2(KEYINPUT13), .A3(new_n590), .ZN(new_n594));
  OAI21_X1  g408(.A(G134), .B1(new_n589), .B2(KEYINPUT13), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n591), .B(new_n593), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G122), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G116), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n371), .B1(new_n598), .B2(KEYINPUT14), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n592), .ZN(new_n600));
  INV_X1    g414(.A(new_n591), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n194), .B1(new_n589), .B2(new_n590), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT9), .B(G234), .ZN(new_n605));
  INV_X1    g419(.A(G217), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n605), .A2(new_n606), .A3(G953), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n596), .A2(new_n603), .A3(new_n607), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G478), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(KEYINPUT15), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n611), .B(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n588), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n526), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(G221), .B1(new_n605), .B2(G902), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n456), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n539), .A2(new_n544), .ZN(new_n621));
  INV_X1    g435(.A(G110), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT23), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n236), .B2(G128), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n249), .A2(KEYINPUT23), .A3(G119), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n624), .B(new_n625), .C1(G119), .C2(new_n249), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT80), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n627), .B2(new_n626), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT24), .B(G110), .Z(new_n630));
  XNOR2_X1  g444(.A(G119), .B(G128), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT79), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n621), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT83), .B(G110), .ZN(new_n635));
  OAI22_X1  g449(.A1(new_n626), .A2(new_n635), .B1(new_n631), .B2(new_n630), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n539), .B(new_n636), .C1(G146), .C2(new_n562), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT22), .B(G137), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n634), .A2(new_n637), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(G902), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT25), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n606), .B1(G234), .B2(new_n333), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n645), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n648), .A2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n364), .A2(new_n620), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G101), .ZN(G3));
  AOI211_X1 g470(.A(G469), .B(G902), .C1(new_n442), .C2(new_n444), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n430), .A2(new_n433), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n367), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n440), .B1(new_n451), .B2(new_n452), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n415), .A2(KEYINPUT92), .ZN(new_n661));
  OAI211_X1 g475(.A(G469), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(G469), .A2(G902), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n619), .B1(new_n657), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n309), .B2(G902), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n312), .A2(new_n666), .A3(new_n319), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n665), .A2(new_n653), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n457), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n503), .A2(new_n522), .ZN(new_n670));
  INV_X1    g484(.A(new_n523), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n503), .A2(new_n522), .A3(new_n523), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n611), .A2(new_n612), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n612), .A2(new_n333), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n609), .A2(new_n610), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT33), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT33), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n609), .A2(new_n680), .A3(new_n610), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n675), .B(new_n677), .C1(new_n682), .C2(new_n612), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n588), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n674), .A2(new_n466), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n668), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT34), .B(G104), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G6));
  INV_X1    g503(.A(new_n586), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n584), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n556), .A2(new_n565), .ZN(new_n692));
  INV_X1    g506(.A(new_n567), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(G902), .B1(new_n694), .B2(new_n568), .ZN(new_n695));
  INV_X1    g509(.A(G475), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT102), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n571), .A2(new_n698), .A3(G475), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n691), .A2(new_n700), .A3(new_n466), .A4(new_n615), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(KEYINPUT103), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(KEYINPUT103), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n674), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n668), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT35), .B(G107), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G9));
  INV_X1    g522(.A(new_n619), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n447), .B2(new_n455), .ZN(new_n710));
  INV_X1    g524(.A(new_n667), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n642), .A2(KEYINPUT36), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n638), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n651), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n649), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n710), .A2(new_n618), .A3(new_n711), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT104), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT37), .B(G110), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G12));
  INV_X1    g533(.A(new_n462), .ZN(new_n720));
  INV_X1    g534(.A(new_n464), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n720), .B1(G900), .B2(new_n721), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n691), .A2(new_n700), .A3(new_n615), .A4(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n723), .B(new_n457), .C1(new_n524), .C2(new_n525), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT105), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n672), .A2(new_n673), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n457), .A4(new_n723), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n729), .A2(new_n710), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n364), .A3(new_n715), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G128), .ZN(G30));
  NAND2_X1  g546(.A1(new_n362), .A2(KEYINPUT32), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n352), .A2(new_n285), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n333), .B1(new_n327), .B2(new_n193), .ZN(new_n735));
  OAI21_X1  g549(.A(G472), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n324), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n715), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n722), .B(KEYINPUT39), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n710), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n742), .A2(KEYINPUT40), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(KEYINPUT40), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n726), .B(KEYINPUT38), .Z(new_n745));
  AND3_X1   g559(.A1(new_n587), .A2(new_n457), .A3(new_n615), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n740), .A2(new_n743), .A3(new_n744), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n262), .ZN(G45));
  NAND2_X1  g564(.A1(new_n675), .A2(new_n677), .ZN(new_n751));
  INV_X1    g565(.A(new_n682), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(G478), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(new_n587), .A3(new_n722), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n754), .B(new_n457), .C1(new_n524), .C2(new_n525), .ZN(new_n755));
  AOI211_X1 g569(.A(new_n709), .B(new_n755), .C1(new_n447), .C2(new_n455), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n364), .A2(new_n715), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G146), .ZN(G48));
  AND3_X1   g572(.A1(new_n415), .A2(new_n430), .A3(new_n443), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n449), .B1(new_n414), .B2(new_n408), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n443), .B1(new_n760), .B2(new_n432), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n759), .B1(new_n431), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(G469), .B1(new_n762), .B2(G902), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n619), .A3(new_n447), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n364), .A2(new_n654), .A3(new_n686), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT41), .B(G113), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT106), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n766), .B(new_n768), .ZN(G15));
  NOR2_X1   g583(.A1(new_n764), .A2(new_n704), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n364), .A2(new_n770), .A3(new_n654), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G116), .ZN(G18));
  AND4_X1   g586(.A1(new_n674), .A2(new_n763), .A3(new_n619), .A4(new_n447), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n617), .A2(new_n465), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n364), .A2(new_n715), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G119), .ZN(G21));
  NOR2_X1   g590(.A1(new_n316), .A2(new_n317), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n193), .B1(new_n328), .B2(new_n329), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n310), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n666), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n653), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n747), .B1(new_n672), .B2(new_n673), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n765), .A2(new_n466), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G122), .ZN(G24));
  INV_X1    g598(.A(new_n780), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n715), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n753), .A2(new_n587), .A3(new_n722), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT107), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n773), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G125), .ZN(G27));
  INV_X1    g605(.A(KEYINPUT42), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT108), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n672), .A2(new_n794), .A3(new_n457), .A4(new_n673), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT108), .B1(new_n726), .B2(new_n669), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n710), .A2(new_n793), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n358), .A2(new_n359), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n361), .A3(G472), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n313), .B1(new_n309), .B2(new_n311), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n349), .A2(new_n733), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n654), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n796), .A2(new_n795), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n665), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n788), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n364), .A2(new_n805), .A3(new_n654), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n808));
  AOI21_X1  g622(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n206), .ZN(G33));
  NAND4_X1  g624(.A1(new_n364), .A2(new_n805), .A3(new_n654), .A4(new_n723), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G134), .ZN(G36));
  AND2_X1   g626(.A1(new_n454), .A2(KEYINPUT45), .ZN(new_n813));
  OAI21_X1  g627(.A(G469), .B1(new_n454), .B2(KEYINPUT45), .ZN(new_n814));
  OAI221_X1 g628(.A(new_n663), .B1(new_n813), .B2(new_n814), .C1(KEYINPUT46), .C2(new_n657), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(KEYINPUT110), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n709), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n813), .A2(new_n814), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(new_n663), .ZN(new_n819));
  OAI211_X1 g633(.A(KEYINPUT110), .B(new_n815), .C1(new_n819), .C2(KEYINPUT46), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n804), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT111), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n587), .A2(new_n683), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT43), .Z(new_n826));
  INV_X1    g640(.A(new_n715), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n711), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(KEYINPUT44), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n823), .A2(KEYINPUT111), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n826), .A2(new_n827), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(KEYINPUT44), .A3(new_n667), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n824), .A2(new_n829), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n822), .A2(new_n741), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G137), .ZN(G39));
  NOR4_X1   g649(.A1(new_n364), .A2(new_n654), .A3(new_n787), .A4(new_n804), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n838), .A2(KEYINPUT47), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(KEYINPUT47), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n821), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n817), .A2(new_n820), .A3(new_n838), .A4(KEYINPUT47), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(new_n535), .ZN(G42));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n826), .A2(new_n720), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n781), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n830), .A2(new_n824), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n841), .A2(new_n842), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n763), .A2(new_n447), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(new_n709), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n764), .A2(new_n804), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n846), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT115), .Z(new_n856));
  INV_X1    g670(.A(new_n786), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n739), .A2(new_n654), .A3(new_n854), .A4(new_n462), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n588), .A2(new_n683), .ZN(new_n860));
  OR3_X1    g674(.A1(new_n859), .A2(KEYINPUT116), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n848), .A2(new_n669), .A3(new_n745), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n862), .A2(KEYINPUT50), .A3(new_n764), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT116), .B1(new_n859), .B2(new_n860), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT50), .B1(new_n862), .B2(new_n764), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n861), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n845), .B1(new_n853), .B2(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT51), .Z(new_n869));
  INV_X1    g683(.A(new_n802), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n856), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT48), .Z(new_n872));
  AOI21_X1  g686(.A(new_n461), .B1(new_n848), .B2(new_n773), .ZN(new_n873));
  INV_X1    g687(.A(new_n684), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n873), .B1(new_n859), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n722), .B(new_n746), .C1(new_n524), .C2(new_n525), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n709), .B(new_n878), .C1(new_n447), .C2(new_n455), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n738), .A2(new_n879), .A3(new_n827), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n731), .A2(new_n757), .A3(new_n790), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n349), .A2(new_n733), .A3(new_n799), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n827), .B1(new_n884), .B2(new_n324), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n730), .B2(new_n756), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(KEYINPUT52), .A3(new_n790), .A4(new_n880), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT113), .B1(new_n526), .B2(new_n874), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n674), .A2(new_n891), .A3(new_n466), .A4(new_n684), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n674), .A2(new_n466), .A3(new_n588), .A4(new_n615), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(new_n654), .A3(new_n710), .A4(new_n711), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n775), .A2(new_n655), .A3(new_n783), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n766), .A2(new_n771), .A3(new_n716), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n805), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n691), .A2(new_n700), .A3(new_n616), .A4(new_n722), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n322), .A2(new_n323), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n363), .A2(new_n349), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n715), .B(new_n900), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n789), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n811), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n809), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n898), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n877), .B1(new_n889), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT54), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n809), .A2(new_n906), .A3(new_n905), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n888), .A2(new_n912), .A3(KEYINPUT53), .A4(new_n898), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n913), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT54), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n876), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  OAI22_X1  g731(.A1(new_n869), .A2(new_n917), .B1(G952), .B2(G953), .ZN(new_n918));
  AND4_X1   g732(.A1(new_n654), .A2(new_n457), .A3(new_n619), .A4(new_n825), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n739), .A2(new_n745), .A3(new_n919), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n851), .B(KEYINPUT49), .Z(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G75));
  AOI21_X1  g736(.A(new_n333), .B1(new_n910), .B2(new_n913), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n923), .A2(G210), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n924), .A2(KEYINPUT56), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n497), .B1(new_n500), .B2(new_n502), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n473), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT55), .Z(new_n928));
  AND2_X1   g742(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n458), .A2(G953), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT117), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n925), .B2(new_n928), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n929), .A2(new_n932), .ZN(G51));
  INV_X1    g747(.A(new_n931), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n663), .B(KEYINPUT57), .Z(new_n935));
  INV_X1    g749(.A(KEYINPUT118), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n916), .B2(new_n914), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n936), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n935), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n445), .ZN(new_n942));
  INV_X1    g756(.A(new_n818), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n923), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT119), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n934), .B1(new_n942), .B2(new_n945), .ZN(G54));
  NAND3_X1  g760(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(new_n581), .Z(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(new_n934), .ZN(G60));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n676), .B(KEYINPUT59), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n752), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n914), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n911), .B1(new_n910), .B2(new_n913), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT118), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n956), .B2(new_n939), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n951), .B1(new_n916), .B2(new_n914), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n931), .B1(new_n958), .B2(new_n682), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n950), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n951), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n954), .B2(new_n955), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n934), .B1(new_n962), .B2(new_n752), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n952), .B1(new_n937), .B2(new_n940), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT120), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n960), .A2(new_n965), .ZN(G63));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT60), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n789), .B1(new_n885), .B2(new_n900), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n811), .B1(new_n970), .B2(new_n899), .ZN(new_n971));
  NOR4_X1   g785(.A1(new_n971), .A2(new_n809), .A3(new_n896), .A4(new_n897), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT53), .B1(new_n972), .B2(new_n888), .ZN(new_n973));
  AND4_X1   g787(.A1(KEYINPUT53), .A2(new_n888), .A3(new_n912), .A4(new_n898), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n934), .B1(new_n975), .B2(new_n645), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT121), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT61), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n968), .B1(new_n910), .B2(new_n913), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n931), .B1(new_n979), .B2(new_n650), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n915), .A2(new_n713), .A3(new_n969), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT122), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT122), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n979), .A2(new_n713), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n976), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n978), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n977), .B(new_n931), .C1(new_n979), .C2(new_n650), .ZN(new_n988));
  AOI22_X1  g802(.A1(new_n982), .A2(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n986), .A2(new_n989), .ZN(G66));
  XOR2_X1   g804(.A(new_n898), .B(KEYINPUT123), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n189), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(G953), .B1(new_n463), .B2(new_n471), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n926), .B1(G898), .B2(new_n189), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G69));
  AND2_X1   g812(.A1(new_n886), .A2(new_n790), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n749), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n843), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n874), .B1(new_n587), .B2(new_n616), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n364), .A2(new_n654), .A3(new_n823), .A4(new_n1004), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n1005), .A2(new_n742), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1002), .A2(new_n1003), .A3(new_n834), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n189), .ZN(new_n1008));
  INV_X1    g822(.A(new_n543), .ZN(new_n1009));
  AOI22_X1  g823(.A1(new_n1009), .A2(KEYINPUT19), .B1(new_n573), .B2(new_n574), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n294), .B(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(KEYINPUT125), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n870), .A2(new_n782), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n822), .A2(new_n741), .A3(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n999), .A2(new_n811), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n834), .A2(new_n1015), .A3(new_n1016), .A4(new_n908), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n189), .B1(new_n1017), .B2(new_n843), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n189), .A2(G900), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1018), .A2(KEYINPUT126), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1011), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(KEYINPUT126), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1012), .B(new_n1013), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT126), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1028), .A2(new_n1021), .A3(new_n1020), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1013), .B1(new_n1029), .B2(new_n1012), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1025), .A2(new_n1030), .ZN(G72));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT63), .Z(new_n1033));
  XNOR2_X1  g847(.A(new_n1033), .B(KEYINPUT127), .ZN(new_n1034));
  OR2_X1    g848(.A1(new_n1017), .A2(new_n843), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1034), .B1(new_n1035), .B2(new_n991), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1036), .A2(new_n285), .A3(new_n352), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1034), .B1(new_n1007), .B2(new_n991), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n734), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n339), .A2(new_n295), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n915), .A2(new_n1033), .A3(new_n1040), .ZN(new_n1041));
  AND4_X1   g855(.A1(new_n931), .A2(new_n1037), .A3(new_n1039), .A4(new_n1041), .ZN(G57));
endmodule


