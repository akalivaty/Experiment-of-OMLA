//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(G8gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G8gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  XOR2_X1   g014(.A(KEYINPUT97), .B(G36gat), .Z(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(KEYINPUT15), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n213), .B(new_n211), .C1(new_n216), .C2(new_n215), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(new_n217), .A3(new_n218), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n226), .B1(new_n219), .B2(new_n223), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n209), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n223), .A2(new_n219), .B1(new_n206), .B2(new_n207), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n224), .B(new_n208), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT98), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n229), .B(KEYINPUT13), .Z(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n224), .A2(new_n208), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n239), .B2(new_n230), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT98), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n229), .A4(new_n231), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n234), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT96), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT11), .B(G169gat), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n234), .A2(new_n242), .A3(new_n243), .A4(new_n250), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(G71gat), .A2(G78gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G71gat), .A2(G78gat), .ZN(new_n257));
  AND2_X1   g056(.A1(G57gat), .A2(G64gat), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n256), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n261));
  INV_X1    g060(.A(G64gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n257), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(KEYINPUT9), .B2(new_n255), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n260), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G127gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n209), .B1(new_n267), .B2(new_n266), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(G155gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G183gat), .B(G211gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n273), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G190gat), .B(G218gat), .Z(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G85gat), .A2(G92gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT7), .ZN(new_n283));
  NAND2_X1  g082(.A1(G99gat), .A2(G106gat), .ZN(new_n284));
  INV_X1    g083(.A(G85gat), .ZN(new_n285));
  INV_X1    g084(.A(G92gat), .ZN(new_n286));
  AOI22_X1  g085(.A1(KEYINPUT8), .A2(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G99gat), .B(G106gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT101), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n283), .A2(new_n289), .A3(new_n287), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n292), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n289), .B1(new_n283), .B2(new_n287), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n225), .B2(new_n227), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n294), .ZN(new_n300));
  NAND2_X1  g099(.A1(G232gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n224), .A2(new_n300), .B1(KEYINPUT41), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n281), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n299), .A2(new_n281), .A3(new_n303), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n302), .A2(KEYINPUT41), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT100), .ZN(new_n308));
  XNOR2_X1  g107(.A(G134gat), .B(G162gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT102), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n305), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n305), .A2(new_n306), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT102), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n279), .A2(new_n318), .A3(KEYINPUT103), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT103), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n278), .B2(new_n317), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n297), .A2(new_n294), .A3(new_n266), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n266), .A2(new_n296), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT104), .A3(new_n293), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT104), .B1(new_n323), .B2(new_n293), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G230gat), .A2(G233gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g129(.A1(new_n330), .A2(KEYINPUT106), .ZN(new_n331));
  XNOR2_X1  g130(.A(G120gat), .B(G148gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G176gat), .B(G204gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(KEYINPUT106), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT10), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n337), .B(new_n322), .C1(new_n325), .C2(new_n326), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n266), .A2(new_n337), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n300), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n329), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT105), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n341), .A2(KEYINPUT105), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n336), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n341), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n334), .B1(new_n346), .B2(new_n330), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n319), .A2(new_n321), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  OR2_X1    g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(G197gat), .A2(G204gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G211gat), .A2(G218gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT22), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G211gat), .ZN(new_n358));
  INV_X1    g157(.A(G218gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n360), .A2(new_n361), .A3(new_n354), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n360), .B2(new_n354), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n357), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n354), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT78), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n351), .A2(new_n352), .B1(new_n355), .B2(new_n354), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n360), .A2(new_n361), .A3(new_n354), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n364), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT2), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(KEYINPUT83), .A3(KEYINPUT2), .ZN(new_n378));
  INV_X1    g177(.A(G141gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G148gat), .ZN(new_n380));
  INV_X1    g179(.A(G148gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G141gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n377), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n374), .A2(KEYINPUT81), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(G155gat), .A3(G162gat), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n385), .A2(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n381), .A3(G141gat), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT84), .B1(new_n379), .B2(G148gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n379), .A2(G148gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n374), .A2(new_n399), .A3(KEYINPUT2), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n375), .A2(KEYINPUT85), .ZN(new_n401));
  XNOR2_X1  g200(.A(G155gat), .B(G162gat), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n398), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n393), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n373), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT88), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n373), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n357), .A2(new_n362), .A3(new_n363), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n364), .A2(new_n369), .A3(KEYINPUT79), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n393), .A2(new_n403), .A3(new_n372), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n370), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n406), .A2(new_n408), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G22gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n419), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n404), .A2(KEYINPUT86), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n393), .A2(new_n403), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n373), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n417), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n420), .A2(new_n421), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT89), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT31), .B(G50gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n405), .A2(KEYINPUT88), .B1(new_n414), .B2(new_n416), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n422), .B1(new_n434), .B2(new_n408), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n417), .A2(new_n422), .A3(new_n426), .ZN(new_n436));
  OAI21_X1  g235(.A(G22gat), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n430), .A2(new_n433), .B1(new_n428), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n437), .A2(new_n428), .A3(KEYINPUT89), .A4(new_n433), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n423), .A2(KEYINPUT3), .A3(new_n425), .ZN(new_n442));
  NOR2_X1   g241(.A1(G127gat), .A2(G134gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT71), .B(G127gat), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(G134gat), .ZN(new_n445));
  INV_X1    g244(.A(G113gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(G120gat), .ZN(new_n447));
  INV_X1    g246(.A(G120gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G113gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n449), .A3(KEYINPUT72), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT1), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT72), .B1(new_n447), .B2(new_n449), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n445), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT73), .B(G120gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n447), .B1(new_n455), .B2(new_n446), .ZN(new_n456));
  INV_X1    g255(.A(new_n443), .ZN(new_n457));
  NAND2_X1  g256(.A1(G127gat), .A2(G134gat), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT1), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n461), .A2(new_n415), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT4), .B1(new_n461), .B2(new_n404), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT72), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n448), .A2(G113gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n446), .A2(G120gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(new_n451), .A3(new_n450), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n469), .A2(new_n445), .B1(new_n456), .B2(new_n459), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n401), .A2(new_n400), .A3(new_n402), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n471), .A2(new_n398), .B1(new_n384), .B2(new_n392), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT4), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n464), .A2(new_n474), .A3(KEYINPUT87), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n470), .A2(new_n472), .A3(new_n476), .A4(new_n473), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n463), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n423), .A2(new_n461), .A3(new_n425), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n470), .A2(new_n472), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n479), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT39), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G1gat), .B(G29gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT0), .ZN(new_n489));
  XNOR2_X1  g288(.A(G57gat), .B(G85gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT91), .B(KEYINPUT39), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n480), .A3(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n487), .A2(KEYINPUT40), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT4), .B(new_n479), .C1(new_n461), .C2(new_n404), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n442), .A2(new_n462), .B1(new_n496), .B2(new_n474), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT5), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n480), .A2(KEYINPUT5), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n463), .A2(new_n475), .A3(new_n477), .A4(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n491), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT40), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n494), .A2(new_n492), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n485), .B1(new_n480), .B2(new_n478), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT92), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT92), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G169gat), .A2(G176gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(G169gat), .A2(G176gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT26), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT70), .ZN(new_n518));
  INV_X1    g317(.A(G169gat), .ZN(new_n519));
  INV_X1    g318(.A(G176gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n518), .B1(new_n521), .B2(KEYINPUT26), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n515), .A2(KEYINPUT70), .A3(new_n516), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n514), .B(new_n517), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT69), .ZN(new_n526));
  XOR2_X1   g325(.A(KEYINPUT27), .B(G183gat), .Z(new_n527));
  OR2_X1    g326(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n526), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G183gat), .A2(G190gat), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n528), .A2(new_n529), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G183gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n524), .A2(new_n531), .A3(new_n532), .A4(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT23), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT23), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT67), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n541), .A3(new_n514), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT66), .B(G176gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n540), .A2(G169gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n542), .A2(new_n521), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(G183gat), .A2(G190gat), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT65), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT65), .ZN(new_n552));
  AND3_X1   g351(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT64), .ZN(new_n554));
  NAND3_X1  g353(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT64), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n549), .A2(new_n552), .A3(new_n554), .A4(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT25), .B1(new_n545), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n553), .A2(new_n547), .ZN(new_n560));
  INV_X1    g359(.A(G183gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n528), .A2(new_n561), .A3(new_n529), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n542), .A2(new_n521), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n544), .B2(new_n520), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n537), .B1(new_n559), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(G226gat), .A2(G233gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n414), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n568), .A2(new_n370), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n569), .ZN(new_n573));
  XNOR2_X1  g372(.A(G8gat), .B(G36gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(G64gat), .B(G92gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  AOI21_X1  g375(.A(new_n569), .B1(new_n568), .B2(new_n370), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT80), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n570), .B1(new_n572), .B2(new_n569), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n578), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n573), .B(new_n576), .C1(new_n581), .C2(new_n571), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT30), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n570), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n578), .B1(new_n585), .B2(new_n577), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT80), .B1(new_n572), .B2(new_n569), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n571), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n573), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(KEYINPUT30), .A3(new_n576), .ZN(new_n591));
  INV_X1    g390(.A(new_n576), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n588), .B2(new_n589), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n584), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n441), .B1(new_n513), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n496), .A2(new_n474), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n463), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n482), .A2(new_n483), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n597), .B(KEYINPUT5), .C1(new_n479), .C2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT6), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n502), .A4(new_n491), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n492), .A2(KEYINPUT6), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n491), .A2(new_n600), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n602), .B(new_n603), .C1(new_n500), .C2(new_n503), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n582), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n576), .A2(KEYINPUT38), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n573), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n606), .B1(new_n588), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n414), .B1(new_n586), .B2(new_n587), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT37), .B1(new_n580), .B2(new_n571), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT93), .B1(new_n605), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n604), .A2(new_n601), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n585), .A2(new_n577), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n607), .B1(new_n616), .B2(new_n414), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n581), .B2(new_n414), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT37), .B1(new_n616), .B2(new_n571), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n581), .B2(new_n571), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n620), .A3(new_n606), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT93), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n615), .A2(new_n621), .A3(new_n622), .A4(new_n582), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n590), .A2(new_n607), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n592), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT38), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n614), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n595), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n595), .B2(new_n627), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n568), .A2(new_n470), .ZN(new_n631));
  NAND2_X1  g430(.A1(G227gat), .A2(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n461), .B(new_n537), .C1(new_n559), .C2(new_n567), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n636));
  XNOR2_X1  g435(.A(G15gat), .B(G43gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G71gat), .B(G99gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n635), .B(KEYINPUT32), .C1(new_n636), .C2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n639), .B1(new_n635), .B2(KEYINPUT32), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT74), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n635), .A2(new_n636), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n641), .B2(new_n643), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT77), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n633), .B1(new_n631), .B2(new_n634), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT76), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT34), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n649), .B1(new_n648), .B2(new_n651), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n646), .A2(new_n647), .A3(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n658), .B(new_n640), .C1(new_n645), .C2(new_n644), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n647), .B1(new_n646), .B2(new_n656), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT36), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT90), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n438), .B2(new_n440), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n437), .A2(new_n428), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n436), .B1(new_n419), .B2(new_n418), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT89), .B1(new_n666), .B2(new_n421), .ZN(new_n667));
  INV_X1    g466(.A(new_n433), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(KEYINPUT90), .A3(new_n439), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n604), .A2(new_n601), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n584), .A2(new_n591), .A3(new_n671), .A4(new_n593), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n664), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n646), .A2(new_n656), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT36), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n662), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n629), .A2(new_n630), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n661), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n669), .A2(new_n439), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n657), .A4(new_n659), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT35), .B1(new_n681), .B2(new_n672), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n659), .A2(new_n674), .ZN(new_n683));
  INV_X1    g482(.A(new_n672), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n680), .A4(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n254), .B(new_n350), .C1(new_n678), .C2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n682), .A2(new_n686), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n595), .A2(new_n627), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT94), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n595), .A2(new_n627), .A3(new_n628), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n691), .B1(new_n695), .B2(new_n677), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n696), .A2(KEYINPUT107), .A3(new_n254), .A4(new_n350), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n615), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G1gat), .ZN(G1324gat));
  INV_X1    g499(.A(G8gat), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n698), .B2(new_n594), .ZN(new_n702));
  INV_X1    g501(.A(new_n594), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT16), .B(G8gat), .ZN(new_n704));
  AOI211_X1 g503(.A(new_n703), .B(new_n704), .C1(new_n690), .C2(new_n697), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n698), .A2(new_n594), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n709), .B2(new_n704), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n706), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n707), .B1(new_n706), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(G1325gat));
  INV_X1    g512(.A(new_n698), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n662), .A2(new_n676), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G15gat), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(G15gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n698), .A2(new_n718), .A3(new_n683), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1326gat));
  NAND2_X1  g519(.A1(new_n664), .A2(new_n670), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n698), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(KEYINPUT109), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(KEYINPUT109), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT43), .B(G22gat), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n725), .B2(new_n726), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(G1327gat));
  AND2_X1   g529(.A1(new_n696), .A2(new_n317), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT44), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n696), .A2(new_n317), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n233), .A2(new_n232), .B1(new_n238), .B2(new_n241), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n250), .B1(new_n738), .B2(new_n243), .ZN(new_n739));
  INV_X1    g538(.A(new_n253), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n252), .A2(KEYINPUT110), .A3(new_n253), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n348), .A2(new_n278), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n736), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G29gat), .B1(new_n746), .B2(new_n671), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n696), .A2(new_n254), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n744), .A2(new_n318), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n748), .A2(G29gat), .A3(new_n671), .A4(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT45), .Z(new_n752));
  NAND2_X1  g551(.A1(new_n747), .A2(new_n752), .ZN(G1328gat));
  INV_X1    g552(.A(new_n216), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n746), .B2(new_n703), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n748), .A2(new_n754), .A3(new_n703), .A4(new_n750), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(G1329gat));
  NOR2_X1   g557(.A1(new_n750), .A2(G43gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n683), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n748), .A2(new_n760), .B1(new_n761), .B2(KEYINPUT47), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n732), .A2(new_n715), .A3(new_n735), .A4(new_n745), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(G43gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(KEYINPUT47), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n764), .B(new_n765), .Z(G1330gat));
  INV_X1    g565(.A(G50gat), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n736), .A2(new_n745), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(new_n441), .ZN(new_n769));
  NOR4_X1   g568(.A1(new_n748), .A2(G50gat), .A3(new_n721), .A4(new_n750), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n736), .A2(new_n722), .A3(new_n745), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n770), .B1(new_n773), .B2(G50gat), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n769), .A2(new_n772), .B1(new_n774), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g574(.A(new_n348), .ZN(new_n776));
  AND4_X1   g575(.A1(new_n321), .A2(new_n319), .A3(new_n776), .A4(new_n743), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n696), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n615), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n594), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT49), .B(G64gat), .Z(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(G1333gat));
  INV_X1    g583(.A(G71gat), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n778), .B2(new_n715), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n683), .A2(new_n785), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g588(.A1(new_n778), .A2(new_n722), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G78gat), .ZN(G1335gat));
  INV_X1    g590(.A(new_n743), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n279), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n731), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT51), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n731), .A2(new_n796), .A3(new_n793), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n795), .A2(new_n776), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n285), .A3(new_n615), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n792), .A2(new_n279), .A3(new_n348), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n736), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n615), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n802), .B2(new_n285), .ZN(G1336gat));
  NOR2_X1   g602(.A1(new_n703), .A2(G92gat), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n795), .A2(new_n776), .A3(new_n797), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n732), .A2(new_n594), .A3(new_n735), .A4(new_n800), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G92gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(KEYINPUT112), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT52), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n805), .B(new_n807), .C1(KEYINPUT112), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1337gat));
  AOI21_X1  g612(.A(G99gat), .B1(new_n798), .B2(new_n683), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n715), .A2(G99gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n801), .B2(new_n815), .ZN(G1338gat));
  NOR2_X1   g615(.A1(new_n680), .A2(G106gat), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n795), .A2(new_n776), .A3(new_n797), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n732), .A2(new_n441), .A3(new_n735), .A4(new_n800), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G106gat), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n732), .A2(new_n722), .A3(new_n735), .A4(new_n800), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n798), .A2(new_n817), .B1(G106gat), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n824), .B2(new_n821), .ZN(G1339gat));
  INV_X1    g624(.A(KEYINPUT105), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n346), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n338), .A2(new_n340), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n830), .B2(new_n329), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(new_n831), .A3(new_n342), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n334), .B1(new_n341), .B2(new_n828), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n345), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n836), .A2(new_n741), .A3(new_n742), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n229), .B1(new_n228), .B2(new_n231), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n235), .A2(new_n237), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n249), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n253), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n347), .B2(new_n345), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n317), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n834), .A2(new_n835), .ZN(new_n845));
  INV_X1    g644(.A(new_n345), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n846), .A3(new_n837), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n842), .A2(new_n317), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n278), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n350), .A2(new_n743), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n722), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n683), .A2(new_n615), .A3(new_n703), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT113), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(KEYINPUT113), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n254), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n857), .A2(new_n446), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n671), .B1(new_n850), .B2(new_n851), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n681), .A2(new_n594), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(G113gat), .B1(new_n863), .B2(new_n792), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n859), .A2(new_n864), .ZN(G1340gat));
  OAI21_X1  g664(.A(G120gat), .B1(new_n857), .B2(new_n348), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n348), .A2(new_n455), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n862), .B2(new_n867), .ZN(G1341gat));
  NAND4_X1  g667(.A1(new_n855), .A2(new_n444), .A3(new_n279), .A4(new_n856), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n444), .B1(new_n863), .B2(new_n279), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G1342gat));
  OAI21_X1  g672(.A(G134gat), .B1(new_n857), .B2(new_n318), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n318), .A2(G134gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n862), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n874), .A2(new_n880), .ZN(G1343gat));
  NOR3_X1   g680(.A1(new_n715), .A2(new_n594), .A3(new_n680), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n860), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(G141gat), .A3(new_n858), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n680), .B1(new_n850), .B2(new_n851), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n715), .A2(new_n671), .A3(new_n594), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n845), .A2(new_n254), .A3(new_n846), .A4(new_n837), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n317), .B1(new_n889), .B2(new_n843), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n890), .A2(new_n891), .B1(new_n847), .B2(new_n848), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n278), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n721), .B1(new_n894), .B2(new_n851), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n887), .B(new_n888), .C1(new_n895), .C2(new_n886), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n792), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n884), .B1(new_n898), .B2(G141gat), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n379), .B1(new_n897), .B2(new_n254), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n884), .A2(KEYINPUT58), .ZN(new_n902));
  OAI22_X1  g701(.A1(new_n899), .A2(new_n900), .B1(new_n901), .B2(new_n902), .ZN(G1344gat));
  NAND4_X1  g702(.A1(new_n860), .A2(new_n381), .A3(new_n776), .A4(new_n882), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n776), .ZN(new_n906));
  AOI211_X1 g705(.A(new_n886), .B(new_n680), .C1(new_n850), .C2(new_n851), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n278), .B1(new_n890), .B2(new_n849), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n254), .B2(new_n349), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n722), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT117), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n885), .A2(KEYINPUT57), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n906), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n381), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n906), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n909), .A2(new_n722), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n886), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n913), .B1(new_n920), .B2(new_n912), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n907), .A2(KEYINPUT117), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT118), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n905), .B1(new_n917), .B2(new_n924), .ZN(new_n925));
  AOI211_X1 g724(.A(KEYINPUT59), .B(new_n381), .C1(new_n897), .C2(new_n776), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n904), .B1(new_n925), .B2(new_n926), .ZN(G1345gat));
  OAI21_X1  g726(.A(G155gat), .B1(new_n896), .B2(new_n278), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n278), .A2(G155gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n883), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT119), .ZN(G1346gat));
  NOR3_X1   g730(.A1(new_n883), .A2(G162gat), .A3(new_n318), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT120), .ZN(new_n933));
  OAI21_X1  g732(.A(G162gat), .B1(new_n896), .B2(new_n318), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT121), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1347gat));
  AOI21_X1  g738(.A(new_n615), .B1(new_n850), .B2(new_n851), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n681), .A2(new_n703), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n519), .A3(new_n792), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n683), .A2(new_n671), .A3(new_n594), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT122), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n852), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G169gat), .B1(new_n947), .B2(new_n858), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n944), .B1(new_n950), .B2(new_n951), .ZN(G1348gat));
  OR3_X1    g751(.A1(new_n947), .A2(new_n543), .A3(new_n348), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  AOI21_X1  g755(.A(G176gat), .B1(new_n943), .B2(new_n776), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(G1349gat));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n527), .A3(new_n278), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT125), .ZN(new_n960));
  OAI21_X1  g759(.A(G183gat), .B1(new_n947), .B2(new_n278), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT60), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT60), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n960), .A2(new_n964), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n943), .A2(new_n533), .A3(new_n317), .ZN(new_n967));
  OAI21_X1  g766(.A(G190gat), .B1(new_n947), .B2(new_n318), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  NAND3_X1  g770(.A1(new_n716), .A2(new_n594), .A3(new_n441), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n940), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(G197gat), .B1(new_n976), .B2(new_n792), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n911), .A2(new_n914), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n715), .A2(new_n615), .A3(new_n703), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n254), .A2(G197gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(G1352gat));
  OAI21_X1  g782(.A(G204gat), .B1(new_n980), .B2(new_n348), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n975), .A2(G204gat), .A3(new_n348), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(G1353gat));
  NAND3_X1  g786(.A1(new_n978), .A2(new_n279), .A3(new_n979), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(G211gat), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT63), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT63), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n988), .A2(new_n991), .A3(G211gat), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n358), .A3(new_n279), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  OAI211_X1 g795(.A(new_n990), .B(new_n992), .C1(new_n995), .C2(new_n996), .ZN(G1354gat));
  OAI21_X1  g796(.A(G218gat), .B1(new_n980), .B2(new_n318), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n976), .A2(new_n359), .A3(new_n317), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1355gat));
endmodule


