

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U551 ( .A(KEYINPUT66), .B(n537), .ZN(n586) );
  INV_X1 U552 ( .A(KEYINPUT30), .ZN(n720) );
  INV_X1 U553 ( .A(n733), .ZN(n711) );
  INV_X1 U554 ( .A(KEYINPUT102), .ZN(n724) );
  INV_X1 U555 ( .A(KEYINPUT100), .ZN(n717) );
  NAND2_X1 U556 ( .A1(n680), .A2(n776), .ZN(n733) );
  NAND2_X1 U557 ( .A1(G8), .A2(n733), .ZN(n806) );
  XNOR2_X1 U558 ( .A(KEYINPUT70), .B(KEYINPUT12), .ZN(n556) );
  NOR2_X1 U559 ( .A1(G1384), .A2(G164), .ZN(n679) );
  XNOR2_X1 U560 ( .A(n557), .B(n556), .ZN(n559) );
  OR2_X1 U561 ( .A1(n678), .A2(n677), .ZN(n775) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n633) );
  NOR2_X1 U563 ( .A1(G651), .A2(n619), .ZN(n634) );
  INV_X1 U564 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U565 ( .A1(n522), .A2(G2104), .ZN(n518) );
  XNOR2_X2 U566 ( .A(n518), .B(KEYINPUT65), .ZN(n1004) );
  NAND2_X1 U567 ( .A1(n1004), .A2(G102), .ZN(n521) );
  AND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n999) );
  NAND2_X1 U569 ( .A1(G114), .A2(n999), .ZN(n519) );
  XOR2_X1 U570 ( .A(KEYINPUT85), .B(n519), .Z(n520) );
  NAND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U572 ( .A1(G2104), .A2(n522), .ZN(n1000) );
  NAND2_X1 U573 ( .A1(G126), .A2(n1000), .ZN(n525) );
  NOR2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n523), .Z(n1003) );
  NAND2_X1 U576 ( .A1(G138), .A2(n1003), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n527), .A2(n526), .ZN(G164) );
  NAND2_X1 U579 ( .A1(G101), .A2(n1004), .ZN(n528) );
  XOR2_X1 U580 ( .A(KEYINPUT23), .B(n528), .Z(n674) );
  NAND2_X1 U581 ( .A1(n1003), .A2(G137), .ZN(n673) );
  NAND2_X1 U582 ( .A1(G113), .A2(n999), .ZN(n530) );
  NAND2_X1 U583 ( .A1(G125), .A2(n1000), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n675) );
  INV_X1 U585 ( .A(n675), .ZN(n531) );
  AND2_X1 U586 ( .A1(n673), .A2(n531), .ZN(n532) );
  AND2_X1 U587 ( .A1(n674), .A2(n532), .ZN(G160) );
  NAND2_X1 U588 ( .A1(G85), .A2(n633), .ZN(n534) );
  XOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .Z(n619) );
  INV_X1 U590 ( .A(G651), .ZN(n535) );
  NOR2_X1 U591 ( .A1(n619), .A2(n535), .ZN(n637) );
  NAND2_X1 U592 ( .A1(G72), .A2(n637), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G47), .A2(n634), .ZN(n539) );
  NOR2_X1 U595 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n536), .Z(n537) );
  NAND2_X1 U597 ( .A1(G60), .A2(n586), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U599 ( .A1(n541), .A2(n540), .ZN(G290) );
  XNOR2_X1 U600 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U602 ( .A(G108), .ZN(G238) );
  NAND2_X1 U603 ( .A1(n637), .A2(G76), .ZN(n542) );
  XNOR2_X1 U604 ( .A(KEYINPUT72), .B(n542), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n633), .A2(G89), .ZN(n543) );
  XNOR2_X1 U606 ( .A(KEYINPUT4), .B(n543), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U608 ( .A(n546), .B(KEYINPUT5), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n634), .A2(G51), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT73), .B(n547), .Z(n549) );
  NAND2_X1 U611 ( .A1(G63), .A2(n586), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(n550), .Z(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U615 ( .A(n553), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U619 ( .A(G223), .B(KEYINPUT69), .ZN(n832) );
  NAND2_X1 U620 ( .A1(n832), .A2(G567), .ZN(n555) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(n555), .Z(G234) );
  NAND2_X1 U622 ( .A1(G81), .A2(n633), .ZN(n557) );
  NAND2_X1 U623 ( .A1(G68), .A2(n637), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(KEYINPUT13), .ZN(n562) );
  NAND2_X1 U626 ( .A1(G43), .A2(n634), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n586), .A2(G56), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(n563), .Z(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X2 U631 ( .A(KEYINPUT71), .B(n566), .Z(n923) );
  NAND2_X1 U632 ( .A1(n923), .A2(G860), .ZN(G153) );
  NAND2_X1 U633 ( .A1(G52), .A2(n634), .ZN(n568) );
  NAND2_X1 U634 ( .A1(G64), .A2(n586), .ZN(n567) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G90), .A2(n633), .ZN(n570) );
  NAND2_X1 U637 ( .A1(G77), .A2(n637), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U639 ( .A(KEYINPUT9), .B(n571), .Z(n572) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT67), .B(n574), .ZN(G301) );
  NAND2_X1 U642 ( .A1(G868), .A2(G301), .ZN(n583) );
  NAND2_X1 U643 ( .A1(G92), .A2(n633), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G79), .A2(n637), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G54), .A2(n634), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G66), .A2(n586), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U650 ( .A(KEYINPUT15), .B(n581), .ZN(n1023) );
  INV_X1 U651 ( .A(G868), .ZN(n653) );
  NAND2_X1 U652 ( .A1(n1023), .A2(n653), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U654 ( .A1(G91), .A2(n633), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G78), .A2(n637), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n586), .A2(G65), .ZN(n587) );
  XOR2_X1 U658 ( .A(KEYINPUT68), .B(n587), .Z(n588) );
  NOR2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n634), .A2(G53), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(G299) );
  NOR2_X1 U662 ( .A1(G286), .A2(n653), .ZN(n593) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n592) );
  NOR2_X1 U664 ( .A1(n593), .A2(n592), .ZN(G297) );
  INV_X1 U665 ( .A(G559), .ZN(n596) );
  NOR2_X1 U666 ( .A1(G860), .A2(n596), .ZN(n594) );
  NOR2_X1 U667 ( .A1(n1023), .A2(n594), .ZN(n595) );
  XOR2_X1 U668 ( .A(KEYINPUT16), .B(n595), .Z(G148) );
  INV_X1 U669 ( .A(n1023), .ZN(n687) );
  NAND2_X1 U670 ( .A1(n596), .A2(n687), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n597), .A2(G868), .ZN(n599) );
  INV_X1 U672 ( .A(n923), .ZN(n683) );
  NAND2_X1 U673 ( .A1(n683), .A2(n653), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U675 ( .A1(G111), .A2(n999), .ZN(n601) );
  NAND2_X1 U676 ( .A1(G99), .A2(n1004), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U678 ( .A(KEYINPUT74), .B(n602), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n1000), .A2(G123), .ZN(n603) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(n603), .Z(n604) );
  NOR2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n1003), .A2(G135), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U684 ( .A(KEYINPUT75), .B(n608), .ZN(n1018) );
  XNOR2_X1 U685 ( .A(n1018), .B(G2096), .ZN(n609) );
  INV_X1 U686 ( .A(G2100), .ZN(n970) );
  NAND2_X1 U687 ( .A1(n609), .A2(n970), .ZN(G156) );
  NAND2_X1 U688 ( .A1(n687), .A2(G559), .ZN(n651) );
  XOR2_X1 U689 ( .A(n923), .B(n651), .Z(n610) );
  NOR2_X1 U690 ( .A1(G860), .A2(n610), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G93), .A2(n633), .ZN(n612) );
  NAND2_X1 U692 ( .A1(G80), .A2(n637), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G55), .A2(n634), .ZN(n614) );
  NAND2_X1 U695 ( .A1(G67), .A2(n586), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n615) );
  OR2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n654) );
  XOR2_X1 U698 ( .A(n654), .B(KEYINPUT76), .Z(n617) );
  XNOR2_X1 U699 ( .A(n618), .B(n617), .ZN(G145) );
  NAND2_X1 U700 ( .A1(G87), .A2(n619), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G74), .A2(G651), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n586), .A2(n622), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n634), .A2(G49), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U706 ( .A1(G50), .A2(n634), .ZN(n625) );
  XOR2_X1 U707 ( .A(KEYINPUT78), .B(n625), .Z(n630) );
  NAND2_X1 U708 ( .A1(G88), .A2(n633), .ZN(n627) );
  NAND2_X1 U709 ( .A1(G75), .A2(n637), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U711 ( .A(KEYINPUT79), .B(n628), .Z(n629) );
  NOR2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G62), .A2(n586), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(G303) );
  INV_X1 U715 ( .A(G303), .ZN(G166) );
  NAND2_X1 U716 ( .A1(G61), .A2(n586), .ZN(n642) );
  NAND2_X1 U717 ( .A1(G86), .A2(n633), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G48), .A2(n634), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n637), .A2(G73), .ZN(n638) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n638), .Z(n639) );
  NOR2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U724 ( .A(KEYINPUT77), .B(n643), .Z(G305) );
  XOR2_X1 U725 ( .A(KEYINPUT80), .B(KEYINPUT19), .Z(n644) );
  XNOR2_X1 U726 ( .A(G288), .B(n644), .ZN(n645) );
  XOR2_X1 U727 ( .A(G299), .B(n645), .Z(n648) );
  XOR2_X1 U728 ( .A(n654), .B(G290), .Z(n646) );
  XOR2_X1 U729 ( .A(n646), .B(G166), .Z(n647) );
  XNOR2_X1 U730 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U731 ( .A(n649), .B(n923), .Z(n650) );
  XNOR2_X1 U732 ( .A(n650), .B(G305), .ZN(n1022) );
  XNOR2_X1 U733 ( .A(n1022), .B(n651), .ZN(n652) );
  NOR2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n656) );
  NOR2_X1 U735 ( .A1(G868), .A2(n654), .ZN(n655) );
  NOR2_X1 U736 ( .A1(n656), .A2(n655), .ZN(G295) );
  XOR2_X1 U737 ( .A(KEYINPUT81), .B(KEYINPUT21), .Z(n660) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n657) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U740 ( .A1(n658), .A2(G2090), .ZN(n659) );
  XNOR2_X1 U741 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U742 ( .A1(G2072), .A2(n661), .ZN(G158) );
  NAND2_X1 U743 ( .A1(G120), .A2(G69), .ZN(n662) );
  NOR2_X1 U744 ( .A1(G238), .A2(n662), .ZN(n663) );
  NAND2_X1 U745 ( .A1(G57), .A2(n663), .ZN(n957) );
  NAND2_X1 U746 ( .A1(G567), .A2(n957), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n664), .B(KEYINPUT83), .ZN(n670) );
  XOR2_X1 U748 ( .A(KEYINPUT82), .B(KEYINPUT22), .Z(n666) );
  NAND2_X1 U749 ( .A1(G132), .A2(G82), .ZN(n665) );
  XNOR2_X1 U750 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n667), .A2(G96), .ZN(n668) );
  OR2_X1 U752 ( .A1(G218), .A2(n668), .ZN(n958) );
  AND2_X1 U753 ( .A1(G2106), .A2(n958), .ZN(n669) );
  NOR2_X1 U754 ( .A1(n670), .A2(n669), .ZN(G319) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n671) );
  INV_X1 U756 ( .A(G319), .ZN(n1027) );
  NOR2_X1 U757 ( .A1(n671), .A2(n1027), .ZN(n672) );
  XNOR2_X1 U758 ( .A(n672), .B(KEYINPUT84), .ZN(n835) );
  NAND2_X1 U759 ( .A1(G36), .A2(n835), .ZN(G176) );
  XNOR2_X1 U760 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n831) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n678) );
  INV_X1 U762 ( .A(G40), .ZN(n676) );
  OR2_X1 U763 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U764 ( .A(KEYINPUT93), .B(n775), .ZN(n680) );
  XNOR2_X1 U765 ( .A(n679), .B(KEYINPUT64), .ZN(n776) );
  AND2_X1 U766 ( .A1(n711), .A2(G1996), .ZN(n681) );
  XOR2_X1 U767 ( .A(n681), .B(KEYINPUT26), .Z(n685) );
  AND2_X1 U768 ( .A1(n733), .A2(G1341), .ZN(n682) );
  NOR2_X1 U769 ( .A1(n683), .A2(n682), .ZN(n684) );
  AND2_X1 U770 ( .A1(n685), .A2(n684), .ZN(n688) );
  NOR2_X1 U771 ( .A1(n687), .A2(n688), .ZN(n686) );
  XNOR2_X1 U772 ( .A(KEYINPUT99), .B(n686), .ZN(n695) );
  NAND2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n692) );
  NOR2_X1 U774 ( .A1(G2067), .A2(n733), .ZN(n690) );
  NOR2_X1 U775 ( .A1(n711), .A2(G1348), .ZN(n689) );
  NOR2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U777 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U778 ( .A(n693), .B(KEYINPUT98), .ZN(n694) );
  NAND2_X1 U779 ( .A1(n695), .A2(n694), .ZN(n704) );
  INV_X1 U780 ( .A(G299), .ZN(n706) );
  INV_X1 U781 ( .A(KEYINPUT97), .ZN(n702) );
  XOR2_X1 U782 ( .A(KEYINPUT95), .B(KEYINPUT27), .Z(n697) );
  NAND2_X1 U783 ( .A1(G2072), .A2(n711), .ZN(n696) );
  XNOR2_X1 U784 ( .A(n697), .B(n696), .ZN(n700) );
  NAND2_X1 U785 ( .A1(G1956), .A2(n733), .ZN(n698) );
  XOR2_X1 U786 ( .A(KEYINPUT96), .B(n698), .Z(n699) );
  NOR2_X1 U787 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U788 ( .A(n702), .B(n701), .ZN(n705) );
  NAND2_X1 U789 ( .A1(n706), .A2(n705), .ZN(n703) );
  NAND2_X1 U790 ( .A1(n704), .A2(n703), .ZN(n709) );
  NOR2_X1 U791 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U792 ( .A(n707), .B(KEYINPUT28), .Z(n708) );
  NAND2_X1 U793 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U794 ( .A(n710), .B(KEYINPUT29), .ZN(n716) );
  NAND2_X1 U795 ( .A1(G1961), .A2(n733), .ZN(n713) );
  XOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .Z(n846) );
  NAND2_X1 U797 ( .A1(n711), .A2(n846), .ZN(n712) );
  NAND2_X1 U798 ( .A1(n713), .A2(n712), .ZN(n726) );
  NOR2_X1 U799 ( .A1(G301), .A2(n726), .ZN(n714) );
  XNOR2_X1 U800 ( .A(n714), .B(KEYINPUT94), .ZN(n715) );
  NOR2_X1 U801 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U802 ( .A(n718), .B(n717), .ZN(n731) );
  NOR2_X1 U803 ( .A1(G1966), .A2(n806), .ZN(n745) );
  NOR2_X1 U804 ( .A1(G2084), .A2(n733), .ZN(n742) );
  NOR2_X1 U805 ( .A1(n745), .A2(n742), .ZN(n719) );
  AND2_X1 U806 ( .A1(n719), .A2(G8), .ZN(n721) );
  XNOR2_X1 U807 ( .A(n721), .B(n720), .ZN(n722) );
  XOR2_X1 U808 ( .A(KEYINPUT101), .B(n722), .Z(n723) );
  NOR2_X1 U809 ( .A1(G168), .A2(n723), .ZN(n725) );
  XNOR2_X1 U810 ( .A(n725), .B(n724), .ZN(n728) );
  NAND2_X1 U811 ( .A1(G301), .A2(n726), .ZN(n727) );
  NAND2_X1 U812 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U813 ( .A(KEYINPUT31), .B(n729), .ZN(n730) );
  NAND2_X1 U814 ( .A1(n731), .A2(n730), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n743), .A2(G286), .ZN(n740) );
  INV_X1 U816 ( .A(G8), .ZN(n738) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n806), .ZN(n732) );
  XNOR2_X1 U818 ( .A(KEYINPUT103), .B(n732), .ZN(n736) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U820 ( .A1(G166), .A2(n734), .ZN(n735) );
  NAND2_X1 U821 ( .A1(n736), .A2(n735), .ZN(n737) );
  OR2_X1 U822 ( .A1(n738), .A2(n737), .ZN(n739) );
  AND2_X1 U823 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U824 ( .A(n741), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U825 ( .A1(G8), .A2(n742), .ZN(n747) );
  INV_X1 U826 ( .A(n743), .ZN(n744) );
  NOR2_X1 U827 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U828 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U829 ( .A1(n749), .A2(n748), .ZN(n805) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n934) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n931) );
  NOR2_X1 U832 ( .A1(n934), .A2(n931), .ZN(n751) );
  INV_X1 U833 ( .A(KEYINPUT33), .ZN(n750) );
  AND2_X1 U834 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U835 ( .A1(n805), .A2(n752), .ZN(n797) );
  INV_X1 U836 ( .A(n806), .ZN(n753) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n935) );
  AND2_X1 U838 ( .A1(n753), .A2(n935), .ZN(n754) );
  NOR2_X1 U839 ( .A1(KEYINPUT33), .A2(n754), .ZN(n757) );
  NAND2_X1 U840 ( .A1(n934), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n755), .A2(n806), .ZN(n756) );
  NOR2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n781) );
  XOR2_X1 U843 ( .A(G1981), .B(G305), .Z(n927) );
  NAND2_X1 U844 ( .A1(G131), .A2(n1003), .ZN(n759) );
  NAND2_X1 U845 ( .A1(G95), .A2(n1004), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U847 ( .A(KEYINPUT90), .B(n760), .ZN(n764) );
  NAND2_X1 U848 ( .A1(G107), .A2(n999), .ZN(n762) );
  NAND2_X1 U849 ( .A1(G119), .A2(n1000), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n1010) );
  INV_X1 U852 ( .A(G1991), .ZN(n984) );
  NOR2_X1 U853 ( .A1(n1010), .A2(n984), .ZN(n774) );
  NAND2_X1 U854 ( .A1(G117), .A2(n999), .ZN(n766) );
  NAND2_X1 U855 ( .A1(G129), .A2(n1000), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n770) );
  NAND2_X1 U857 ( .A1(G105), .A2(n1004), .ZN(n767) );
  XNOR2_X1 U858 ( .A(n767), .B(KEYINPUT38), .ZN(n768) );
  XNOR2_X1 U859 ( .A(n768), .B(KEYINPUT91), .ZN(n769) );
  NOR2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n1003), .A2(G141), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n1014) );
  AND2_X1 U863 ( .A1(G1996), .A2(n1014), .ZN(n773) );
  NOR2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n884) );
  NOR2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n777), .B(KEYINPUT86), .ZN(n826) );
  XOR2_X1 U867 ( .A(KEYINPUT92), .B(n826), .Z(n778) );
  NOR2_X1 U868 ( .A1(n884), .A2(n778), .ZN(n819) );
  INV_X1 U869 ( .A(n819), .ZN(n779) );
  AND2_X1 U870 ( .A1(n927), .A2(n779), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n795) );
  NAND2_X1 U872 ( .A1(n1004), .A2(G104), .ZN(n782) );
  XOR2_X1 U873 ( .A(KEYINPUT87), .B(n782), .Z(n784) );
  NAND2_X1 U874 ( .A1(n1003), .A2(G140), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n785), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G116), .A2(n999), .ZN(n787) );
  NAND2_X1 U878 ( .A1(G128), .A2(n1000), .ZN(n786) );
  NAND2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U880 ( .A(n788), .B(KEYINPUT35), .Z(n789) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U882 ( .A(KEYINPUT36), .B(n791), .Z(n792) );
  XOR2_X1 U883 ( .A(KEYINPUT88), .B(n792), .Z(n1017) );
  XNOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  OR2_X1 U885 ( .A1(n1017), .A2(n824), .ZN(n793) );
  XNOR2_X1 U886 ( .A(n793), .B(KEYINPUT89), .ZN(n892) );
  NAND2_X1 U887 ( .A1(n892), .A2(n826), .ZN(n822) );
  INV_X1 U888 ( .A(n822), .ZN(n794) );
  OR2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n813) );
  NOR2_X1 U891 ( .A1(G2090), .A2(G303), .ZN(n798) );
  NAND2_X1 U892 ( .A1(G8), .A2(n798), .ZN(n799) );
  XNOR2_X1 U893 ( .A(n799), .B(KEYINPUT104), .ZN(n803) );
  NOR2_X1 U894 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XOR2_X1 U895 ( .A(n800), .B(KEYINPUT24), .Z(n801) );
  NOR2_X1 U896 ( .A1(n806), .A2(n801), .ZN(n807) );
  INV_X1 U897 ( .A(n807), .ZN(n802) );
  AND2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n804) );
  AND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n811) );
  NOR2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U901 ( .A1(n819), .A2(n808), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n822), .A2(n809), .ZN(n810) );
  NOR2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U905 ( .A(n814), .B(KEYINPUT105), .ZN(n816) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n930) );
  NAND2_X1 U907 ( .A1(n930), .A2(n826), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n829) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n1014), .ZN(n877) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n817) );
  AND2_X1 U911 ( .A1(n984), .A2(n1010), .ZN(n885) );
  NOR2_X1 U912 ( .A1(n817), .A2(n885), .ZN(n818) );
  NOR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U914 ( .A1(n877), .A2(n820), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n1017), .A2(n824), .ZN(n889) );
  NAND2_X1 U918 ( .A1(n825), .A2(n889), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U921 ( .A(n831), .B(n830), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U924 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G120), .B(KEYINPUT109), .ZN(G236) );
  XOR2_X1 U928 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  NAND2_X1 U930 ( .A1(G124), .A2(n1000), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n836), .B(KEYINPUT44), .ZN(n838) );
  NAND2_X1 U932 ( .A1(n999), .A2(G112), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n838), .A2(n837), .ZN(n842) );
  NAND2_X1 U934 ( .A1(G136), .A2(n1003), .ZN(n840) );
  NAND2_X1 U935 ( .A1(G100), .A2(n1004), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n841) );
  NOR2_X1 U937 ( .A1(n842), .A2(n841), .ZN(G162) );
  XNOR2_X1 U938 ( .A(G2090), .B(G35), .ZN(n855) );
  XOR2_X1 U939 ( .A(G25), .B(G1991), .Z(n843) );
  NAND2_X1 U940 ( .A1(n843), .A2(G28), .ZN(n852) );
  XNOR2_X1 U941 ( .A(G2067), .B(G26), .ZN(n845) );
  XNOR2_X1 U942 ( .A(G33), .B(G2072), .ZN(n844) );
  NOR2_X1 U943 ( .A1(n845), .A2(n844), .ZN(n850) );
  XNOR2_X1 U944 ( .A(G1996), .B(G32), .ZN(n848) );
  XNOR2_X1 U945 ( .A(G27), .B(n846), .ZN(n847) );
  NOR2_X1 U946 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U947 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U948 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U949 ( .A(KEYINPUT53), .B(n853), .ZN(n854) );
  NOR2_X1 U950 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U951 ( .A(KEYINPUT120), .B(n856), .ZN(n860) );
  XNOR2_X1 U952 ( .A(KEYINPUT54), .B(G34), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n857), .B(KEYINPUT121), .ZN(n858) );
  XNOR2_X1 U954 ( .A(G2084), .B(n858), .ZN(n859) );
  NAND2_X1 U955 ( .A1(n860), .A2(n859), .ZN(n863) );
  NOR2_X1 U956 ( .A1(G29), .A2(KEYINPUT55), .ZN(n861) );
  NAND2_X1 U957 ( .A1(n863), .A2(n861), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G11), .A2(n862), .ZN(n900) );
  INV_X1 U959 ( .A(KEYINPUT55), .ZN(n894) );
  OR2_X1 U960 ( .A1(n894), .A2(n863), .ZN(n898) );
  XNOR2_X1 U961 ( .A(G164), .B(G2078), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n864), .B(KEYINPUT119), .ZN(n874) );
  NAND2_X1 U963 ( .A1(G139), .A2(n1003), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G103), .A2(n1004), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U966 ( .A1(G115), .A2(n999), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G127), .A2(n1000), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U969 ( .A(KEYINPUT115), .B(n869), .ZN(n870) );
  XNOR2_X1 U970 ( .A(KEYINPUT47), .B(n870), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n996) );
  XOR2_X1 U972 ( .A(G2072), .B(n996), .Z(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(KEYINPUT50), .B(n875), .ZN(n880) );
  XOR2_X1 U975 ( .A(G2090), .B(G162), .Z(n876) );
  NOR2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U977 ( .A(KEYINPUT51), .B(n878), .Z(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n882) );
  XOR2_X1 U979 ( .A(G160), .B(G2084), .Z(n881) );
  NOR2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n888) );
  NOR2_X1 U982 ( .A1(n885), .A2(n1018), .ZN(n886) );
  XOR2_X1 U983 ( .A(KEYINPUT118), .B(n886), .Z(n887) );
  NOR2_X1 U984 ( .A1(n888), .A2(n887), .ZN(n890) );
  NAND2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n891) );
  NOR2_X1 U986 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U987 ( .A(n893), .B(KEYINPUT52), .ZN(n895) );
  NAND2_X1 U988 ( .A1(n895), .A2(n894), .ZN(n896) );
  NAND2_X1 U989 ( .A1(G29), .A2(n896), .ZN(n897) );
  NAND2_X1 U990 ( .A1(n898), .A2(n897), .ZN(n899) );
  NOR2_X1 U991 ( .A1(n900), .A2(n899), .ZN(n955) );
  XNOR2_X1 U992 ( .A(G1348), .B(KEYINPUT59), .ZN(n901) );
  XNOR2_X1 U993 ( .A(n901), .B(G4), .ZN(n905) );
  XNOR2_X1 U994 ( .A(G1341), .B(G19), .ZN(n903) );
  XNOR2_X1 U995 ( .A(G1956), .B(G20), .ZN(n902) );
  NOR2_X1 U996 ( .A1(n903), .A2(n902), .ZN(n904) );
  NAND2_X1 U997 ( .A1(n905), .A2(n904), .ZN(n908) );
  XOR2_X1 U998 ( .A(G6), .B(G1981), .Z(n906) );
  XNOR2_X1 U999 ( .A(KEYINPUT125), .B(n906), .ZN(n907) );
  NOR2_X1 U1000 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(KEYINPUT60), .B(n909), .ZN(n913) );
  XNOR2_X1 U1002 ( .A(G1966), .B(G21), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(G5), .B(G1961), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1005 ( .A1(n913), .A2(n912), .ZN(n920) );
  XNOR2_X1 U1006 ( .A(G1971), .B(G22), .ZN(n915) );
  XNOR2_X1 U1007 ( .A(G23), .B(G1976), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(n915), .A2(n914), .ZN(n917) );
  XOR2_X1 U1009 ( .A(G1986), .B(G24), .Z(n916) );
  NAND2_X1 U1010 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1011 ( .A(KEYINPUT58), .B(n918), .ZN(n919) );
  NOR2_X1 U1012 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1013 ( .A(KEYINPUT61), .B(n921), .Z(n922) );
  NOR2_X1 U1014 ( .A1(G16), .A2(n922), .ZN(n952) );
  XOR2_X1 U1015 ( .A(KEYINPUT56), .B(G16), .Z(n950) );
  XNOR2_X1 U1016 ( .A(n923), .B(G1341), .ZN(n925) );
  XOR2_X1 U1017 ( .A(G301), .B(G1961), .Z(n924) );
  NAND2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n947) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G168), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(n926), .B(KEYINPUT122), .ZN(n928) );
  NAND2_X1 U1021 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1022 ( .A(n929), .B(KEYINPUT57), .ZN(n945) );
  NOR2_X1 U1023 ( .A1(n931), .A2(n930), .ZN(n941) );
  XOR2_X1 U1024 ( .A(G299), .B(G1956), .Z(n933) );
  NAND2_X1 U1025 ( .A1(G1971), .A2(G303), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n939) );
  INV_X1 U1027 ( .A(n934), .ZN(n936) );
  NAND2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1029 ( .A(KEYINPUT123), .B(n937), .Z(n938) );
  NOR2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1031 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1032 ( .A(n1023), .B(G1348), .ZN(n942) );
  NOR2_X1 U1033 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1034 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1035 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1036 ( .A(KEYINPUT124), .B(n948), .ZN(n949) );
  NOR2_X1 U1037 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1038 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(n953), .B(KEYINPUT126), .ZN(n954) );
  NAND2_X1 U1040 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1041 ( .A(KEYINPUT62), .B(n956), .Z(G311) );
  XNOR2_X1 U1042 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1043 ( .A(G132), .ZN(G219) );
  INV_X1 U1044 ( .A(G96), .ZN(G221) );
  INV_X1 U1045 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1046 ( .A1(n958), .A2(n957), .ZN(G325) );
  INV_X1 U1047 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1048 ( .A(G2443), .B(G2430), .Z(n960) );
  XNOR2_X1 U1049 ( .A(G1348), .B(G2451), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(n960), .B(n959), .ZN(n967) );
  XOR2_X1 U1051 ( .A(G2438), .B(KEYINPUT107), .Z(n962) );
  XNOR2_X1 U1052 ( .A(G1341), .B(G2454), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(n962), .B(n961), .ZN(n963) );
  XOR2_X1 U1054 ( .A(n963), .B(G2435), .Z(n965) );
  XNOR2_X1 U1055 ( .A(G2446), .B(G2427), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(n965), .B(n964), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n967), .B(n966), .ZN(n968) );
  NAND2_X1 U1058 ( .A1(n968), .A2(G14), .ZN(n969) );
  XOR2_X1 U1059 ( .A(KEYINPUT108), .B(n969), .Z(G401) );
  XNOR2_X1 U1060 ( .A(KEYINPUT42), .B(n970), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(G2067), .B(G2084), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n972), .B(n971), .ZN(n973) );
  XOR2_X1 U1063 ( .A(n973), .B(G2678), .Z(n975) );
  XNOR2_X1 U1064 ( .A(G2090), .B(KEYINPUT111), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n975), .B(n974), .ZN(n979) );
  XOR2_X1 U1066 ( .A(G2096), .B(KEYINPUT43), .Z(n977) );
  XNOR2_X1 U1067 ( .A(G2072), .B(G2078), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n977), .B(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(n979), .B(n978), .Z(G227) );
  XOR2_X1 U1070 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n981) );
  XNOR2_X1 U1071 ( .A(G1981), .B(G1976), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n981), .B(n980), .ZN(n992) );
  XOR2_X1 U1073 ( .A(KEYINPUT41), .B(G2474), .Z(n983) );
  XNOR2_X1 U1074 ( .A(G1986), .B(KEYINPUT114), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n983), .B(n982), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(n984), .B(G1971), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G1956), .B(G1961), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n986), .B(n985), .ZN(n987) );
  XOR2_X1 U1079 ( .A(n988), .B(n987), .Z(n990) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G1996), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(n992), .B(n991), .ZN(G229) );
  XOR2_X1 U1083 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n994) );
  XNOR2_X1 U1084 ( .A(KEYINPUT46), .B(KEYINPUT116), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(n994), .B(n993), .ZN(n995) );
  XOR2_X1 U1086 ( .A(n995), .B(G162), .Z(n998) );
  XNOR2_X1 U1087 ( .A(G164), .B(n996), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n998), .B(n997), .ZN(n1013) );
  NAND2_X1 U1089 ( .A1(G118), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(G130), .A2(n1000), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1009) );
  NAND2_X1 U1092 ( .A1(G142), .A2(n1003), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(G106), .A2(n1004), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(n1007), .B(KEYINPUT45), .Z(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XOR2_X1 U1097 ( .A(n1011), .B(n1010), .Z(n1012) );
  XOR2_X1 U1098 ( .A(n1013), .B(n1012), .Z(n1016) );
  XOR2_X1 U1099 ( .A(G160), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1100 ( .A(n1016), .B(n1015), .ZN(n1020) );
  XOR2_X1 U1101 ( .A(n1018), .B(n1017), .Z(n1019) );
  XNOR2_X1 U1102 ( .A(n1020), .B(n1019), .ZN(n1021) );
  NOR2_X1 U1103 ( .A1(G37), .A2(n1021), .ZN(G395) );
  INV_X1 U1104 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1105 ( .A(n1022), .B(G286), .Z(n1025) );
  XOR2_X1 U1106 ( .A(n1023), .B(G171), .Z(n1024) );
  XNOR2_X1 U1107 ( .A(n1025), .B(n1024), .ZN(n1026) );
  NOR2_X1 U1108 ( .A1(G37), .A2(n1026), .ZN(G397) );
  OR2_X1 U1109 ( .A1(G401), .A2(n1027), .ZN(n1030) );
  NOR2_X1 U1110 ( .A1(G227), .A2(G229), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(KEYINPUT49), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1112 ( .A1(n1030), .A2(n1029), .ZN(n1032) );
  NOR2_X1 U1113 ( .A1(G395), .A2(G397), .ZN(n1031) );
  NAND2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(G225) );
  INV_X1 U1115 ( .A(G225), .ZN(G308) );
  INV_X1 U1116 ( .A(G57), .ZN(G237) );
endmodule

