

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740;

  NOR2_X1 U371 ( .A1(n502), .A2(n512), .ZN(n503) );
  XNOR2_X1 U372 ( .A(n416), .B(G472), .ZN(n483) );
  XNOR2_X1 U373 ( .A(n365), .B(n364), .ZN(n625) );
  INV_X1 U374 ( .A(n360), .ZN(n351) );
  XNOR2_X1 U375 ( .A(n435), .B(n376), .ZN(n464) );
  BUF_X1 U376 ( .A(G128), .Z(n350) );
  AND2_X4 U377 ( .A1(n650), .A2(n355), .ZN(n698) );
  XNOR2_X2 U378 ( .A(n475), .B(n351), .ZN(n359) );
  XNOR2_X2 U379 ( .A(n440), .B(n391), .ZN(n475) );
  XOR2_X1 U380 ( .A(n685), .B(n684), .Z(n352) );
  BUF_X2 U381 ( .A(n483), .Z(n583) );
  XNOR2_X2 U382 ( .A(n404), .B(n403), .ZN(n582) );
  XNOR2_X2 U383 ( .A(n504), .B(KEYINPUT1), .ZN(n358) );
  INV_X1 U384 ( .A(KEYINPUT69), .ZN(n360) );
  NAND2_X1 U385 ( .A1(n605), .A2(n603), .ZN(n355) );
  XNOR2_X1 U386 ( .A(n366), .B(n388), .ZN(n484) );
  XNOR2_X1 U387 ( .A(n415), .B(n400), .ZN(n694) );
  INV_X1 U388 ( .A(G953), .ZN(n730) );
  BUF_X1 U389 ( .A(n698), .Z(n353) );
  NOR2_X2 U390 ( .A1(n554), .A2(n591), .ZN(n556) );
  NOR2_X2 U391 ( .A1(n369), .A2(n367), .ZN(n650) );
  NOR2_X1 U392 ( .A1(n680), .A2(G902), .ZN(n366) );
  INV_X1 U393 ( .A(KEYINPUT68), .ZN(n364) );
  NAND2_X1 U394 ( .A1(n484), .A2(n620), .ZN(n365) );
  INV_X1 U395 ( .A(G146), .ZN(n395) );
  XNOR2_X1 U396 ( .A(G110), .B(G107), .ZN(n396) );
  INV_X1 U397 ( .A(KEYINPUT39), .ZN(n451) );
  XNOR2_X1 U398 ( .A(G116), .B(G113), .ZN(n406) );
  XOR2_X1 U399 ( .A(G104), .B(KEYINPUT11), .Z(n454) );
  XNOR2_X1 U400 ( .A(n381), .B(n372), .ZN(n383) );
  XNOR2_X1 U401 ( .A(n373), .B(KEYINPUT96), .ZN(n372) );
  XNOR2_X1 U402 ( .A(KEYINPUT24), .B(G110), .ZN(n373) );
  NAND2_X1 U403 ( .A1(n668), .A2(n371), .ZN(n368) );
  XNOR2_X1 U404 ( .A(n563), .B(KEYINPUT33), .ZN(n641) );
  NAND2_X1 U405 ( .A1(n363), .A2(n362), .ZN(n361) );
  INV_X1 U406 ( .A(n590), .ZN(n362) );
  XNOR2_X1 U407 ( .A(n541), .B(KEYINPUT110), .ZN(n363) );
  NOR2_X1 U408 ( .A1(n588), .A2(n621), .ZN(n541) );
  XNOR2_X1 U409 ( .A(n428), .B(KEYINPUT75), .ZN(n508) );
  NAND2_X1 U410 ( .A1(n427), .A2(n354), .ZN(n428) );
  NOR2_X1 U411 ( .A1(n730), .A2(G952), .ZN(n704) );
  NOR2_X1 U412 ( .A1(G953), .A2(n609), .ZN(n645) );
  XNOR2_X1 U413 ( .A(n570), .B(n569), .ZN(n667) );
  XNOR2_X1 U414 ( .A(n556), .B(n555), .ZN(n666) );
  INV_X1 U415 ( .A(KEYINPUT32), .ZN(n555) );
  XNOR2_X1 U416 ( .A(n361), .B(KEYINPUT78), .ZN(n554) );
  INV_X1 U417 ( .A(n557), .ZN(n356) );
  AND2_X1 U418 ( .A1(n426), .A2(n486), .ZN(n354) );
  INV_X1 U419 ( .A(n358), .ZN(n588) );
  NAND2_X1 U420 ( .A1(n606), .A2(n355), .ZN(n607) );
  NAND2_X1 U421 ( .A1(n358), .A2(n625), .ZN(n579) );
  AND2_X1 U422 ( .A1(n588), .A2(n356), .ZN(n558) );
  AND2_X1 U423 ( .A1(n588), .A2(n357), .ZN(n626) );
  INV_X1 U424 ( .A(n625), .ZN(n357) );
  NOR2_X1 U425 ( .A1(n530), .A2(n358), .ZN(n531) );
  NAND2_X1 U426 ( .A1(n505), .A2(n358), .ZN(n725) );
  XNOR2_X2 U427 ( .A(n728), .B(n395), .ZN(n415) );
  XNOR2_X2 U428 ( .A(n359), .B(n394), .ZN(n728) );
  NAND2_X1 U429 ( .A1(n368), .A2(n444), .ZN(n367) );
  AND2_X2 U430 ( .A1(n370), .A2(n371), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n648), .B(KEYINPUT73), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n602), .B(n601), .ZN(n668) );
  INV_X1 U433 ( .A(KEYINPUT2), .ZN(n371) );
  BUF_X1 U434 ( .A(n484), .Z(n557) );
  XOR2_X1 U435 ( .A(n410), .B(n409), .Z(n374) );
  XOR2_X1 U436 ( .A(n651), .B(n653), .Z(n375) );
  XNOR2_X1 U437 ( .A(n374), .B(n412), .ZN(n413) );
  XNOR2_X1 U438 ( .A(n429), .B(n413), .ZN(n414) );
  XNOR2_X1 U439 ( .A(n415), .B(n414), .ZN(n651) );
  XNOR2_X1 U440 ( .A(n397), .B(G101), .ZN(n398) );
  OR2_X1 U441 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U442 ( .A(G902), .ZN(n480) );
  XNOR2_X1 U443 ( .A(n399), .B(n398), .ZN(n400) );
  BUF_X1 U444 ( .A(n648), .Z(n729) );
  INV_X1 U445 ( .A(n704), .ZN(n655) );
  XNOR2_X1 U446 ( .A(n647), .B(n646), .ZN(G75) );
  XNOR2_X1 U447 ( .A(KEYINPUT23), .B(KEYINPUT95), .ZN(n377) );
  XNOR2_X2 U448 ( .A(G146), .B(G125), .ZN(n435) );
  INV_X1 U449 ( .A(KEYINPUT10), .ZN(n376) );
  XNOR2_X1 U450 ( .A(n377), .B(n464), .ZN(n380) );
  NAND2_X1 U451 ( .A1(G234), .A2(n730), .ZN(n378) );
  XOR2_X1 U452 ( .A(KEYINPUT8), .B(n378), .Z(n476) );
  NAND2_X1 U453 ( .A1(n476), .A2(G221), .ZN(n379) );
  XNOR2_X1 U454 ( .A(n380), .B(n379), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n350), .B(G140), .ZN(n381) );
  XNOR2_X1 U456 ( .A(G119), .B(G137), .ZN(n382) );
  XNOR2_X1 U457 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U458 ( .A(n385), .B(n384), .ZN(n680) );
  XNOR2_X1 U459 ( .A(G902), .B(KEYINPUT15), .ZN(n649) );
  NAND2_X1 U460 ( .A1(G234), .A2(n649), .ZN(n386) );
  XNOR2_X1 U461 ( .A(KEYINPUT20), .B(n386), .ZN(n389) );
  NAND2_X1 U462 ( .A1(G217), .A2(n389), .ZN(n387) );
  XNOR2_X1 U463 ( .A(KEYINPUT25), .B(n387), .ZN(n388) );
  AND2_X1 U464 ( .A1(n389), .A2(G221), .ZN(n390) );
  XNOR2_X1 U465 ( .A(n390), .B(KEYINPUT21), .ZN(n620) );
  XNOR2_X2 U466 ( .A(G143), .B(G128), .ZN(n440) );
  INV_X1 U467 ( .A(G134), .ZN(n391) );
  INV_X1 U468 ( .A(KEYINPUT65), .ZN(n393) );
  XNOR2_X1 U469 ( .A(n393), .B(KEYINPUT4), .ZN(n436) );
  XNOR2_X1 U470 ( .A(G137), .B(n436), .ZN(n394) );
  XNOR2_X1 U471 ( .A(n396), .B(G104), .ZN(n431) );
  XOR2_X1 U472 ( .A(G131), .B(G140), .Z(n465) );
  XNOR2_X1 U473 ( .A(n431), .B(n465), .ZN(n399) );
  NAND2_X1 U474 ( .A1(G227), .A2(n730), .ZN(n397) );
  NAND2_X1 U475 ( .A1(n694), .A2(n480), .ZN(n402) );
  XOR2_X1 U476 ( .A(KEYINPUT71), .B(G469), .Z(n401) );
  XNOR2_X2 U477 ( .A(n402), .B(n401), .ZN(n504) );
  NAND2_X1 U478 ( .A1(n625), .A2(n504), .ZN(n404) );
  INV_X1 U479 ( .A(KEYINPUT97), .ZN(n403) );
  INV_X1 U480 ( .A(n582), .ZN(n427) );
  INV_X1 U481 ( .A(G119), .ZN(n405) );
  XNOR2_X1 U482 ( .A(n406), .B(n405), .ZN(n408) );
  XNOR2_X1 U483 ( .A(G101), .B(KEYINPUT3), .ZN(n407) );
  XNOR2_X1 U484 ( .A(n408), .B(n407), .ZN(n429) );
  XOR2_X1 U485 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n410) );
  XNOR2_X1 U486 ( .A(G131), .B(KEYINPUT98), .ZN(n409) );
  NOR2_X1 U487 ( .A1(G237), .A2(G953), .ZN(n411) );
  XNOR2_X1 U488 ( .A(n411), .B(KEYINPUT74), .ZN(n461) );
  NAND2_X1 U489 ( .A1(G210), .A2(n461), .ZN(n412) );
  NAND2_X1 U490 ( .A1(n651), .A2(n480), .ZN(n416) );
  NOR2_X1 U491 ( .A1(G237), .A2(G902), .ZN(n417) );
  XNOR2_X1 U492 ( .A(n417), .B(KEYINPUT72), .ZN(n446) );
  INV_X1 U493 ( .A(G214), .ZN(n418) );
  OR2_X1 U494 ( .A1(n446), .A2(n418), .ZN(n613) );
  NAND2_X1 U495 ( .A1(n483), .A2(n613), .ZN(n420) );
  XNOR2_X1 U496 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n419) );
  XNOR2_X1 U497 ( .A(n420), .B(n419), .ZN(n426) );
  NAND2_X1 U498 ( .A1(G234), .A2(G237), .ZN(n421) );
  XNOR2_X1 U499 ( .A(n421), .B(KEYINPUT14), .ZN(n423) );
  NAND2_X1 U500 ( .A1(G952), .A2(n423), .ZN(n638) );
  NOR2_X1 U501 ( .A1(n638), .A2(G953), .ZN(n422) );
  XOR2_X1 U502 ( .A(n422), .B(KEYINPUT92), .Z(n545) );
  NAND2_X1 U503 ( .A1(G902), .A2(n423), .ZN(n543) );
  NOR2_X1 U504 ( .A1(G900), .A2(n543), .ZN(n424) );
  NAND2_X1 U505 ( .A1(G953), .A2(n424), .ZN(n425) );
  NAND2_X1 U506 ( .A1(n545), .A2(n425), .ZN(n486) );
  INV_X1 U507 ( .A(n429), .ZN(n433) );
  XNOR2_X1 U508 ( .A(KEYINPUT16), .B(G122), .ZN(n430) );
  XNOR2_X1 U509 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U510 ( .A(n433), .B(n432), .ZN(n676) );
  XNOR2_X1 U511 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n434) );
  XNOR2_X1 U512 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U513 ( .A(n437), .B(n436), .ZN(n442) );
  NAND2_X1 U514 ( .A1(n730), .A2(G224), .ZN(n438) );
  XNOR2_X1 U515 ( .A(n438), .B(KEYINPUT90), .ZN(n439) );
  XNOR2_X1 U516 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U517 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U518 ( .A(n676), .B(n443), .ZN(n701) );
  INV_X1 U519 ( .A(n649), .ZN(n444) );
  OR2_X1 U520 ( .A1(n701), .A2(n444), .ZN(n450) );
  INV_X1 U521 ( .A(G210), .ZN(n445) );
  OR2_X1 U522 ( .A1(n446), .A2(n445), .ZN(n448) );
  INV_X1 U523 ( .A(KEYINPUT91), .ZN(n447) );
  XNOR2_X1 U524 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X2 U525 ( .A(n450), .B(n449), .ZN(n533) );
  XNOR2_X1 U526 ( .A(n533), .B(KEYINPUT38), .ZN(n614) );
  NAND2_X1 U527 ( .A1(n508), .A2(n614), .ZN(n452) );
  XNOR2_X2 U528 ( .A(n452), .B(n451), .ZN(n529) );
  XNOR2_X1 U529 ( .A(G143), .B(KEYINPUT103), .ZN(n453) );
  XNOR2_X1 U530 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U531 ( .A(n455), .B(G122), .Z(n460) );
  XOR2_X1 U532 ( .A(KEYINPUT102), .B(KEYINPUT104), .Z(n457) );
  XNOR2_X1 U533 ( .A(KEYINPUT101), .B(KEYINPUT12), .ZN(n456) );
  XNOR2_X1 U534 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U535 ( .A(G113), .B(n458), .ZN(n459) );
  XNOR2_X1 U536 ( .A(n460), .B(n459), .ZN(n463) );
  NAND2_X1 U537 ( .A1(n461), .A2(G214), .ZN(n462) );
  XNOR2_X1 U538 ( .A(n463), .B(n462), .ZN(n466) );
  XOR2_X1 U539 ( .A(n465), .B(n464), .Z(n727) );
  XNOR2_X1 U540 ( .A(n466), .B(n727), .ZN(n687) );
  NAND2_X1 U541 ( .A1(n687), .A2(n480), .ZN(n468) );
  XNOR2_X1 U542 ( .A(KEYINPUT13), .B(G475), .ZN(n467) );
  XNOR2_X1 U543 ( .A(n468), .B(n467), .ZN(n516) );
  XOR2_X1 U544 ( .A(KEYINPUT7), .B(G107), .Z(n470) );
  XNOR2_X1 U545 ( .A(G116), .B(G122), .ZN(n469) );
  XNOR2_X1 U546 ( .A(n470), .B(n469), .ZN(n474) );
  XOR2_X1 U547 ( .A(KEYINPUT105), .B(KEYINPUT9), .Z(n472) );
  XNOR2_X1 U548 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n471) );
  XNOR2_X1 U549 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U550 ( .A(n474), .B(n473), .Z(n479) );
  AND2_X1 U551 ( .A1(G217), .A2(n476), .ZN(n477) );
  XNOR2_X1 U552 ( .A(n475), .B(n477), .ZN(n478) );
  XNOR2_X1 U553 ( .A(n479), .B(n478), .ZN(n685) );
  NAND2_X1 U554 ( .A1(n685), .A2(n480), .ZN(n481) );
  XNOR2_X1 U555 ( .A(n481), .B(G478), .ZN(n515) );
  OR2_X1 U556 ( .A1(n516), .A2(n515), .ZN(n720) );
  NOR2_X2 U557 ( .A1(n529), .A2(n720), .ZN(n482) );
  XNOR2_X1 U558 ( .A(n482), .B(KEYINPUT40), .ZN(n738) );
  INV_X1 U559 ( .A(n620), .ZN(n485) );
  NOR2_X1 U560 ( .A1(n485), .A2(n557), .ZN(n487) );
  NAND2_X1 U561 ( .A1(n487), .A2(n486), .ZN(n499) );
  INV_X1 U562 ( .A(n499), .ZN(n488) );
  NAND2_X1 U563 ( .A1(n583), .A2(n488), .ZN(n489) );
  XNOR2_X1 U564 ( .A(n489), .B(KEYINPUT28), .ZN(n491) );
  INV_X1 U565 ( .A(n504), .ZN(n490) );
  OR2_X1 U566 ( .A1(n491), .A2(n490), .ZN(n510) );
  NAND2_X1 U567 ( .A1(n614), .A2(n613), .ZN(n493) );
  INV_X1 U568 ( .A(KEYINPUT113), .ZN(n492) );
  XNOR2_X1 U569 ( .A(n493), .B(n492), .ZN(n612) );
  INV_X1 U570 ( .A(n516), .ZN(n506) );
  OR2_X1 U571 ( .A1(n506), .A2(n515), .ZN(n615) );
  OR2_X1 U572 ( .A1(n612), .A2(n615), .ZN(n495) );
  INV_X1 U573 ( .A(KEYINPUT41), .ZN(n494) );
  XNOR2_X1 U574 ( .A(n495), .B(n494), .ZN(n639) );
  NOR2_X1 U575 ( .A1(n510), .A2(n639), .ZN(n496) );
  XNOR2_X1 U576 ( .A(n496), .B(KEYINPUT42), .ZN(n661) );
  NOR2_X1 U577 ( .A1(n738), .A2(n661), .ZN(n497) );
  XNOR2_X1 U578 ( .A(n497), .B(KEYINPUT46), .ZN(n526) );
  INV_X1 U579 ( .A(KEYINPUT6), .ZN(n498) );
  XNOR2_X2 U580 ( .A(n583), .B(n498), .ZN(n590) );
  NOR2_X1 U581 ( .A1(n720), .A2(n499), .ZN(n500) );
  NAND2_X1 U582 ( .A1(n590), .A2(n500), .ZN(n530) );
  XNOR2_X1 U583 ( .A(KEYINPUT114), .B(n530), .ZN(n502) );
  INV_X1 U584 ( .A(n613), .ZN(n501) );
  OR2_X2 U585 ( .A1(n533), .A2(n501), .ZN(n512) );
  XNOR2_X1 U586 ( .A(n503), .B(KEYINPUT36), .ZN(n505) );
  XOR2_X1 U587 ( .A(KEYINPUT86), .B(n725), .Z(n524) );
  NAND2_X1 U588 ( .A1(n506), .A2(n515), .ZN(n566) );
  NOR2_X1 U589 ( .A1(n566), .A2(n533), .ZN(n507) );
  NAND2_X1 U590 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U591 ( .A(n509), .B(KEYINPUT112), .ZN(n740) );
  INV_X1 U592 ( .A(n510), .ZN(n513) );
  XNOR2_X1 U593 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n511) );
  XNOR2_X1 U594 ( .A(n512), .B(n511), .ZN(n547) );
  AND2_X1 U595 ( .A1(n513), .A2(n547), .ZN(n722) );
  NOR2_X1 U596 ( .A1(n722), .A2(KEYINPUT47), .ZN(n521) );
  INV_X1 U597 ( .A(n722), .ZN(n519) );
  INV_X1 U598 ( .A(KEYINPUT47), .ZN(n514) );
  NAND2_X1 U599 ( .A1(n514), .A2(KEYINPUT82), .ZN(n517) );
  NAND2_X1 U600 ( .A1(n516), .A2(n515), .ZN(n716) );
  NAND2_X1 U601 ( .A1(n716), .A2(n720), .ZN(n610) );
  XOR2_X1 U602 ( .A(n517), .B(n610), .Z(n518) );
  NOR2_X1 U603 ( .A1(n519), .A2(n518), .ZN(n520) );
  OR2_X1 U604 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U605 ( .A1(n740), .A2(n522), .ZN(n523) );
  NOR2_X1 U606 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U607 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U608 ( .A(KEYINPUT70), .B(KEYINPUT48), .ZN(n527) );
  XNOR2_X2 U609 ( .A(n528), .B(n527), .ZN(n537) );
  OR2_X1 U610 ( .A1(n529), .A2(n716), .ZN(n726) );
  NAND2_X1 U611 ( .A1(n531), .A2(n613), .ZN(n532) );
  XNOR2_X1 U612 ( .A(n532), .B(KEYINPUT43), .ZN(n534) );
  NAND2_X1 U613 ( .A1(n534), .A2(n533), .ZN(n662) );
  NAND2_X1 U614 ( .A1(n726), .A2(n662), .ZN(n535) );
  NOR2_X2 U615 ( .A1(n537), .A2(n535), .ZN(n648) );
  XOR2_X1 U616 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n604) );
  NOR2_X1 U617 ( .A1(n729), .A2(n604), .ZN(n536) );
  XOR2_X1 U618 ( .A(KEYINPUT83), .B(n536), .Z(n608) );
  NAND2_X1 U619 ( .A1(n726), .A2(KEYINPUT2), .ZN(n538) );
  XNOR2_X1 U620 ( .A(n538), .B(KEYINPUT79), .ZN(n539) );
  NAND2_X1 U621 ( .A1(n539), .A2(n662), .ZN(n540) );
  NOR2_X1 U622 ( .A1(n537), .A2(n540), .ZN(n603) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT108), .ZN(n621) );
  XNOR2_X1 U624 ( .A(G898), .B(KEYINPUT93), .ZN(n671) );
  NAND2_X1 U625 ( .A1(n671), .A2(G953), .ZN(n542) );
  XNOR2_X1 U626 ( .A(n542), .B(KEYINPUT94), .ZN(n674) );
  OR2_X1 U627 ( .A1(n674), .A2(n543), .ZN(n544) );
  NAND2_X1 U628 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U629 ( .A1(n547), .A2(n546), .ZN(n549) );
  XNOR2_X1 U630 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n548) );
  XNOR2_X2 U631 ( .A(n549), .B(n548), .ZN(n584) );
  INV_X1 U632 ( .A(n584), .ZN(n552) );
  INV_X1 U633 ( .A(n615), .ZN(n550) );
  NAND2_X1 U634 ( .A1(n550), .A2(n620), .ZN(n551) );
  OR2_X1 U635 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X2 U636 ( .A(n553), .B(KEYINPUT22), .ZN(n591) );
  INV_X1 U637 ( .A(n583), .ZN(n624) );
  NAND2_X1 U638 ( .A1(n624), .A2(n558), .ZN(n559) );
  NOR2_X1 U639 ( .A1(n591), .A2(n559), .ZN(n659) );
  INV_X1 U640 ( .A(KEYINPUT44), .ZN(n560) );
  NOR2_X1 U641 ( .A1(n659), .A2(n560), .ZN(n561) );
  NAND2_X1 U642 ( .A1(n666), .A2(n561), .ZN(n572) );
  INV_X1 U643 ( .A(n579), .ZN(n562) );
  NAND2_X1 U644 ( .A1(n590), .A2(n562), .ZN(n563) );
  NAND2_X1 U645 ( .A1(n641), .A2(n584), .ZN(n565) );
  XNOR2_X1 U646 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n564) );
  XNOR2_X1 U647 ( .A(n565), .B(n564), .ZN(n568) );
  INV_X1 U648 ( .A(n566), .ZN(n567) );
  NAND2_X1 U649 ( .A1(n568), .A2(n567), .ZN(n570) );
  XOR2_X1 U650 ( .A(KEYINPUT76), .B(KEYINPUT35), .Z(n569) );
  NOR2_X1 U651 ( .A1(n667), .A2(KEYINPUT87), .ZN(n571) );
  NOR2_X1 U652 ( .A1(n572), .A2(n571), .ZN(n574) );
  NOR2_X1 U653 ( .A1(KEYINPUT87), .A2(KEYINPUT44), .ZN(n573) );
  NOR2_X1 U654 ( .A1(n574), .A2(n573), .ZN(n599) );
  NOR2_X1 U655 ( .A1(n659), .A2(KEYINPUT44), .ZN(n575) );
  NAND2_X1 U656 ( .A1(n666), .A2(n575), .ZN(n577) );
  INV_X1 U657 ( .A(KEYINPUT87), .ZN(n576) );
  NAND2_X1 U658 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U659 ( .A1(n578), .A2(n667), .ZN(n597) );
  NOR2_X1 U660 ( .A1(n624), .A2(n579), .ZN(n630) );
  NAND2_X1 U661 ( .A1(n630), .A2(n584), .ZN(n581) );
  XOR2_X1 U662 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n580) );
  XNOR2_X1 U663 ( .A(n581), .B(n580), .ZN(n664) );
  NOR2_X1 U664 ( .A1(n582), .A2(n583), .ZN(n585) );
  NAND2_X1 U665 ( .A1(n585), .A2(n584), .ZN(n713) );
  NAND2_X1 U666 ( .A1(n664), .A2(n713), .ZN(n587) );
  XNOR2_X1 U667 ( .A(n610), .B(KEYINPUT82), .ZN(n586) );
  NAND2_X1 U668 ( .A1(n587), .A2(n586), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n621), .A2(n588), .ZN(n589) );
  NOR2_X1 U670 ( .A1(n590), .A2(n589), .ZN(n593) );
  INV_X1 U671 ( .A(n591), .ZN(n592) );
  NAND2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n658) );
  NAND2_X1 U673 ( .A1(n594), .A2(n658), .ZN(n595) );
  XNOR2_X1 U674 ( .A(n595), .B(KEYINPUT109), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n602) );
  XNOR2_X1 U677 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n600) );
  XNOR2_X1 U678 ( .A(n600), .B(KEYINPUT64), .ZN(n601) );
  INV_X1 U679 ( .A(n668), .ZN(n605) );
  NOR2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  INV_X1 U681 ( .A(n610), .ZN(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n618) );
  NOR2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n616) );
  NOR2_X1 U684 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U686 ( .A1(n619), .A2(n641), .ZN(n635) );
  NOR2_X1 U687 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U688 ( .A(n622), .B(KEYINPUT49), .ZN(n623) );
  NAND2_X1 U689 ( .A1(n624), .A2(n623), .ZN(n628) );
  XNOR2_X1 U690 ( .A(n626), .B(KEYINPUT50), .ZN(n627) );
  NOR2_X1 U691 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U692 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U693 ( .A(KEYINPUT51), .B(n631), .Z(n632) );
  NOR2_X1 U694 ( .A1(n632), .A2(n639), .ZN(n633) );
  XOR2_X1 U695 ( .A(n633), .B(KEYINPUT118), .Z(n634) );
  NAND2_X1 U696 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U697 ( .A(KEYINPUT52), .B(n636), .Z(n637) );
  NOR2_X1 U698 ( .A1(n638), .A2(n637), .ZN(n643) );
  INV_X1 U699 ( .A(n639), .ZN(n640) );
  AND2_X1 U700 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U701 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U702 ( .A1(n645), .A2(n644), .ZN(n647) );
  XNOR2_X1 U703 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n646) );
  NAND2_X1 U704 ( .A1(n698), .A2(G472), .ZN(n654) );
  XNOR2_X1 U705 ( .A(KEYINPUT88), .B(KEYINPUT115), .ZN(n652) );
  XNOR2_X1 U706 ( .A(n652), .B(KEYINPUT62), .ZN(n653) );
  XNOR2_X1 U707 ( .A(n654), .B(n375), .ZN(n656) );
  NAND2_X1 U708 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U709 ( .A(n657), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U710 ( .A(n658), .B(G101), .ZN(G3) );
  XOR2_X1 U711 ( .A(G110), .B(n659), .Z(G12) );
  XNOR2_X1 U712 ( .A(G137), .B(KEYINPUT125), .ZN(n660) );
  XNOR2_X1 U713 ( .A(n661), .B(n660), .ZN(G39) );
  XNOR2_X1 U714 ( .A(n662), .B(G140), .ZN(G42) );
  NOR2_X1 U715 ( .A1(n664), .A2(n720), .ZN(n663) );
  XOR2_X1 U716 ( .A(G113), .B(n663), .Z(G15) );
  NOR2_X1 U717 ( .A1(n664), .A2(n716), .ZN(n665) );
  XOR2_X1 U718 ( .A(G116), .B(n665), .Z(G18) );
  XNOR2_X1 U719 ( .A(n666), .B(G119), .ZN(G21) );
  XNOR2_X1 U720 ( .A(n667), .B(G122), .ZN(G24) );
  NOR2_X1 U721 ( .A1(n668), .A2(G953), .ZN(n673) );
  NAND2_X1 U722 ( .A1(G953), .A2(G224), .ZN(n669) );
  XOR2_X1 U723 ( .A(KEYINPUT61), .B(n669), .Z(n670) );
  NOR2_X1 U724 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U725 ( .A1(n673), .A2(n672), .ZN(n679) );
  INV_X1 U726 ( .A(n674), .ZN(n675) );
  NOR2_X1 U727 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U728 ( .A(n677), .B(KEYINPUT123), .ZN(n678) );
  XNOR2_X1 U729 ( .A(n679), .B(n678), .ZN(G69) );
  NAND2_X1 U730 ( .A1(n353), .A2(G217), .ZN(n682) );
  XNOR2_X1 U731 ( .A(n680), .B(KEYINPUT122), .ZN(n681) );
  XNOR2_X1 U732 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U733 ( .A1(n683), .A2(n704), .ZN(G66) );
  NAND2_X1 U734 ( .A1(n698), .A2(G478), .ZN(n684) );
  NOR2_X1 U735 ( .A1(n352), .A2(n704), .ZN(G63) );
  NAND2_X1 U736 ( .A1(n698), .A2(G475), .ZN(n689) );
  XOR2_X1 U737 ( .A(KEYINPUT89), .B(KEYINPUT59), .Z(n686) );
  XNOR2_X1 U738 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U739 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X2 U740 ( .A1(n690), .A2(n704), .ZN(n692) );
  XOR2_X1 U741 ( .A(KEYINPUT121), .B(KEYINPUT60), .Z(n691) );
  XNOR2_X1 U742 ( .A(n692), .B(n691), .ZN(G60) );
  NAND2_X1 U743 ( .A1(n353), .A2(G469), .ZN(n696) );
  XNOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n693) );
  XNOR2_X1 U745 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U746 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U747 ( .A1(n697), .A2(n704), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n698), .A2(G210), .ZN(n703) );
  XOR2_X1 U749 ( .A(KEYINPUT80), .B(KEYINPUT54), .Z(n699) );
  XNOR2_X1 U750 ( .A(n699), .B(KEYINPUT55), .ZN(n700) );
  XNOR2_X1 U751 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U752 ( .A(n703), .B(n702), .ZN(n705) );
  NOR2_X2 U753 ( .A1(n705), .A2(n704), .ZN(n708) );
  XNOR2_X1 U754 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n706) );
  XOR2_X1 U755 ( .A(n706), .B(KEYINPUT85), .Z(n707) );
  XNOR2_X1 U756 ( .A(n708), .B(n707), .ZN(G51) );
  OR2_X1 U757 ( .A1(n713), .A2(n720), .ZN(n709) );
  XNOR2_X1 U758 ( .A(n709), .B(G104), .ZN(G6) );
  XOR2_X1 U759 ( .A(KEYINPUT117), .B(KEYINPUT27), .Z(n711) );
  XNOR2_X1 U760 ( .A(G107), .B(KEYINPUT26), .ZN(n710) );
  XNOR2_X1 U761 ( .A(n711), .B(n710), .ZN(n712) );
  XOR2_X1 U762 ( .A(KEYINPUT116), .B(n712), .Z(n715) );
  OR2_X1 U763 ( .A1(n713), .A2(n716), .ZN(n714) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(G9) );
  XOR2_X1 U765 ( .A(n350), .B(KEYINPUT29), .Z(n719) );
  INV_X1 U766 ( .A(n716), .ZN(n717) );
  NAND2_X1 U767 ( .A1(n722), .A2(n717), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(G30) );
  INV_X1 U769 ( .A(n720), .ZN(n721) );
  NAND2_X1 U770 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n723), .B(G146), .ZN(G48) );
  XOR2_X1 U772 ( .A(G125), .B(KEYINPUT37), .Z(n724) );
  XNOR2_X1 U773 ( .A(n725), .B(n724), .ZN(G27) );
  XNOR2_X1 U774 ( .A(G134), .B(n726), .ZN(G36) );
  XNOR2_X1 U775 ( .A(n728), .B(n727), .ZN(n732) );
  XOR2_X1 U776 ( .A(n732), .B(n729), .Z(n731) );
  NAND2_X1 U777 ( .A1(n731), .A2(n730), .ZN(n737) );
  XNOR2_X1 U778 ( .A(G227), .B(n732), .ZN(n733) );
  NAND2_X1 U779 ( .A1(n733), .A2(G900), .ZN(n734) );
  XNOR2_X1 U780 ( .A(KEYINPUT124), .B(n734), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U782 ( .A1(n737), .A2(n736), .ZN(G72) );
  XOR2_X1 U783 ( .A(G131), .B(KEYINPUT126), .Z(n739) );
  XNOR2_X1 U784 ( .A(n738), .B(n739), .ZN(G33) );
  XNOR2_X1 U785 ( .A(G143), .B(n740), .ZN(G45) );
endmodule

