//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OR2_X1    g0009(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n211));
  AND3_X1   g0011(.A1(new_n210), .A2(G50), .A3(new_n211), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n212), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n209), .B(new_n213), .C1(new_n220), .C2(KEYINPUT1), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0022(.A(G238), .B(G244), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(G232), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT2), .B(G226), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n226), .B(new_n229), .Z(G358));
  XOR2_X1   g0030(.A(G58), .B(G77), .Z(new_n231));
  XNOR2_X1  g0031(.A(G50), .B(G68), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XNOR2_X1  g0034(.A(G107), .B(G116), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G351));
  INV_X1    g0037(.A(G1), .ZN(new_n238));
  OAI21_X1  g0038(.A(new_n238), .B1(G41), .B2(G45), .ZN(new_n239));
  INV_X1    g0039(.A(G274), .ZN(new_n240));
  NOR2_X1   g0040(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(KEYINPUT66), .ZN(new_n242));
  NAND2_X1  g0042(.A1(G33), .A2(G41), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n243), .A2(G1), .A3(G13), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT66), .ZN(new_n245));
  OAI211_X1 g0045(.A(new_n245), .B(new_n238), .C1(G41), .C2(G45), .ZN(new_n246));
  AND3_X1   g0046(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n241), .B1(new_n247), .B2(G238), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  OAI211_X1 g0051(.A(G226), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  OAI211_X1 g0052(.A(G232), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G97), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT77), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT77), .A4(new_n254), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n244), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT78), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n248), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI211_X1 g0061(.A(KEYINPUT78), .B(new_n244), .C1(new_n257), .C2(new_n258), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT13), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n258), .ZN(new_n264));
  INV_X1    g0064(.A(new_n244), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT78), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT13), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n259), .A2(new_n260), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .A4(new_n248), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n263), .A2(new_n270), .A3(G190), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G1), .A2(G13), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n272), .A2(KEYINPUT67), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT67), .B1(new_n272), .B2(new_n273), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G68), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n277), .A2(G50), .B1(G20), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  INV_X1    g0080(.A(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT11), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n238), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n278), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT12), .ZN(new_n289));
  INV_X1    g0089(.A(new_n275), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n272), .A2(KEYINPUT67), .A3(new_n273), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(new_n291), .B1(new_n238), .B2(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G68), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n285), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n271), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n263), .B2(new_n270), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT79), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n248), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n266), .B2(KEYINPUT78), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n268), .B1(new_n301), .B2(new_n269), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n261), .A2(KEYINPUT13), .A3(new_n262), .ZN(new_n303));
  OAI21_X1  g0103(.A(G200), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT79), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(new_n295), .A4(new_n271), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT3), .B(G33), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(G222), .A3(new_n249), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(G223), .A3(G1698), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n310), .B(new_n311), .C1(new_n280), .C2(new_n309), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n265), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n241), .B1(new_n247), .B2(G226), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n315), .A2(G169), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT69), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n203), .A2(new_n317), .A3(G20), .ZN(new_n318));
  NOR3_X1   g0118(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT69), .B1(new_n319), .B2(new_n281), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n277), .A2(G150), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT68), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT68), .ZN(new_n325));
  INV_X1    g0125(.A(G58), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT8), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n324), .A2(new_n281), .A3(G33), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n276), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n286), .A2(G50), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n292), .B2(G50), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g0133(.A(KEYINPUT70), .B(G179), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n315), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n316), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT9), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(new_n337), .A3(new_n332), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n290), .A2(new_n291), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n322), .B2(new_n328), .ZN(new_n340));
  OAI221_X1 g0140(.A(G50), .B1(G1), .B2(new_n281), .C1(new_n274), .C2(new_n275), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G50), .B2(new_n286), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT9), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n313), .A2(new_n314), .A3(G190), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n297), .B1(new_n313), .B2(new_n314), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT10), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(new_n344), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n336), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G20), .A2(G77), .ZN(new_n352));
  INV_X1    g0152(.A(new_n277), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n352), .B1(new_n323), .B2(new_n353), .C1(new_n282), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n276), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n292), .A2(G77), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n286), .A2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT73), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n309), .A2(G238), .A3(G1698), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n309), .A2(G232), .A3(new_n249), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n250), .A2(new_n251), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT71), .B(G107), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n265), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n241), .B1(new_n247), .B2(G244), .ZN(new_n368));
  AOI21_X1  g0168(.A(G169), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT76), .B1(new_n360), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT76), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n367), .A2(new_n368), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(new_n372), .C1(new_n373), .C2(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n367), .A2(new_n368), .A3(new_n334), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(KEYINPUT75), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(KEYINPUT75), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n297), .B1(new_n367), .B2(new_n368), .ZN(new_n381));
  OR3_X1    g0181(.A1(new_n381), .A2(new_n372), .A3(KEYINPUT74), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n373), .A2(G190), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT72), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT74), .B1(new_n381), .B2(new_n372), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n373), .A2(KEYINPUT72), .A3(G190), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n380), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n351), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT3), .ZN(new_n391));
  INV_X1    g0191(.A(G33), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT3), .A2(G33), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n281), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT7), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n393), .A2(new_n397), .A3(new_n281), .A4(new_n394), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(G68), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  XNOR2_X1  g0200(.A(G58), .B(G68), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(G20), .B1(G159), .B2(new_n277), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n400), .B1(new_n399), .B2(new_n402), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n276), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n324), .A2(new_n327), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n238), .B2(G20), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n276), .A2(new_n287), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n407), .A2(new_n408), .B1(new_n287), .B2(new_n406), .ZN(new_n409));
  INV_X1    g0209(.A(new_n241), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n242), .A2(G232), .A3(new_n244), .A4(new_n246), .ZN(new_n411));
  INV_X1    g0211(.A(G87), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n392), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G223), .A2(G1698), .ZN(new_n414));
  INV_X1    g0214(.A(G226), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(G1698), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n413), .B1(new_n416), .B2(new_n309), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n410), .B(new_n411), .C1(new_n417), .C2(new_n244), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n297), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(G1698), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(G223), .B2(G1698), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n421), .A2(new_n363), .B1(new_n392), .B2(new_n412), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n265), .ZN(new_n423));
  INV_X1    g0223(.A(G190), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n410), .A4(new_n411), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n405), .A2(new_n409), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n405), .A2(new_n426), .A3(KEYINPUT17), .A4(new_n409), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G169), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n418), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n423), .A2(new_n410), .A3(new_n334), .A4(new_n411), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n399), .A2(new_n402), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT16), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n339), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n407), .A2(new_n408), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n406), .A2(new_n287), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n435), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT18), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n405), .A2(new_n409), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n435), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n431), .A2(KEYINPUT80), .A3(new_n444), .A4(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n444), .A2(new_n447), .A3(new_n429), .A4(new_n430), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n390), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(G169), .B1(new_n302), .B2(new_n303), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n302), .A2(new_n303), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n453), .A2(KEYINPUT14), .B1(new_n454), .B2(G179), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT14), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(G169), .C1(new_n302), .C2(new_n303), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n295), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n308), .A2(new_n452), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G41), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n238), .B(G45), .C1(new_n460), .C2(KEYINPUT5), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT81), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G41), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n465), .A2(KEYINPUT81), .A3(new_n238), .A4(G45), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n460), .A2(KEYINPUT5), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G270), .A3(new_n244), .ZN(new_n469));
  OAI211_X1 g0269(.A(G264), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n470));
  OAI211_X1 g0270(.A(G257), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n393), .A2(G303), .A3(new_n394), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n265), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n461), .A2(new_n462), .B1(KEYINPUT5), .B2(new_n460), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(G274), .A3(new_n244), .A4(new_n466), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n469), .A2(new_n474), .A3(G179), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT85), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n287), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n272), .A2(new_n273), .B1(G20), .B2(new_n479), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n482), .B(new_n281), .C1(G33), .C2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(KEYINPUT20), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT20), .B1(new_n481), .B2(new_n484), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n480), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n238), .A2(G33), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n286), .B(new_n489), .C1(new_n274), .C2(new_n275), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n479), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n478), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n487), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n485), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n339), .A2(G116), .A3(new_n286), .A4(new_n489), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT85), .A4(new_n480), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n477), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G169), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n492), .B2(new_n496), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n500), .B2(KEYINPUT21), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n492), .A2(new_n496), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n504), .B2(new_n499), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n498), .A2(G200), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n469), .A2(new_n474), .A3(G190), .A4(new_n476), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n506), .A2(new_n492), .A3(new_n496), .A4(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n508), .A2(KEYINPUT86), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(KEYINPUT86), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n501), .B(new_n505), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G244), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n309), .A2(KEYINPUT4), .A3(G244), .A4(new_n249), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n309), .A2(G250), .A3(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n482), .A4(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n518), .A2(new_n265), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n468), .A2(G257), .A3(new_n244), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n476), .ZN(new_n521));
  OAI21_X1  g0321(.A(G200), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT82), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n265), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n525), .A2(G190), .A3(new_n476), .A4(new_n520), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n286), .A2(G97), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n490), .B2(new_n483), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  AND2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n396), .A2(new_n398), .A3(new_n364), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n529), .B1(new_n539), .B2(new_n276), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n526), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n525), .A2(new_n476), .A3(new_n520), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(KEYINPUT82), .A3(G200), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n524), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n432), .B1(new_n519), .B2(new_n521), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n520), .A2(new_n476), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(new_n334), .A3(new_n525), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n539), .A2(new_n276), .ZN(new_n548));
  INV_X1    g0348(.A(new_n529), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n552));
  OAI211_X1 g0352(.A(G238), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G116), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n265), .ZN(new_n556));
  INV_X1    g0356(.A(G45), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT83), .B1(new_n557), .B2(G1), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT83), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(new_n238), .A3(G45), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n244), .A2(new_n558), .A3(new_n560), .A4(G250), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n238), .A2(G45), .A3(G274), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n561), .A2(KEYINPUT84), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT84), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n556), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n282), .B2(new_n483), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n281), .A2(G68), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n363), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(KEYINPUT71), .A2(G107), .ZN(new_n571));
  NOR2_X1   g0371(.A1(KEYINPUT71), .A2(G107), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G87), .A2(G97), .ZN(new_n574));
  NAND3_X1  g0374(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n573), .A2(new_n574), .B1(new_n281), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n276), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n339), .A2(G87), .A3(new_n286), .A4(new_n489), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n354), .A2(new_n287), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n556), .B(G190), .C1(new_n563), .C2(new_n564), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n566), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n556), .B(new_n334), .C1(new_n563), .C2(new_n564), .ZN(new_n583));
  INV_X1    g0383(.A(new_n354), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n339), .A2(new_n286), .A3(new_n584), .A4(new_n489), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n577), .A2(new_n585), .A3(new_n579), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n561), .A2(new_n562), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT84), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n561), .A2(KEYINPUT84), .A3(new_n562), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n589), .A2(new_n590), .B1(new_n265), .B2(new_n555), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n583), .B(new_n586), .C1(new_n591), .C2(G169), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n582), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n544), .A2(new_n551), .A3(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(KEYINPUT22), .B(G87), .C1(new_n250), .C2(new_n251), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT23), .B1(new_n571), .B2(new_n572), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n595), .A2(new_n596), .B1(new_n597), .B2(G20), .ZN(new_n598));
  OAI21_X1  g0398(.A(G87), .B1(new_n250), .B2(new_n251), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT22), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT24), .B1(new_n598), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT24), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n599), .A2(new_n600), .B1(G20), .B2(new_n602), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n595), .A2(new_n596), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n281), .B1(new_n364), .B2(KEYINPUT23), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n606), .B(new_n607), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n276), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n286), .A2(G107), .ZN(new_n613));
  XOR2_X1   g0413(.A(new_n613), .B(KEYINPUT25), .Z(new_n614));
  INV_X1    g0414(.A(new_n490), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(G107), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(G250), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n618));
  OAI211_X1 g0418(.A(G257), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n619));
  XOR2_X1   g0419(.A(KEYINPUT87), .B(G294), .Z(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n392), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n265), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n468), .A2(G264), .A3(new_n244), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(new_n476), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT88), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n625), .A3(G169), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n265), .B1(new_n475), .B2(new_n466), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(G264), .B1(new_n621), .B2(new_n265), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(G179), .A3(new_n476), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n625), .B1(new_n624), .B2(G169), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n617), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(G200), .B1(new_n628), .B2(new_n476), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n624), .A2(G190), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n612), .B(new_n616), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n594), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n459), .A2(new_n512), .A3(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n336), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT91), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n433), .A2(new_n434), .ZN(new_n641));
  AOI211_X1 g0441(.A(KEYINPUT18), .B(new_n641), .C1(new_n405), .C2(new_n409), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n446), .B1(new_n445), .B2(new_n435), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n444), .A2(KEYINPUT91), .A3(new_n447), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n453), .A2(KEYINPUT14), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n454), .A2(G179), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n457), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n304), .A2(new_n295), .A3(new_n271), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n370), .A2(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n649), .A2(new_n294), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n431), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n646), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n349), .A2(new_n350), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n639), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n501), .A2(new_n505), .A3(new_n632), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n545), .A2(new_n550), .A3(new_n547), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT82), .B1(new_n542), .B2(G200), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n526), .A2(new_n540), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n658), .B1(new_n543), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT89), .B1(new_n591), .B2(new_n297), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT89), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n565), .A2(new_n664), .A3(G200), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n663), .A2(new_n581), .A3(new_n580), .A4(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n635), .A2(new_n666), .A3(new_n592), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n657), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n658), .A2(new_n666), .A3(new_n669), .A4(new_n592), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n582), .A2(new_n592), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT26), .B1(new_n671), .B2(new_n551), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n592), .B(KEYINPUT90), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n668), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n459), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n656), .A2(new_n676), .ZN(G369));
  NAND3_X1  g0477(.A1(new_n238), .A2(new_n281), .A3(G13), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT92), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G213), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n678), .B2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g0484(.A(KEYINPUT93), .B(G343), .Z(new_n685));
  OR3_X1    g0485(.A1(new_n684), .A2(KEYINPUT94), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT94), .B1(new_n684), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n503), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT95), .Z(new_n690));
  NAND2_X1  g0490(.A1(new_n501), .A2(new_n505), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n511), .B2(new_n690), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n688), .A2(new_n617), .ZN(new_n695));
  INV_X1    g0495(.A(new_n688), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n636), .A2(new_n695), .B1(new_n632), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n688), .B1(new_n501), .B2(new_n505), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n632), .A3(new_n635), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n632), .A2(new_n688), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n698), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n207), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n573), .A2(new_n479), .A3(new_n574), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n708), .A3(G1), .ZN(new_n709));
  INV_X1    g0509(.A(new_n212), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n706), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(new_n674), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n297), .B1(new_n546), .B2(new_n525), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n540), .B(new_n526), .C1(new_n714), .C2(KEYINPUT82), .ZN(new_n715));
  INV_X1    g0515(.A(new_n543), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n551), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n635), .A2(new_n666), .A3(new_n592), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n713), .B1(new_n719), .B2(new_n657), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n688), .B1(new_n720), .B2(new_n673), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT96), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n675), .A2(new_n696), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT96), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n671), .A2(new_n551), .A3(KEYINPUT26), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n658), .A2(new_n592), .A3(new_n666), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n727), .B1(KEYINPUT26), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n688), .B1(new_n720), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n722), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n546), .A2(new_n591), .A3(new_n628), .A4(new_n525), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(new_n477), .ZN(new_n735));
  INV_X1    g0535(.A(new_n542), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n622), .A2(new_n623), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n565), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n477), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n736), .A2(new_n738), .A3(new_n739), .A4(KEYINPUT30), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n565), .A2(new_n334), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n741), .A2(new_n498), .A3(new_n624), .A4(new_n542), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n735), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n743), .A2(new_n744), .A3(new_n688), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(new_n743), .B2(new_n688), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n512), .A2(new_n637), .A3(new_n696), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n732), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n712), .B1(new_n752), .B2(G1), .ZN(G364));
  NAND2_X1  g0553(.A1(new_n281), .A2(G13), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT97), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G45), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G1), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n705), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n694), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G330), .B2(new_n693), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n309), .A2(new_n207), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n207), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n233), .A2(new_n557), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n704), .A2(new_n309), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n212), .B2(new_n557), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n273), .B1(G20), .B2(new_n432), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n758), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n334), .A2(new_n281), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n424), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n297), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n777), .A2(G200), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n278), .A2(new_n779), .B1(new_n781), .B2(new_n280), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n281), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G87), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(new_n424), .A3(G200), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n309), .C1(new_n534), .C2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n424), .A2(G179), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n281), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n483), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n783), .A2(new_n424), .A3(new_n297), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G159), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n782), .A2(new_n788), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n776), .A2(G190), .ZN(new_n797));
  OR3_X1    g0597(.A1(new_n797), .A2(KEYINPUT99), .A3(new_n297), .ZN(new_n798));
  OAI21_X1  g0598(.A(KEYINPUT99), .B1(new_n797), .B2(new_n297), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OR3_X1    g0601(.A1(new_n797), .A2(KEYINPUT98), .A3(G200), .ZN(new_n802));
  OAI21_X1  g0602(.A(KEYINPUT98), .B1(new_n797), .B2(G200), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n796), .B1(new_n202), .B2(new_n801), .C1(new_n326), .C2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n778), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n781), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G303), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n363), .B1(new_n784), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n811), .A2(KEYINPUT100), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(KEYINPUT100), .ZN(new_n813));
  INV_X1    g0613(.A(new_n787), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n814), .A2(G283), .B1(new_n793), .B2(G329), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n620), .B2(new_n790), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n809), .A2(new_n812), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G322), .ZN(new_n818));
  INV_X1    g0618(.A(G326), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n804), .C1(new_n819), .C2(new_n801), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n805), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n775), .B1(new_n821), .B2(new_n772), .ZN(new_n822));
  INV_X1    g0622(.A(new_n771), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n693), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n760), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  OAI211_X1 g0626(.A(new_n380), .B(new_n388), .C1(new_n360), .C2(new_n696), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT102), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n360), .B1(new_n686), .B2(new_n687), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(new_n651), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n651), .A2(new_n828), .A3(new_n829), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n723), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n832), .B1(new_n827), .B2(new_n830), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n675), .A2(new_n836), .A3(new_n696), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n758), .B1(new_n838), .B2(new_n751), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n751), .B2(new_n838), .ZN(new_n840));
  INV_X1    g0640(.A(new_n758), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n772), .A2(new_n769), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n280), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n801), .A2(new_n810), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n309), .B1(new_n814), .B2(G87), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n534), .B2(new_n784), .C1(new_n808), .C2(new_n792), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n791), .B(new_n846), .C1(new_n780), .C2(G116), .ZN(new_n847));
  INV_X1    g0647(.A(G283), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n779), .ZN(new_n849));
  INV_X1    g0649(.A(new_n804), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n844), .B(new_n849), .C1(G294), .C2(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G150), .A2(new_n778), .B1(new_n780), .B2(G159), .ZN(new_n852));
  INV_X1    g0652(.A(G143), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n804), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G137), .B2(new_n800), .ZN(new_n855));
  XNOR2_X1  g0655(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n855), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n309), .B1(new_n784), .B2(new_n202), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n814), .A2(G68), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n860), .B2(new_n792), .ZN(new_n861));
  INV_X1    g0661(.A(new_n790), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n858), .B(new_n861), .C1(G58), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n851), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n772), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n843), .B1(new_n836), .B2(new_n770), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n840), .A2(new_n866), .ZN(G384));
  NOR3_X1   g0667(.A1(new_n273), .A2(new_n281), .A3(new_n479), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n536), .B(KEYINPUT103), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT35), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT36), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n280), .B(new_n710), .C1(G58), .C2(G68), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n875), .A2(KEYINPUT104), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n875), .A2(KEYINPUT104), .B1(new_n202), .B2(G68), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n238), .B(G13), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT105), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n684), .B1(new_n405), .B2(new_n409), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n449), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n449), .A2(new_n880), .A3(new_n881), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n443), .A2(new_n427), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n885), .B2(new_n881), .ZN(new_n886));
  INV_X1    g0686(.A(new_n881), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n443), .A4(new_n427), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n884), .A4(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n644), .A2(new_n431), .A3(new_n645), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n881), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n893), .A2(new_n890), .ZN(new_n894));
  XNOR2_X1  g0694(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n647), .A2(new_n457), .A3(new_n648), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n307), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n688), .A2(new_n294), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n650), .A2(new_n899), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n294), .B2(new_n649), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n834), .B1(new_n748), .B2(new_n749), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n896), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT40), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n884), .A2(new_n890), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n882), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n891), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n905), .A2(new_n909), .A3(new_n913), .A4(new_n906), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n915), .A2(new_n459), .A3(new_n750), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n459), .B2(new_n750), .ZN(new_n917));
  INV_X1    g0717(.A(G330), .ZN(new_n918));
  OR3_X1    g0718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n911), .A2(new_n910), .A3(new_n882), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n895), .B1(new_n893), .B2(new_n890), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n458), .A2(new_n696), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n912), .A2(new_n891), .A3(KEYINPUT39), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n380), .A2(new_n688), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n837), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n905), .A2(new_n913), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n684), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n646), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n927), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n722), .A2(new_n459), .A3(new_n726), .A4(new_n731), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n656), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n919), .A2(new_n937), .B1(new_n238), .B2(new_n755), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT107), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n919), .A2(new_n937), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n938), .B2(new_n939), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n879), .B1(new_n940), .B2(new_n942), .ZN(G367));
  NAND2_X1  g0743(.A1(new_n229), .A2(new_n765), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n944), .B(new_n773), .C1(new_n207), .C2(new_n354), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT109), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n758), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n945), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT110), .Z(new_n949));
  AOI22_X1  g0749(.A1(new_n785), .A2(G58), .B1(new_n814), .B2(G77), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n862), .A2(G68), .ZN(new_n951));
  XOR2_X1   g0751(.A(KEYINPUT112), .B(G137), .Z(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n363), .B1(new_n953), .B2(new_n793), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n950), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n781), .A2(new_n202), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(G159), .C2(new_n778), .ZN(new_n957));
  INV_X1    g0757(.A(G150), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n957), .B1(new_n853), .B2(new_n801), .C1(new_n958), .C2(new_n804), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n785), .A2(KEYINPUT46), .A3(G116), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT46), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n784), .B2(new_n479), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n962), .C1(new_n779), .C2(new_n620), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT111), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n808), .B2(new_n801), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n309), .B1(new_n814), .B2(G97), .ZN(new_n966));
  INV_X1    g0766(.A(G317), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n966), .B1(new_n967), .B2(new_n792), .C1(new_n573), .C2(new_n790), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G283), .B2(new_n780), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n804), .B2(new_n810), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n959), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT47), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n865), .B1(new_n971), .B2(new_n972), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n949), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n666), .A2(new_n592), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n696), .A2(new_n580), .ZN(new_n977));
  MUX2_X1   g0777(.A(new_n976), .B(new_n674), .S(new_n977), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n771), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n662), .B1(new_n540), .B2(new_n696), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n658), .A2(new_n688), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(new_n700), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n551), .B1(new_n981), .B2(new_n632), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n985), .A2(KEYINPUT42), .B1(new_n696), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(KEYINPUT42), .B2(new_n985), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT43), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n978), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n978), .A2(new_n989), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n990), .B(new_n991), .Z(new_n992));
  NOR2_X1   g0792(.A1(new_n698), .A2(new_n984), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n992), .B(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n757), .B(KEYINPUT108), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n702), .A2(new_n983), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT45), .Z(new_n999));
  NOR2_X1   g0799(.A1(new_n702), .A2(new_n983), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1002), .A2(new_n694), .A3(new_n697), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n698), .A3(new_n1001), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n700), .B1(new_n697), .B2(new_n699), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n694), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n752), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n752), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n705), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n997), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n980), .B1(new_n995), .B2(new_n1012), .ZN(G387));
  NAND2_X1  g0813(.A1(new_n862), .A2(G283), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G303), .A2(new_n780), .B1(new_n778), .B2(G311), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n804), .B2(new_n967), .C1(new_n818), .C2(new_n801), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1014), .B1(new_n620), .B2(new_n784), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT49), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n363), .B1(new_n792), .B2(new_n819), .C1(new_n479), .C2(new_n787), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1019), .B2(KEYINPUT49), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G77), .A2(new_n785), .B1(new_n793), .B2(G150), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n862), .A2(new_n584), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n363), .B1(new_n814), .B2(G97), .ZN(new_n1026));
  AND3_X1   g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n781), .B2(new_n278), .C1(new_n406), .C2(new_n779), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G159), .B2(new_n800), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n202), .B2(new_n804), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n865), .B1(new_n1023), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n323), .A2(G50), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT114), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g0834(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n708), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1033), .A2(KEYINPUT50), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n765), .B1(new_n226), .B2(new_n557), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(G107), .B2(new_n207), .C1(new_n708), .C2(new_n761), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n841), .B1(new_n1039), .B2(new_n773), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n697), .B2(new_n823), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1031), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1007), .A2(new_n997), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT113), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1007), .A2(KEYINPUT113), .A3(new_n997), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n706), .B1(new_n752), .B2(new_n1007), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n752), .B2(new_n1007), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(G393));
  NAND2_X1  g0850(.A1(new_n1005), .A2(KEYINPUT115), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT115), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1003), .A2(new_n1052), .A3(new_n1004), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n997), .A3(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n773), .B1(new_n483), .B2(new_n207), .C1(new_n236), .C2(new_n766), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n758), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT116), .Z(new_n1057));
  AOI22_X1  g0857(.A1(new_n850), .A2(G159), .B1(G150), .B2(new_n800), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT51), .Z(new_n1059));
  NOR2_X1   g0859(.A1(new_n779), .A2(new_n202), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n790), .A2(new_n280), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n309), .B1(new_n787), .B2(new_n412), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n784), .A2(new_n278), .B1(new_n792), .B2(new_n853), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1059), .B(new_n1064), .C1(new_n323), .C2(new_n781), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n801), .A2(new_n967), .B1(new_n804), .B2(new_n808), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n309), .B1(new_n814), .B2(G107), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n848), .B2(new_n784), .C1(new_n818), .C2(new_n792), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT117), .Z(new_n1070));
  NAND2_X1  g0870(.A1(new_n778), .A2(G303), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n780), .A2(G294), .B1(G116), .B2(new_n862), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1065), .A2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1057), .B1(new_n823), .B2(new_n983), .C1(new_n1074), .C2(new_n865), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n705), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1054), .B(new_n1075), .C1(new_n1076), .C2(new_n1077), .ZN(G390));
  NOR4_X1   g0878(.A1(new_n511), .A2(new_n594), .A3(new_n636), .A4(new_n688), .ZN(new_n1079));
  OAI211_X1 g0879(.A(G330), .B(new_n836), .C1(new_n1079), .C2(new_n747), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n901), .B2(new_n904), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n675), .A2(new_n836), .A3(new_n696), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n899), .B1(new_n307), .B2(new_n897), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1082), .A2(new_n928), .B1(new_n1083), .B2(new_n903), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1084), .A2(new_n924), .B1(new_n923), .B2(new_n926), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n924), .B1(new_n921), .B2(new_n922), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n730), .A2(new_n836), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n929), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1086), .B1(new_n1088), .B2(new_n905), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1081), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n906), .B(G330), .C1(new_n1083), .C2(new_n903), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n928), .B1(new_n730), .B2(new_n836), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1083), .A2(new_n903), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n924), .B(new_n896), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n923), .A2(new_n926), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n925), .B1(new_n905), .B2(new_n930), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1091), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n459), .A2(G330), .A3(new_n750), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n935), .A2(new_n1098), .A3(new_n656), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n901), .A2(new_n904), .A3(new_n1080), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n930), .B1(new_n1101), .B2(new_n1081), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1093), .A2(new_n1080), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1091), .A2(new_n1103), .A3(new_n1092), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1090), .A2(new_n1097), .A3(new_n1100), .A4(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1106), .A2(new_n705), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT119), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT118), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1090), .A2(new_n1097), .A3(KEYINPUT118), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1105), .A2(new_n1100), .ZN(new_n1113));
  AND4_X1   g0913(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1099), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1108), .B1(new_n1116), .B2(new_n1112), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1107), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n793), .A2(G294), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n786), .A2(new_n859), .A3(new_n1119), .A4(new_n363), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1061), .B(new_n1120), .C1(new_n778), .C2(new_n364), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n483), .B2(new_n781), .C1(new_n479), .C2(new_n804), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G283), .B2(new_n800), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT120), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n780), .A2(new_n1125), .B1(new_n778), .B2(new_n953), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n784), .A2(new_n958), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT53), .ZN(new_n1128));
  INV_X1    g0928(.A(G125), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n309), .B1(new_n792), .B2(new_n1129), .C1(new_n202), .C2(new_n787), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G159), .B2(new_n862), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1126), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n804), .A2(new_n860), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(G128), .C2(new_n800), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n772), .B1(new_n1123), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n841), .B1(new_n406), .B2(new_n842), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(new_n1095), .C2(new_n770), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT121), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1090), .A2(new_n1097), .A3(new_n997), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1118), .A2(new_n1141), .ZN(G378));
  NAND2_X1  g0942(.A1(new_n333), .A2(new_n932), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n351), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n351), .A2(new_n1144), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OR3_X1    g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n934), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n927), .A2(new_n931), .A3(new_n933), .A4(new_n1152), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n915), .A2(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n918), .B1(new_n908), .B2(new_n914), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n1155), .A3(new_n1154), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1153), .A2(new_n769), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n842), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n758), .B1(G50), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G50), .B1(new_n394), .B2(new_n460), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n778), .A2(G97), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G41), .B(new_n309), .C1(new_n785), .C2(G77), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n814), .A2(G58), .B1(new_n793), .B2(G283), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1166), .A2(new_n951), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n584), .B2(new_n780), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n534), .B2(new_n804), .C1(new_n479), .C2(new_n801), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT58), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1165), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n850), .A2(G128), .B1(G125), .B2(new_n800), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n778), .A2(G132), .B1(G150), .B2(new_n862), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT122), .B1(new_n1125), .B2(new_n785), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1125), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT122), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1177), .A2(new_n1178), .A3(new_n784), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1176), .B(new_n1179), .C1(G137), .C2(new_n780), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1174), .A2(new_n1175), .A3(new_n1180), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n814), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1173), .B1(new_n1172), .B2(new_n1171), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1164), .B1(new_n1189), .B2(new_n772), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1161), .A2(new_n997), .B1(new_n1162), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1106), .A2(new_n1100), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1160), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1159), .B1(new_n1155), .B2(new_n1154), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1192), .B(KEYINPUT57), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n705), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1158), .A2(new_n1160), .B1(new_n1106), .B2(new_n1100), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(KEYINPUT57), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1191), .B1(new_n1196), .B2(new_n1198), .ZN(G375));
  NAND3_X1  g0999(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1113), .A2(new_n1011), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n363), .B1(new_n787), .B2(new_n280), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n784), .A2(new_n483), .B1(new_n792), .B2(new_n810), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n584), .C2(new_n862), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n781), .B2(new_n573), .C1(new_n479), .C2(new_n779), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n804), .A2(new_n848), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(G294), .C2(new_n800), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G128), .A2(new_n793), .B1(new_n785), .B2(G159), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT124), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(KEYINPUT124), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n309), .B1(new_n787), .B2(new_n326), .C1(new_n790), .C2(new_n202), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G150), .A2(new_n780), .B1(new_n778), .B2(new_n1125), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n860), .C2(new_n801), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n850), .B2(new_n953), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n772), .B1(new_n1207), .B2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n758), .C1(G68), .C2(new_n1163), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1093), .B2(new_n769), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1105), .B2(new_n997), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1201), .A2(new_n1220), .ZN(G381));
  NAND2_X1  g1021(.A1(new_n1116), .A2(new_n1112), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT119), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1116), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1140), .B1(new_n1225), .B2(new_n1107), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1161), .A2(new_n997), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1162), .A2(new_n1190), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n706), .B1(new_n1197), .B2(KEYINPUT57), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1161), .A2(new_n1192), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT57), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1229), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1226), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(G390), .ZN(new_n1236));
  INV_X1    g1036(.A(G384), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OR4_X1    g1039(.A1(G387), .A2(new_n1235), .A3(G381), .A4(new_n1239), .ZN(G407));
  INV_X1    g1040(.A(new_n685), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(new_n682), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1235), .A2(new_n1243), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT125), .Z(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1046(.A1(new_n1197), .A2(new_n1011), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1118), .A2(new_n1141), .A3(new_n1191), .A4(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1248), .B(new_n1243), .C1(new_n1226), .C2(new_n1234), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1242), .A2(G2897), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT127), .Z(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1200), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .A4(KEYINPUT60), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(new_n705), .A3(new_n1113), .A4(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(G384), .A3(new_n1220), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G384), .B1(new_n1255), .B2(new_n1220), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1256), .B1(new_n1257), .B2(KEYINPUT126), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT126), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1259), .B(G384), .C1(new_n1255), .C2(new_n1220), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1251), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1220), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1237), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1259), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1251), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1256), .A4(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1261), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1249), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G378), .A2(G375), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(new_n1243), .A3(new_n1248), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1191), .A2(new_n1247), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1242), .B1(new_n1226), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1269), .A2(new_n1273), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1238), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G390), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n992), .B(new_n993), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1012), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1283), .A2(new_n1284), .B1(new_n979), .B2(new_n975), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1279), .A2(G390), .A3(new_n1280), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1282), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1285), .B1(new_n1282), .B2(new_n1286), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1278), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1272), .A2(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1275), .A2(KEYINPUT63), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1269), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(G405));
  NAND2_X1  g1096(.A1(new_n1235), .A2(new_n1270), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1271), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1235), .B(new_n1270), .C1(new_n1260), .C2(new_n1258), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1300), .B(new_n1291), .ZN(G402));
endmodule


