//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n187));
  OAI21_X1  g001(.A(G214), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  OAI21_X1  g003(.A(G210), .B1(G237), .B2(G902), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G122), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT68), .A2(G119), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT68), .A2(G119), .ZN(new_n195));
  OAI21_X1  g009(.A(G116), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT67), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT2), .B(G113), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(KEYINPUT67), .A3(new_n201), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G107), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT77), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n206), .A2(new_n209), .A3(new_n211), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G101), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(G101), .A3(new_n214), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n203), .A2(new_n204), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n208), .A2(KEYINPUT78), .A3(G104), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n208), .B2(G104), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n205), .A2(G107), .ZN(new_n224));
  OAI211_X1 g038(.A(G101), .B(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n212), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n196), .A2(KEYINPUT5), .A3(new_n198), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT68), .B(G119), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G116), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(G113), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n202), .A2(new_n196), .A3(new_n198), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n193), .B1(new_n220), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n203), .A2(new_n204), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n218), .A2(new_n219), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n192), .A3(new_n234), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n240), .A3(KEYINPUT6), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(G146), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT64), .A3(G143), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n249), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G125), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT1), .B1(new_n243), .B2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G128), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n248), .A2(new_n259), .B1(new_n253), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G224), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT80), .ZN(new_n266));
  OR3_X1    g080(.A1(new_n257), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n257), .B2(new_n263), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n270), .B(new_n193), .C1(new_n220), .C2(new_n235), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n241), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G902), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT82), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT81), .B(KEYINPUT8), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n192), .B(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n227), .B1(new_n232), .B2(new_n233), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n275), .B(new_n277), .C1(new_n235), .C2(new_n278), .ZN(new_n279));
  OR3_X1    g093(.A1(new_n257), .A2(new_n263), .A3(KEYINPUT7), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT7), .B(new_n266), .C1(new_n257), .C2(new_n263), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n232), .A2(new_n233), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n226), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n234), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n275), .B1(new_n285), .B2(new_n277), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n220), .A2(new_n235), .A3(new_n193), .ZN(new_n287));
  INV_X1    g101(.A(new_n267), .ZN(new_n288));
  NOR4_X1   g102(.A1(new_n282), .A2(new_n286), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n191), .B1(new_n274), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n282), .ZN(new_n291));
  INV_X1    g105(.A(new_n286), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n291), .A2(new_n267), .A3(new_n240), .A4(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n293), .A2(new_n273), .A3(new_n190), .A4(new_n272), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n189), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(G234), .A2(G237), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(G952), .A3(new_n264), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT21), .B(G898), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(KEYINPUT90), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(G902), .A3(G953), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G469), .ZN(new_n302));
  XNOR2_X1  g116(.A(G110), .B(G140), .ZN(new_n303));
  INV_X1    g117(.A(G227), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(G953), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n303), .B(new_n305), .Z(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n246), .A2(G143), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n261), .A2(new_n308), .A3(new_n245), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n260), .B1(new_n308), .B2(KEYINPUT1), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(new_n253), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n212), .A3(new_n225), .ZN(new_n312));
  INV_X1    g126(.A(new_n262), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n312), .B1(new_n313), .B2(new_n227), .ZN(new_n314));
  INV_X1    g128(.A(G134), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT65), .B1(new_n315), .B2(G137), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT11), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(G137), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT11), .ZN(new_n319));
  OAI211_X1 g133(.A(KEYINPUT65), .B(new_n319), .C1(new_n315), .C2(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G131), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n317), .A2(new_n323), .A3(new_n318), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n314), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n314), .A2(KEYINPUT12), .A3(new_n325), .ZN(new_n329));
  INV_X1    g143(.A(new_n255), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n238), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT10), .B1(new_n262), .B2(new_n226), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT10), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n311), .A2(new_n333), .A3(new_n212), .A4(new_n225), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n325), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n331), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT79), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n331), .A2(new_n335), .A3(new_n339), .A4(new_n336), .ZN(new_n340));
  AOI221_X4 g154(.A(new_n307), .B1(new_n328), .B2(new_n329), .C1(new_n338), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n340), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n331), .A2(new_n335), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n325), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n306), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n302), .B(new_n273), .C1(new_n341), .C2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n344), .A3(new_n306), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n338), .A2(new_n340), .B1(new_n329), .B2(new_n328), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n347), .B(G469), .C1(new_n306), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(G469), .A2(G902), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G221), .ZN(new_n352));
  XOR2_X1   g166(.A(KEYINPUT9), .B(G234), .Z(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n353), .B2(new_n273), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n295), .A2(new_n301), .A3(new_n351), .A4(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G475), .ZN(new_n357));
  XNOR2_X1  g171(.A(G113), .B(G122), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(new_n205), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(KEYINPUT69), .A2(G237), .ZN(new_n361));
  NOR2_X1   g175(.A1(KEYINPUT69), .A2(G237), .ZN(new_n362));
  OAI211_X1 g176(.A(G214), .B(new_n264), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  XOR2_X1   g177(.A(KEYINPUT83), .B(G143), .Z(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT69), .B(G237), .ZN(new_n366));
  NOR2_X1   g180(.A1(KEYINPUT83), .A2(G143), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n366), .A2(G214), .A3(new_n264), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n323), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n368), .A3(G131), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(KEYINPUT85), .A3(new_n323), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT17), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT17), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n256), .A2(KEYINPUT16), .A3(G140), .ZN(new_n378));
  XNOR2_X1  g192(.A(G125), .B(G140), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(KEYINPUT16), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G146), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT16), .ZN(new_n382));
  OR2_X1    g196(.A1(G125), .A2(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(G125), .A2(G140), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n246), .B1(new_n385), .B2(new_n378), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT86), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n381), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n375), .A2(new_n377), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n372), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT18), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n379), .B(KEYINPUT84), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G146), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n379), .A2(KEYINPUT73), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n383), .A2(new_n398), .A3(new_n384), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n246), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n369), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n394), .A2(new_n402), .A3(new_n404), .A4(new_n370), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n360), .B1(new_n392), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n372), .A2(new_n371), .ZN(new_n408));
  AOI21_X1  g222(.A(G131), .B1(new_n365), .B2(new_n368), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n374), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n376), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n377), .ZN(new_n413));
  INV_X1    g227(.A(new_n391), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n359), .A3(new_n405), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n407), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n357), .B1(new_n417), .B2(new_n273), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT19), .B1(new_n397), .B2(new_n399), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(KEYINPUT19), .B2(new_n395), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n246), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n421), .A2(new_n374), .A3(new_n373), .A4(new_n381), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n359), .B1(new_n422), .B2(new_n405), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(G475), .A2(G902), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT20), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n428));
  INV_X1    g242(.A(new_n426), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n428), .B(new_n429), .C1(new_n416), .C2(new_n424), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n418), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G122), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G116), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(G116), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT14), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n197), .A2(G122), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT88), .B1(new_n439), .B2(KEYINPUT14), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n438), .B(G107), .C1(new_n436), .C2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G128), .B(G143), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(new_n315), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n433), .A2(new_n439), .A3(new_n208), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(KEYINPUT13), .ZN(new_n446));
  OR3_X1    g260(.A1(new_n260), .A2(KEYINPUT13), .A3(G143), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(G134), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT87), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n433), .A2(new_n439), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G107), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n451), .A2(new_n444), .B1(new_n315), .B2(new_n442), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n446), .A2(new_n453), .A3(G134), .A4(new_n447), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n445), .B2(new_n455), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n353), .A2(G217), .A3(new_n264), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n460), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n445), .A2(new_n455), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT89), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n464), .B2(new_n457), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n273), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G478), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(KEYINPUT15), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n460), .B1(new_n458), .B2(new_n459), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n464), .A2(new_n462), .A3(new_n457), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n472), .B(new_n273), .C1(KEYINPUT15), .C2(new_n467), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n431), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n187), .B1(new_n356), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n415), .A2(new_n359), .A3(new_n405), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n359), .B1(new_n415), .B2(new_n405), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n273), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G475), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n373), .A2(new_n374), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n377), .B1(new_n482), .B2(new_n376), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n406), .B1(new_n483), .B2(new_n414), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n423), .B1(new_n484), .B2(new_n359), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n428), .B1(new_n485), .B2(new_n429), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n425), .A2(KEYINPUT20), .A3(new_n426), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n481), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(new_n474), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n351), .A2(new_n355), .ZN(new_n490));
  INV_X1    g304(.A(new_n301), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n491), .B(new_n189), .C1(new_n290), .C2(new_n294), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT91), .A4(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT22), .ZN(new_n496));
  INV_X1    g310(.A(G137), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT22), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n495), .B(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(G137), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n494), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(G137), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n496), .A2(new_n497), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT74), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n401), .A2(new_n381), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n229), .A2(G128), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n260), .A2(G119), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(KEYINPUT23), .A3(new_n509), .ZN(new_n510));
  OR4_X1    g324(.A1(KEYINPUT23), .A2(new_n194), .A3(new_n195), .A4(G128), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G110), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n508), .A2(new_n509), .ZN(new_n515));
  XOR2_X1   g329(.A(KEYINPUT24), .B(G110), .Z(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n507), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n508), .A2(new_n509), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n516), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n510), .A2(new_n511), .A3(G110), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n521), .A2(new_n522), .A3(new_n387), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n506), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n518), .ZN(new_n525));
  AOI21_X1  g339(.A(G110), .B1(new_n510), .B2(new_n511), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n401), .B(new_n381), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n498), .A2(new_n501), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n521), .A2(new_n522), .A3(new_n387), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n524), .A2(new_n273), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT75), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT25), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G234), .ZN(new_n536));
  OAI21_X1  g350(.A(G217), .B1(new_n536), .B2(G902), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT25), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n273), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT76), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n524), .A3(new_n530), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G472), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  INV_X1    g362(.A(new_n237), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n255), .B1(new_n322), .B2(new_n324), .ZN(new_n550));
  INV_X1    g364(.A(new_n324), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n497), .A2(KEYINPUT66), .A3(G134), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT66), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n497), .B2(G134), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n315), .A2(G137), .ZN(new_n555));
  OAI211_X1 g369(.A(G131), .B(new_n552), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n551), .A2(new_n262), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT71), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n550), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n325), .A2(new_n330), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n313), .A2(new_n324), .A3(new_n556), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT71), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n548), .B(new_n549), .C1(new_n560), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n366), .A2(G210), .A3(new_n264), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT26), .B(G101), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n549), .A2(new_n561), .A3(new_n562), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n237), .B1(new_n550), .B2(new_n558), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(KEYINPUT28), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n564), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT30), .B1(new_n550), .B2(new_n558), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT30), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n561), .A2(new_n575), .A3(new_n562), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n549), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n570), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n577), .A2(new_n578), .A3(new_n569), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT31), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n573), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n550), .A2(new_n558), .A3(KEYINPUT30), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n575), .B1(new_n561), .B2(new_n562), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n237), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n569), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n570), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(KEYINPUT31), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n547), .B(new_n273), .C1(new_n581), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT32), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n579), .A2(new_n580), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(KEYINPUT31), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n573), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT32), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n547), .A4(new_n273), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n564), .ZN(new_n596));
  INV_X1    g410(.A(new_n572), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n585), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT29), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(KEYINPUT29), .B(new_n585), .C1(new_n596), .C2(new_n597), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n273), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G472), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n546), .B1(new_n595), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n477), .A2(new_n493), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT92), .B(G101), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  OAI21_X1  g422(.A(new_n273), .B1(new_n581), .B2(new_n587), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G472), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n588), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n356), .A2(new_n546), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n472), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT33), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n614), .A2(G478), .A3(new_n273), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n466), .A2(new_n467), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n488), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND4_X1  g437(.A1(new_n481), .A2(new_n474), .A3(new_n486), .A4(new_n487), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n612), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  INV_X1    g442(.A(new_n611), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT93), .B1(new_n519), .B2(new_n523), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT93), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n527), .A2(new_n631), .A3(new_n529), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n506), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT36), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n633), .A2(new_n636), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n544), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n540), .A2(new_n639), .A3(KEYINPUT94), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT94), .B1(new_n540), .B2(new_n639), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n477), .A2(new_n493), .A3(new_n629), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT37), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n513), .ZN(G12));
  AOI22_X1  g459(.A1(new_n589), .A2(new_n594), .B1(new_n603), .B2(G472), .ZN(new_n646));
  INV_X1    g460(.A(new_n295), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n351), .A2(new_n355), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT96), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n297), .B(KEYINPUT95), .Z(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n652), .B1(G900), .B2(new_n300), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n431), .A2(new_n650), .A3(new_n474), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n653), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT96), .B1(new_n624), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n649), .A2(new_n657), .A3(new_n642), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  NAND2_X1  g473(.A1(new_n570), .A2(new_n571), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n569), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n661), .A2(KEYINPUT97), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(KEYINPUT97), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n586), .A3(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n664), .A2(new_n273), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n595), .B1(new_n547), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT98), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n290), .A2(new_n294), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT38), .Z(new_n669));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n653), .B(KEYINPUT39), .Z(new_n672));
  NOR2_X1   g486(.A1(new_n648), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n189), .B1(new_n674), .B2(KEYINPUT40), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT94), .ZN(new_n676));
  INV_X1    g490(.A(new_n539), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT25), .B1(new_n531), .B2(new_n532), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n677), .A2(new_n678), .A3(new_n541), .ZN(new_n679));
  INV_X1    g493(.A(new_n638), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n633), .A2(new_n636), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n543), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n676), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n540), .A2(new_n639), .A3(KEYINPUT94), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n427), .A2(new_n430), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n475), .B1(new_n686), .B2(new_n481), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n673), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n675), .A2(new_n685), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n671), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  NOR2_X1   g506(.A1(new_n619), .A2(new_n655), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n649), .A2(new_n642), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NOR2_X1   g509(.A1(new_n341), .A2(new_n345), .ZN(new_n696));
  OAI21_X1  g510(.A(G469), .B1(new_n696), .B2(G902), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n355), .A3(new_n346), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n605), .A2(new_n492), .A3(new_n620), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n605), .A2(new_n492), .A3(new_n625), .A4(new_n699), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  NOR2_X1   g518(.A1(new_n476), .A2(new_n491), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n595), .A2(new_n604), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n647), .A2(new_n698), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n705), .A2(new_n706), .A3(new_n642), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  INV_X1    g523(.A(KEYINPUT99), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n573), .B(new_n710), .C1(new_n579), .C2(new_n580), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n590), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n710), .B1(new_n591), .B2(new_n573), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n547), .B(new_n273), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n610), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n546), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n698), .A2(new_n491), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n488), .A2(new_n295), .A3(new_n474), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(KEYINPUT100), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT100), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n687), .B2(new_n295), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n716), .B(new_n717), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT101), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n715), .B2(new_n685), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n642), .A2(KEYINPUT102), .A3(new_n610), .A4(new_n714), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n693), .A3(new_n707), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n731));
  INV_X1    g545(.A(new_n546), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n706), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n350), .B(KEYINPUT103), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n346), .A2(new_n349), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT104), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n346), .A2(new_n349), .A3(new_n737), .A4(new_n734), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n355), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT105), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n736), .A2(new_n741), .A3(new_n355), .A4(new_n738), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n733), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n619), .A2(new_n189), .A3(new_n668), .A4(new_n655), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT42), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n740), .A2(new_n742), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(KEYINPUT42), .A3(new_n605), .A4(new_n744), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n731), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n605), .A3(new_n744), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT106), .A3(new_n747), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  NOR2_X1   g569(.A1(new_n668), .A2(new_n189), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n743), .A2(new_n657), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n347), .B1(new_n348), .B2(new_n306), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(G469), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT107), .Z(new_n763));
  INV_X1    g577(.A(new_n734), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n346), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n763), .A2(new_n759), .A3(new_n764), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n355), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(new_n672), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n488), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(KEYINPUT43), .A3(new_n618), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n431), .A2(new_n618), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n685), .B1(new_n778), .B2(KEYINPUT110), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n772), .B(new_n773), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n776), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n779), .A2(new_n611), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n769), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n756), .C1(new_n786), .C2(new_n785), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n768), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT47), .B(new_n355), .C1(new_n766), .C2(new_n767), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n744), .A2(new_n546), .A3(new_n646), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT111), .Z(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  AND2_X1   g611(.A1(new_n667), .A2(new_n355), .ZN(new_n798));
  INV_X1    g612(.A(new_n697), .ZN(new_n799));
  INV_X1    g613(.A(new_n346), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT49), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n188), .A2(new_n802), .A3(new_n669), .A4(new_n771), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n798), .A2(new_n732), .A3(new_n618), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n782), .A2(new_n651), .A3(new_n699), .A4(new_n716), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n669), .A2(new_n189), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n716), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n778), .A2(new_n652), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n808), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(KEYINPUT50), .A3(new_n699), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n728), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n699), .A2(new_n756), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n778), .A2(new_n652), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n297), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n816), .A2(new_n546), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n667), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n488), .A3(new_n618), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n814), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT119), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n814), .A2(new_n826), .A3(new_n818), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n801), .A2(new_n354), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n791), .A2(new_n792), .A3(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n830), .A2(new_n756), .A3(new_n811), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n805), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n778), .A2(new_n733), .A3(new_n652), .A4(new_n816), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT48), .Z(new_n834));
  OAI211_X1 g648(.A(G952), .B(new_n264), .C1(new_n821), .C2(new_n619), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n811), .B2(new_n707), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n834), .A2(KEYINPUT122), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n817), .B(new_n822), .C1(new_n809), .C2(new_n813), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n805), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n831), .B1(new_n824), .B2(KEYINPUT120), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n844), .A2(KEYINPUT121), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT121), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n832), .B(new_n841), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n752), .A2(KEYINPUT106), .A3(new_n747), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT106), .B1(new_n752), .B2(new_n747), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n728), .A2(new_n746), .A3(new_n693), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n746), .A2(new_n605), .A3(new_n657), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n476), .A2(new_n685), .A3(new_n655), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n490), .A3(new_n706), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n756), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n722), .A2(new_n703), .A3(new_n708), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n624), .B(KEYINPUT113), .Z(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n612), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n700), .ZN(new_n863));
  INV_X1    g677(.A(new_n643), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n860), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n606), .A2(new_n621), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n606), .A2(new_n621), .A3(KEYINPUT112), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n859), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n850), .B1(new_n853), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n642), .B(new_n649), .C1(new_n657), .C2(new_n693), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n718), .A2(KEYINPUT100), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n687), .A2(new_n720), .A3(new_n295), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n739), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n679), .A2(new_n682), .A3(new_n655), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n666), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n729), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT115), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n729), .A2(new_n873), .A3(new_n879), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT52), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n886), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n722), .A2(new_n703), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n295), .A2(new_n301), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n646), .A2(new_n890), .A3(new_n546), .A4(new_n698), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n891), .A2(new_n620), .B1(new_n861), .B2(new_n612), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n889), .A2(new_n643), .A3(new_n708), .A4(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n606), .A2(new_n621), .A3(KEYINPUT112), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT112), .B1(new_n606), .B2(new_n621), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n754), .A2(new_n897), .A3(KEYINPUT114), .A4(new_n859), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n872), .A2(new_n888), .A3(new_n898), .A4(KEYINPUT53), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n729), .A2(new_n873), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(KEYINPUT52), .A3(new_n879), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n887), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n872), .A2(new_n898), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT53), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n849), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n752), .A2(new_n747), .ZN(new_n910));
  AND4_X1   g724(.A1(new_n910), .A2(new_n859), .A3(new_n865), .A4(new_n870), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n905), .A3(KEYINPUT53), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT117), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n911), .A2(new_n905), .A3(new_n914), .A4(KEYINPUT53), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n872), .A2(new_n888), .A3(new_n898), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n907), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n916), .A2(new_n849), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT118), .B1(new_n909), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n901), .A2(new_n908), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT54), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n923));
  INV_X1    g737(.A(new_n919), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n848), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(G952), .A2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n804), .B1(new_n926), .B2(new_n927), .ZN(G75));
  AOI21_X1  g742(.A(new_n273), .B1(new_n916), .B2(new_n918), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT56), .B1(new_n929), .B2(G210), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n241), .A2(new_n271), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n269), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n930), .A2(new_n933), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n264), .A2(G952), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G51));
  NAND2_X1  g751(.A1(new_n734), .A2(KEYINPUT57), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n734), .A2(KEYINPUT57), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n849), .B1(new_n916), .B2(new_n918), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n938), .B(new_n939), .C1(new_n919), .C2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n696), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n941), .A2(KEYINPUT123), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT123), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n929), .A2(new_n763), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n936), .B1(new_n945), .B2(new_n946), .ZN(G54));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT58), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n357), .ZN(new_n950));
  NAND3_X1  g764(.A1(KEYINPUT124), .A2(KEYINPUT58), .A3(G475), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n929), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(new_n485), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n936), .B1(new_n952), .B2(new_n485), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(G60));
  INV_X1    g771(.A(new_n936), .ZN(new_n958));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT59), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n919), .B2(new_n940), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n614), .A2(new_n615), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n925), .A2(new_n920), .A3(new_n960), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n962), .ZN(G63));
  AND2_X1   g779(.A1(new_n916), .A2(new_n918), .ZN(new_n966));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT60), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n638), .B2(new_n637), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n524), .A2(new_n530), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n966), .B2(new_n968), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n970), .A2(new_n958), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G66));
  AOI21_X1  g789(.A(new_n264), .B1(new_n299), .B2(G224), .ZN(new_n976));
  INV_X1    g790(.A(new_n897), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(new_n264), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n931), .B1(G898), .B2(new_n264), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n978), .B(new_n979), .Z(G69));
  NOR2_X1   g794(.A1(new_n582), .A2(new_n583), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(new_n420), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n691), .A2(new_n903), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT62), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n605), .B1(new_n861), .B2(new_n620), .ZN(new_n986));
  NOR4_X1   g800(.A1(new_n986), .A2(new_n189), .A3(new_n668), .A4(new_n674), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n788), .A3(new_n796), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n983), .B1(new_n990), .B2(G953), .ZN(new_n991));
  INV_X1    g805(.A(new_n769), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n605), .A3(new_n876), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n788), .A2(new_n796), .A3(new_n903), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n754), .A2(new_n757), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n994), .A2(G953), .A3(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(G900), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n982), .B1(new_n997), .B2(new_n264), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n991), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n304), .B2(new_n997), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT126), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n991), .B(new_n1001), .C1(new_n996), .C2(new_n998), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(G72));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n989), .B2(new_n977), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n584), .A2(new_n570), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT127), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1010), .A2(new_n569), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n936), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n994), .A2(new_n977), .A3(new_n995), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1007), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n569), .B(new_n1010), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g830(.A1(new_n901), .A2(new_n908), .B1(new_n586), .B2(new_n600), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1016), .B1(new_n1007), .B2(new_n1017), .ZN(G57));
endmodule


