//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1175, new_n1176, new_n1177;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  INV_X1    g014(.A(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g027(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n453));
  NAND3_X1  g028(.A1(new_n437), .A2(new_n438), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OAI22_X1  g037(.A1(new_n461), .A2(KEYINPUT67), .B1(new_n462), .B2(new_n457), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(KEYINPUT67), .B2(new_n461), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT68), .ZN(G319));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(new_n467), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n478), .A2(KEYINPUT69), .A3(G137), .A4(new_n471), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT70), .Z(G160));
  NAND2_X1  g057(.A1(new_n478), .A2(new_n471), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n471), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT71), .B1(new_n475), .B2(new_n471), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n478), .A2(new_n489), .A3(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n487), .B1(G124), .B2(new_n491), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  AND2_X1   g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n466), .B2(new_n467), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(KEYINPUT72), .B(new_n496), .C1(new_n466), .C2(new_n467), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n471), .C1(new_n466), .C2(new_n467), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n478), .A2(new_n504), .A3(G138), .A4(new_n471), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G166));
  INV_X1    g096(.A(new_n511), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n515), .A2(G89), .ZN(new_n523));
  NAND2_X1  g098(.A1(G63), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n518), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n525), .A2(new_n529), .ZN(G168));
  AOI22_X1  g105(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n513), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G90), .Z(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n516), .A2(new_n533), .B1(new_n518), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n513), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT74), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n516), .A2(new_n540), .B1(new_n518), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT75), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G860), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  INV_X1    g128(.A(G78), .ZN(new_n554));
  INV_X1    g129(.A(G543), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n522), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT79), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n558));
  OAI221_X1 g133(.A(new_n558), .B1(new_n554), .B2(new_n555), .C1(new_n522), .C2(new_n553), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(G651), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n518), .B2(new_n562), .ZN(new_n563));
  OR2_X1    g138(.A1(KEYINPUT6), .A2(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(KEYINPUT6), .A2(G651), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n555), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n566), .A2(new_n561), .A3(new_n567), .A4(G53), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n511), .A2(new_n515), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n563), .A2(new_n568), .B1(G91), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n560), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  AOI22_X1  g148(.A1(new_n569), .A2(G88), .B1(G50), .B2(new_n566), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n574), .B(new_n575), .C1(new_n513), .C2(new_n512), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT80), .B1(new_n514), .B2(new_n520), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(G303));
  AND3_X1   g153(.A1(new_n511), .A2(new_n515), .A3(G87), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n566), .A2(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  INV_X1    g159(.A(G48), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n516), .A2(new_n584), .B1(new_n518), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n511), .A2(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n513), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n513), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n516), .A2(new_n594), .B1(new_n518), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(G171), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT81), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n511), .A2(new_n515), .A3(G92), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT82), .Z(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n602), .B(KEYINPUT82), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n522), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G54), .B2(new_n566), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n605), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n601), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n601), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  XNOR2_X1  g192(.A(G280), .B(KEYINPUT83), .ZN(G297));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n544), .A2(new_n599), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n612), .A2(new_n619), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n621), .B1(new_n623), .B2(new_n599), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n478), .A2(new_n472), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT84), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n491), .A2(G123), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(G111), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(new_n483), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n629), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(G2096), .ZN(new_n640));
  NAND4_X1  g215(.A1(new_n630), .A2(new_n638), .A3(new_n639), .A4(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT88), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT87), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2430), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n645), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT86), .ZN(new_n655));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT89), .Z(G401));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT90), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n665), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT17), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT91), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n666), .B2(new_n670), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT92), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n673), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT93), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT20), .Z(new_n688));
  NOR2_X1   g263(.A1(new_n681), .A2(new_n683), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n690), .A2(new_n686), .A3(new_n684), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n688), .B(new_n691), .C1(new_n686), .C2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  NAND2_X1  g274(.A1(G160), .A2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT94), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(KEYINPUT94), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT24), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(G34), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(G34), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT99), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(G2084), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(G2084), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n701), .A2(G32), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT26), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n472), .A2(G105), .ZN(new_n717));
  INV_X1    g292(.A(G141), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n716), .B(new_n717), .C1(new_n483), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G129), .B2(new_n491), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(new_n701), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT27), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1996), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NOR2_X1   g299(.A1(G168), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n724), .B2(G21), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n635), .A2(G139), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT25), .Z(new_n730));
  AOI22_X1  g305(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n730), .C1(new_n471), .C2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G33), .B(new_n732), .S(G29), .Z(new_n733));
  AOI22_X1  g308(.A1(new_n727), .A2(G1966), .B1(G2072), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n726), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n631), .A2(new_n636), .A3(new_n704), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT30), .B(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  NAND2_X1  g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n738), .A2(new_n701), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n734), .A2(new_n736), .A3(new_n737), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G171), .A2(new_n724), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G5), .B2(new_n724), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G2072), .B2(new_n733), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n704), .A2(G27), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n704), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT100), .B(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n744), .A2(new_n745), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n742), .A2(new_n747), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n712), .A2(new_n713), .A3(new_n723), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT101), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n705), .A2(G25), .ZN(new_n757));
  INV_X1    g332(.A(G131), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n471), .A2(G107), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n760));
  OAI22_X1  g335(.A1(new_n483), .A2(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G119), .B2(new_n491), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n757), .B1(new_n763), .B2(new_n705), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT35), .B(G1991), .Z(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n724), .A2(G24), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n597), .B2(new_n724), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1986), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G23), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT97), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n581), .A2(new_n582), .ZN(new_n775));
  OAI21_X1  g350(.A(KEYINPUT98), .B1(new_n775), .B2(new_n579), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT98), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n580), .A2(new_n777), .A3(new_n581), .A4(new_n582), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(new_n724), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n724), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n724), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n724), .A2(G6), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n590), .B2(new_n724), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT32), .B(G1981), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n780), .A2(new_n781), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n782), .A2(new_n786), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n772), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT36), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n755), .A2(KEYINPUT101), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n705), .A2(G26), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT28), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n491), .A2(G128), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G116), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n635), .B2(G140), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(G29), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2067), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n539), .A2(new_n543), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(new_n724), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n724), .B2(G19), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n808), .B1(new_n812), .B2(G1341), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n704), .A2(G35), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G162), .B2(new_n704), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT29), .Z(new_n816));
  INV_X1    g391(.A(G2090), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n724), .A2(G20), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT23), .Z(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G299), .B2(G16), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1956), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n816), .A2(new_n817), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n818), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n724), .A2(G4), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n612), .B2(new_n724), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1348), .ZN(new_n827));
  INV_X1    g402(.A(G1341), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n811), .A2(new_n828), .ZN(new_n829));
  NOR4_X1   g404(.A1(new_n813), .A2(new_n824), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n756), .A2(new_n797), .A3(new_n798), .A4(new_n830), .ZN(G150));
  INV_X1    g406(.A(G150), .ZN(G311));
  AOI22_X1  g407(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n513), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n516), .A2(new_n835), .B1(new_n518), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(new_n545), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n605), .A2(new_n607), .A3(new_n611), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n619), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT102), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n809), .A2(new_n838), .ZN(new_n845));
  INV_X1    g420(.A(new_n838), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n544), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n844), .B(new_n848), .Z(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n849), .A2(KEYINPUT103), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT103), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n545), .B1(new_n849), .B2(new_n850), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n840), .B1(new_n853), .B2(new_n854), .ZN(G145));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n732), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT104), .Z(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G142), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n471), .A2(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n483), .A2(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G130), .B2(new_n491), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n627), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n762), .ZN(new_n866));
  INV_X1    g441(.A(new_n806), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n720), .B(new_n507), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n866), .B(new_n806), .ZN(new_n871));
  INV_X1    g446(.A(new_n869), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n859), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n868), .A2(new_n869), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n858), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n878));
  XNOR2_X1  g453(.A(G160), .B(new_n637), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(G162), .Z(new_n880));
  NAND4_X1  g455(.A1(new_n874), .A2(new_n877), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n877), .A2(new_n878), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n884), .A2(new_n874), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n883), .B(KEYINPUT40), .C1(new_n885), .C2(new_n880), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n880), .B1(new_n884), .B2(new_n874), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n881), .A2(new_n882), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n886), .A2(new_n890), .ZN(G395));
  NOR2_X1   g466(.A1(new_n838), .A2(G868), .ZN(new_n892));
  XNOR2_X1  g467(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n612), .A2(new_n616), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n841), .A2(G299), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n899), .A3(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n848), .B(new_n622), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n896), .A2(new_n897), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n894), .A2(new_n895), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G305), .B(G166), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n779), .A2(G290), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n597), .A2(new_n776), .A3(new_n778), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT109), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT110), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(KEYINPUT42), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT42), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n904), .A2(new_n907), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  INV_X1    g493(.A(new_n902), .ZN(new_n919));
  INV_X1    g494(.A(new_n905), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n920), .A2(new_n899), .B1(new_n896), .B2(new_n897), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n896), .A2(new_n897), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n912), .A2(KEYINPUT42), .A3(new_n914), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n918), .A2(new_n923), .A3(new_n924), .A4(new_n906), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n917), .A2(new_n925), .A3(G868), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n892), .B1(new_n926), .B2(KEYINPUT111), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n917), .A2(new_n925), .A3(new_n928), .A4(G868), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n927), .A2(KEYINPUT112), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT112), .B1(new_n927), .B2(new_n929), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(G295));
  NAND2_X1  g507(.A1(new_n927), .A2(new_n929), .ZN(G331));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  NOR2_X1   g509(.A1(G171), .A2(KEYINPUT113), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n845), .A2(new_n847), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G286), .B1(G171), .B2(KEYINPUT113), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n936), .B1(new_n845), .B2(new_n847), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n848), .A2(new_n935), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n939), .B1(new_n943), .B2(new_n937), .ZN(new_n944));
  OAI22_X1  g519(.A1(new_n901), .A2(new_n903), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n912), .A2(new_n914), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n938), .B2(new_n941), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n939), .A3(new_n937), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n920), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n921), .A2(new_n922), .B1(new_n947), .B2(new_n948), .ZN(new_n954));
  INV_X1    g529(.A(new_n949), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n946), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n945), .A2(KEYINPUT114), .A3(new_n949), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n952), .A2(new_n959), .A3(new_n882), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n905), .A2(new_n899), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n905), .B2(new_n893), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n948), .B2(new_n947), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n957), .B1(new_n963), .B2(new_n955), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n882), .A3(new_n950), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n934), .B1(new_n960), .B2(new_n966), .ZN(new_n967));
  AND4_X1   g542(.A1(new_n951), .A2(new_n964), .A3(new_n882), .A4(new_n950), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n882), .A3(new_n950), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(KEYINPUT43), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n967), .B1(new_n934), .B2(new_n970), .ZN(G397));
  INV_X1    g546(.A(KEYINPUT63), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n507), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n501), .B2(new_n506), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n473), .A2(G40), .A3(new_n480), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n785), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n473), .A2(G40), .A3(new_n480), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(G2090), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n576), .A2(G8), .A3(new_n577), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT55), .Z(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n989), .A3(G8), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n979), .A2(new_n977), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n776), .A2(new_n778), .A3(G1976), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(G8), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT52), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n979), .B2(new_n977), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n992), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  OAI21_X1  g576(.A(G1981), .B1(new_n586), .B2(new_n589), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n586), .A2(new_n589), .A3(G1981), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1981), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n590), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(new_n1002), .A3(KEYINPUT49), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n996), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1005), .A2(new_n1008), .A3(KEYINPUT118), .A4(new_n996), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1000), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n975), .A2(G1384), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n507), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1015), .B(new_n979), .C1(KEYINPUT45), .C2(new_n977), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n735), .ZN(new_n1017));
  INV_X1    g592(.A(G2084), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n984), .A2(new_n985), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G8), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G286), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n988), .B(KEYINPUT55), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n979), .B1(new_n977), .B2(new_n983), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1026), .A2(new_n817), .B1(new_n980), .B2(new_n785), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1023), .B1(new_n1027), .B2(new_n995), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n990), .A2(new_n1013), .A3(new_n1022), .A4(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1013), .A2(new_n990), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1020), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n987), .A2(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(new_n1023), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n972), .A2(new_n1029), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1013), .A2(G8), .A3(new_n989), .A4(new_n987), .ZN(new_n1035));
  OR2_X1    g610(.A1(G288), .A2(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT119), .B1(new_n1037), .B2(new_n1004), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n996), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1037), .A2(KEYINPUT119), .A3(new_n1004), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n980), .A2(G2078), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n1044));
  AOI21_X1  g619(.A(G171), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT125), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1961), .B1(new_n984), .B2(new_n985), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n974), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1014), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n501), .B2(new_n506), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n982), .ZN(new_n1052));
  INV_X1    g627(.A(G2078), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1044), .B1(new_n1054), .B2(KEYINPUT124), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT124), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1049), .A2(new_n1052), .A3(new_n1056), .A4(new_n1053), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n1046), .B(new_n1047), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT124), .B1(new_n1016), .B2(G2078), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(KEYINPUT53), .A3(new_n1057), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1047), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT125), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1045), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1064));
  OR3_X1    g639(.A1(new_n980), .A2(new_n1044), .A3(G2078), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G171), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(KEYINPUT54), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1013), .A2(new_n990), .A3(new_n1028), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1021), .B(new_n1070), .C1(new_n995), .C2(G168), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1017), .A2(KEYINPUT123), .A3(new_n1019), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT123), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1072), .A2(new_n1073), .A3(G286), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1070), .A2(new_n995), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1071), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(G168), .A2(new_n995), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1069), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1045), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1064), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(G171), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1068), .B(new_n1080), .C1(new_n1083), .C2(KEYINPUT54), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n1085));
  XNOR2_X1  g660(.A(G299), .B(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1956), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT56), .B(G2072), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n976), .A2(new_n978), .A3(new_n979), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1092));
  INV_X1    g667(.A(G1348), .ZN(new_n1093));
  INV_X1    g668(.A(G2067), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n974), .A2(new_n982), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n986), .A2(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(new_n841), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1091), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1091), .B(KEYINPUT120), .C1(new_n1092), .C2(new_n1097), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n841), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1096), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n841), .A2(new_n1103), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1092), .A2(KEYINPUT122), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1086), .A2(KEYINPUT122), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1091), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n1112), .C2(new_n1092), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1107), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  OR3_X1    g689(.A1(new_n980), .A2(KEYINPUT121), .A3(G1996), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT58), .B(G1341), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n991), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT121), .B1(new_n980), .B2(G1996), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n809), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT59), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1122), .A3(new_n809), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1102), .B1(new_n1114), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1042), .B1(new_n1084), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1042), .B(KEYINPUT126), .C1(new_n1084), .C2(new_n1125), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1077), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1079), .ZN(new_n1131));
  OR3_X1    g706(.A1(new_n1130), .A2(KEYINPUT62), .A3(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1082), .A2(G171), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1069), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT62), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1128), .A2(new_n1129), .A3(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n976), .A2(new_n982), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n806), .B(new_n1094), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(KEYINPUT116), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1142), .A2(KEYINPUT116), .ZN(new_n1144));
  INV_X1    g719(.A(G1996), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n720), .B(new_n1145), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n1143), .B(new_n1144), .C1(new_n1138), .C2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n762), .B(new_n766), .Z(new_n1148));
  OAI21_X1  g723(.A(new_n1147), .B1(new_n1139), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n597), .B(G1986), .Z(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1138), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1137), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1139), .B1(new_n720), .B2(new_n1140), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT46), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1138), .A2(new_n1145), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT47), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1139), .A2(G1986), .A3(G290), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT48), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1149), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1147), .A2(new_n763), .A3(new_n766), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n867), .A2(new_n1094), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1139), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1152), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g741(.A1(G319), .A2(new_n660), .A3(new_n678), .ZN(new_n1168));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n1169));
  OR2_X1    g743(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n698), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n888), .A2(new_n889), .ZN(new_n1173));
  NOR3_X1   g747(.A1(new_n970), .A2(new_n1172), .A3(new_n1173), .ZN(G308));
  AND3_X1   g748(.A1(new_n698), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1175));
  INV_X1    g749(.A(new_n1173), .ZN(new_n1176));
  AND2_X1   g750(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n1175), .B(new_n1176), .C1(new_n1177), .C2(new_n968), .ZN(G225));
endmodule


