//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT26), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT69), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n202), .A2(new_n203), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n207), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n204), .A2(new_n205), .A3(new_n206), .A4(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT27), .B(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  OR2_X1    g010(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n212));
  NAND2_X1  g011(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n211), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n213), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n209), .A2(new_n214), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  OAI211_X1 g024(.A(G183gat), .B(G190gat), .C1(KEYINPUT67), .C2(KEYINPUT24), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n202), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT25), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(G176gat), .ZN(new_n235));
  AND2_X1   g034(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT25), .B1(new_n228), .B2(new_n229), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n220), .A2(new_n223), .ZN(new_n242));
  NAND3_X1  g041(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n225), .A3(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n235), .B(KEYINPUT66), .C1(new_n237), .C2(new_n236), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n240), .A2(new_n241), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n221), .A2(new_n233), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G127gat), .B(G134gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(KEYINPUT1), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n248), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n251), .A2(new_n254), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n257), .A2(new_n221), .A3(new_n233), .A4(new_n246), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT64), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G15gat), .B(G43gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(G99gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT72), .B(G71gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT33), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(KEYINPUT32), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT33), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n262), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n261), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(new_n256), .B2(new_n258), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT70), .B1(new_n273), .B2(KEYINPUT33), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(new_n266), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n262), .A2(new_n276), .A3(KEYINPUT32), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT32), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT71), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n268), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n256), .A2(new_n272), .A3(new_n258), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT34), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(new_n272), .B2(KEYINPUT73), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n282), .B(new_n284), .Z(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n285), .B(new_n268), .C1(new_n275), .C2(new_n280), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OR3_X1    g089(.A1(new_n281), .A2(new_n286), .A3(new_n288), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G197gat), .B(G204gat), .ZN(new_n296));
  INV_X1    g095(.A(G211gat), .ZN(new_n297));
  INV_X1    g096(.A(G218gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n296), .B1(KEYINPUT22), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n295), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G155gat), .ZN(new_n303));
  INV_X1    g102(.A(G162gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT2), .ZN(new_n306));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT82), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(G148gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n321));
  OAI21_X1  g120(.A(G141gat), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT83), .B1(new_n322), .B2(new_n317), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n309), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n312), .A2(G141gat), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT2), .B1(new_n317), .B2(new_n326), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n327), .A2(new_n305), .A3(new_n307), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n302), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G228gat), .ZN(new_n335));
  INV_X1    g134(.A(G233gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n316), .B1(new_n315), .B2(new_n318), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n322), .A2(KEYINPUT83), .A3(new_n317), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n308), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(new_n328), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT3), .B1(new_n302), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n334), .B(new_n337), .C1(new_n341), .C2(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n300), .A2(new_n293), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n300), .A2(new_n293), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n332), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n341), .B1(new_n325), .B2(new_n347), .ZN(new_n348));
  OAI22_X1  g147(.A1(new_n333), .A2(new_n348), .B1(new_n335), .B2(new_n336), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G22gat), .ZN(new_n351));
  XOR2_X1   g150(.A(KEYINPUT31), .B(G50gat), .Z(new_n352));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT87), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n355), .B1(new_n350), .B2(G22gat), .ZN(new_n357));
  INV_X1    g156(.A(G22gat), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n344), .A2(new_n349), .A3(new_n358), .A4(new_n354), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n360), .B2(new_n351), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n292), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT3), .B1(new_n340), .B2(new_n328), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(new_n330), .A3(new_n255), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(new_n341), .B2(new_n257), .ZN(new_n367));
  NOR4_X1   g166(.A1(new_n340), .A2(new_n255), .A3(new_n328), .A4(KEYINPUT4), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n364), .B(new_n365), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n324), .A2(new_n329), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n255), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n324), .A2(new_n257), .A3(new_n329), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n365), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(KEYINPUT4), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n324), .A2(new_n257), .A3(new_n366), .A4(new_n329), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n381), .A2(new_n365), .A3(new_n364), .A4(new_n370), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n372), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384));
  INV_X1    g183(.A(G85gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT0), .B(G57gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n372), .A2(new_n388), .A3(new_n378), .A4(new_n382), .ZN(new_n391));
  XOR2_X1   g190(.A(KEYINPUT85), .B(KEYINPUT6), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n391), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n247), .A2(new_n342), .ZN(new_n398));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(KEYINPUT77), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n247), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n302), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n399), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n247), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n401), .B1(new_n247), .B2(new_n332), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n301), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT79), .B(G8gat), .ZN(new_n408));
  INV_X1    g207(.A(G36gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n403), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT81), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT30), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n403), .A2(new_n407), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n412), .B(KEYINPUT80), .Z(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n414), .A2(KEYINPUT81), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT88), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n416), .A2(KEYINPUT88), .A3(new_n419), .A4(new_n421), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n362), .A2(new_n397), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT35), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n287), .A2(new_n289), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n361), .A2(new_n429), .A3(new_n428), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n392), .B1(new_n383), .B2(new_n389), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n431), .A2(KEYINPUT86), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n395), .B1(new_n431), .B2(KEYINPUT86), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n432), .A2(new_n433), .B1(new_n395), .B2(new_n392), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(new_n422), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n427), .A2(new_n428), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(KEYINPUT90), .B(KEYINPUT39), .Z(new_n437));
  INV_X1    g236(.A(KEYINPUT89), .ZN(new_n438));
  AOI211_X1 g237(.A(new_n438), .B(new_n365), .C1(new_n381), .C2(new_n364), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT89), .B1(new_n440), .B2(new_n377), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n437), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n257), .B1(new_n373), .B2(KEYINPUT3), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n330), .A2(new_n443), .B1(new_n379), .B2(new_n380), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n438), .B1(new_n444), .B2(new_n365), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n374), .A2(new_n365), .A3(new_n375), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n446), .A2(KEYINPUT39), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(KEYINPUT89), .A3(new_n377), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n442), .A2(new_n449), .A3(new_n389), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT40), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n442), .A2(new_n449), .A3(KEYINPUT40), .A4(new_n389), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n452), .A2(new_n391), .A3(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n424), .A2(new_n425), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT91), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n417), .A2(KEYINPUT37), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n412), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n417), .A2(KEYINPUT37), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT38), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AND4_X1   g260(.A1(new_n396), .A2(new_n394), .A3(new_n414), .A4(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n460), .A2(KEYINPUT38), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n400), .A2(new_n301), .A3(new_n402), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n302), .B1(new_n405), .B2(new_n406), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT37), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n418), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n361), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n391), .A3(new_n453), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT91), .B1(new_n469), .B2(new_n426), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n457), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n287), .A2(KEYINPUT36), .A3(new_n289), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT74), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n287), .A2(KEYINPUT74), .A3(KEYINPUT36), .A4(new_n289), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n290), .A2(new_n291), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n361), .B1(new_n434), .B2(new_n422), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n471), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n436), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT92), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n436), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT16), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(G1gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(G1gat), .B2(new_n486), .ZN(new_n489));
  INV_X1    g288(.A(G8gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT97), .ZN(new_n492));
  OR3_X1    g291(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n493), .A2(new_n494), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT96), .ZN(new_n497));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT95), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G43gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(G50gat), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT15), .B1(new_n502), .B2(KEYINPUT95), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n497), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G50gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G43gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT94), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n498), .A2(KEYINPUT94), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT15), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n496), .B1(new_n505), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n509), .A2(new_n510), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n498), .A2(KEYINPUT94), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n497), .A3(new_n503), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n517), .A2(KEYINPUT15), .B1(new_n518), .B2(new_n495), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n492), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n513), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n495), .B1(new_n521), .B2(new_n504), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(new_n495), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n513), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(KEYINPUT97), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n491), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(new_n522), .B2(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(new_n525), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(new_n527), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n526), .B1(new_n530), .B2(new_n491), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n532), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n514), .A2(new_n519), .A3(new_n492), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT97), .B1(new_n522), .B2(new_n524), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n527), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n528), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n491), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n526), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n532), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n520), .A2(new_n525), .A3(new_n491), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n532), .B(KEYINPUT13), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n533), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  INV_X1    g348(.A(G197gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT11), .B(G169gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT93), .B(KEYINPUT12), .Z(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  AOI21_X1  g354(.A(KEYINPUT18), .B1(new_n531), .B2(new_n532), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(KEYINPUT98), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n555), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n542), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n533), .A2(new_n542), .A3(new_n547), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n483), .A2(new_n485), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G57gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(G64gat), .ZN(new_n567));
  INV_X1    g366(.A(G64gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G57gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(KEYINPUT9), .B2(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n571), .A2(KEYINPUT99), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n571), .A2(KEYINPUT99), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n574), .A2(KEYINPUT100), .A3(new_n571), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT100), .B1(new_n574), .B2(new_n571), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n578), .B(new_n570), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT101), .B(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT102), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n577), .A2(new_n588), .A3(new_n581), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n577), .B2(new_n581), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT21), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n491), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT103), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n593), .A2(new_n595), .ZN(new_n598));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n601), .ZN(new_n603));
  INV_X1    g402(.A(new_n593), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n594), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n603), .B1(new_n605), .B2(new_n596), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n587), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n601), .B1(new_n597), .B2(new_n598), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n596), .A3(new_n603), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n586), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  INV_X1    g411(.A(G92gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(KEYINPUT8), .A2(new_n612), .B1(new_n385), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(new_n385), .B2(new_n613), .ZN(new_n616));
  NAND3_X1  g415(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G99gat), .B(G106gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n530), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n619), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n618), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n529), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625));
  NAND2_X1  g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT104), .Z(new_n627));
  OAI211_X1 g426(.A(new_n621), .B(new_n624), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n625), .ZN(new_n629));
  XOR2_X1   g428(.A(G134gat), .B(G162gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G190gat), .B(G218gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n628), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(G230gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n336), .ZN(new_n637));
  OAI211_X1 g436(.A(KEYINPUT10), .B(new_n623), .C1(new_n589), .C2(new_n590), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n581), .A3(new_n577), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n582), .A2(new_n620), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT105), .B(KEYINPUT10), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n637), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  AOI211_X1 g442(.A(new_n636), .B(new_n336), .C1(new_n639), .C2(new_n640), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n611), .A2(new_n635), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n565), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n434), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g454(.A1(new_n565), .A2(new_n426), .A3(new_n652), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT16), .B(G8gat), .Z(new_n657));
  AND2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n659), .B(new_n660), .C1(new_n490), .C2(new_n656), .ZN(G1325gat));
  INV_X1    g460(.A(new_n292), .ZN(new_n662));
  AOI21_X1  g461(.A(G15gat), .B1(new_n653), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n479), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n476), .A2(KEYINPUT106), .A3(new_n478), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n663), .B1(new_n653), .B2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n361), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  INV_X1    g472(.A(new_n651), .ZN(new_n674));
  NOR4_X1   g473(.A1(new_n565), .A2(new_n611), .A3(new_n635), .A4(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(G29gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n434), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n427), .A2(new_n428), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n435), .A2(new_n430), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n476), .A2(KEYINPUT106), .A3(new_n478), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT106), .B1(new_n476), .B2(new_n478), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n471), .B(new_n480), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n667), .A2(KEYINPUT108), .A3(new_n480), .A4(new_n471), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n682), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n679), .B1(new_n689), .B2(new_n635), .ZN(new_n690));
  INV_X1    g489(.A(new_n611), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n651), .B(KEYINPUT107), .Z(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n564), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n483), .A2(KEYINPUT44), .A3(new_n485), .A4(new_n634), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n690), .A2(new_n691), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n434), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n678), .A2(new_n699), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n675), .A2(new_n409), .A3(new_n455), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n702));
  OAI21_X1  g501(.A(G36gat), .B1(new_n697), .B2(new_n426), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(G1329gat));
  AND3_X1   g504(.A1(new_n690), .A2(new_n691), .A3(new_n696), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n706), .A2(G43gat), .A3(new_n668), .A4(new_n695), .ZN(new_n707));
  INV_X1    g506(.A(new_n565), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n611), .A2(new_n674), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n708), .A2(new_n662), .A3(new_n634), .A4(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT109), .B1(new_n710), .B2(new_n501), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n707), .A2(KEYINPUT47), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT47), .B1(new_n707), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1330gat));
  NAND4_X1  g513(.A1(new_n706), .A2(G50gat), .A3(new_n361), .A4(new_n695), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n675), .A2(new_n361), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(G50gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n361), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n697), .A2(new_n506), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(G50gat), .B1(new_n675), .B2(new_n361), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT48), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(G1331gat));
  NOR3_X1   g522(.A1(new_n689), .A2(new_n691), .A3(new_n634), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n692), .A2(new_n564), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n698), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n566), .ZN(G1332gat));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n426), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  NAND4_X1  g532(.A1(new_n724), .A2(G71gat), .A3(new_n668), .A4(new_n725), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n726), .A2(new_n292), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(G71gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT50), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n738), .B(new_n734), .C1(new_n735), .C2(G71gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1334gat));
  NOR2_X1   g539(.A1(new_n726), .A2(new_n719), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g541(.A1(new_n698), .A2(G85gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n687), .A2(new_n688), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n635), .B1(new_n744), .B2(new_n436), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n611), .A2(new_n564), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  INV_X1    g547(.A(new_n746), .ZN(new_n749));
  NOR4_X1   g548(.A1(new_n689), .A2(new_n748), .A3(new_n635), .A4(new_n749), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n674), .B(new_n743), .C1(new_n747), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n690), .A2(new_n696), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n651), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n752), .A2(new_n698), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n751), .B1(new_n755), .B2(new_n385), .ZN(G1336gat));
  NOR2_X1   g555(.A1(new_n426), .A2(G92gat), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n693), .B(new_n757), .C1(new_n747), .C2(new_n750), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n690), .A2(new_n455), .A3(new_n696), .A4(new_n753), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G92gat), .ZN(new_n760));
  AOI211_X1 g559(.A(KEYINPUT110), .B(KEYINPUT52), .C1(new_n758), .C2(new_n760), .ZN(new_n761));
  OR2_X1    g560(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n762));
  NAND2_X1  g561(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n763));
  AND4_X1   g562(.A1(new_n762), .A2(new_n758), .A3(new_n763), .A4(new_n760), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n761), .A2(new_n764), .ZN(G1337gat));
  NOR2_X1   g564(.A1(new_n292), .A2(G99gat), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n674), .B(new_n766), .C1(new_n747), .C2(new_n750), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n667), .A3(new_n754), .ZN(new_n768));
  INV_X1    g567(.A(G99gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(G1338gat));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n719), .A2(G106gat), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n693), .B(new_n772), .C1(new_n747), .C2(new_n750), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n690), .A2(new_n361), .A3(new_n696), .A4(new_n753), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G106gat), .ZN(new_n775));
  AOI211_X1 g574(.A(new_n771), .B(KEYINPUT53), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n771), .A2(KEYINPUT53), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n771), .A2(KEYINPUT53), .ZN(new_n778));
  AND4_X1   g577(.A1(new_n777), .A2(new_n773), .A3(new_n778), .A4(new_n775), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n776), .A2(new_n779), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n643), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n638), .A2(new_n642), .A3(new_n637), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT54), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n783), .B(new_n648), .C1(new_n785), .C2(new_n643), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n781), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n785), .A2(new_n643), .ZN(new_n789));
  INV_X1    g588(.A(new_n648), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n643), .B2(new_n782), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n789), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n786), .A2(new_n787), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n788), .A2(new_n792), .A3(new_n649), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n558), .B2(new_n563), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n533), .A2(new_n542), .A3(new_n559), .A4(new_n547), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n531), .A2(new_n532), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n544), .A2(new_n546), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n553), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n651), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n635), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n635), .A2(new_n800), .A3(new_n794), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n611), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n652), .A2(new_n564), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n698), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n361), .A2(new_n429), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n809), .A2(new_n426), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(G113gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n812), .A3(new_n564), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n809), .A2(new_n426), .A3(new_n362), .ZN(new_n814));
  OAI21_X1  g613(.A(G113gat), .B1(new_n814), .B2(new_n694), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(G1340gat));
  INV_X1    g615(.A(G120gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n811), .A2(new_n817), .A3(new_n674), .ZN(new_n818));
  OAI21_X1  g617(.A(G120gat), .B1(new_n814), .B2(new_n692), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1341gat));
  INV_X1    g619(.A(G127gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n814), .A2(new_n821), .A3(new_n691), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n811), .A2(new_n611), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT113), .Z(new_n824));
  AOI21_X1  g623(.A(new_n822), .B1(new_n824), .B2(new_n821), .ZN(G1342gat));
  INV_X1    g624(.A(G134gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n826), .A3(new_n634), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT56), .Z(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n814), .B2(new_n635), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1343gat));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n361), .B1(new_n805), .B2(new_n807), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n667), .A2(new_n434), .A3(new_n426), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND4_X1   g633(.A1(KEYINPUT116), .A2(new_n834), .A3(new_n310), .A4(new_n564), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n788), .A2(new_n792), .A3(new_n649), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n787), .B1(new_n786), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT114), .B1(new_n789), .B2(new_n791), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI211_X1 g639(.A(new_n836), .B(new_n840), .C1(new_n558), .C2(new_n563), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n635), .B1(new_n841), .B2(new_n801), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n611), .B1(new_n842), .B2(new_n804), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT57), .B(new_n361), .C1(new_n843), .C2(new_n807), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n832), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n846), .A3(KEYINPUT115), .ZN(new_n847));
  INV_X1    g646(.A(new_n836), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n564), .B(new_n848), .C1(new_n839), .C2(new_n838), .ZN(new_n849));
  INV_X1    g648(.A(new_n801), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n803), .B1(new_n851), .B2(new_n635), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n808), .B1(new_n852), .B2(new_n611), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT57), .A4(new_n361), .ZN(new_n855));
  INV_X1    g654(.A(new_n833), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n847), .A2(new_n855), .A3(new_n564), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n835), .B1(new_n857), .B2(G141gat), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT58), .B1(new_n858), .B2(KEYINPUT117), .ZN(new_n859));
  NOR4_X1   g658(.A1(new_n832), .A2(new_n833), .A3(G141gat), .A4(new_n694), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(KEYINPUT117), .B2(KEYINPUT58), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n860), .B(new_n862), .C1(new_n857), .C2(G141gat), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n831), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n860), .B1(new_n857), .B2(G141gat), .ZN(new_n865));
  INV_X1    g664(.A(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n868), .B(new_n835), .C1(new_n857), .C2(G141gat), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT118), .B(new_n867), .C1(new_n869), .C2(KEYINPUT58), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n864), .A2(new_n870), .ZN(G1344gat));
  NAND2_X1  g670(.A1(new_n313), .A2(new_n314), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n834), .A2(new_n872), .A3(new_n674), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n847), .A2(new_n855), .A3(new_n856), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n651), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n872), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n853), .B2(new_n361), .ZN(new_n878));
  OAI211_X1 g677(.A(KEYINPUT57), .B(new_n361), .C1(new_n805), .C2(new_n807), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n674), .B(new_n856), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n874), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n873), .B1(new_n877), .B2(new_n882), .ZN(G1345gat));
  NOR3_X1   g682(.A1(new_n875), .A2(new_n303), .A3(new_n691), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n834), .A2(new_n611), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT119), .Z(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n303), .B2(new_n886), .ZN(G1346gat));
  NAND3_X1  g686(.A1(new_n834), .A2(new_n304), .A3(new_n634), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT120), .Z(new_n889));
  OAI21_X1  g688(.A(G162gat), .B1(new_n875), .B2(new_n635), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT121), .ZN(G1347gat));
  NOR2_X1   g691(.A1(new_n434), .A2(new_n426), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n806), .B2(new_n808), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n810), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n236), .A2(new_n237), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(new_n694), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT122), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(new_n362), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n694), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1348gat));
  NOR2_X1   g701(.A1(new_n896), .A2(new_n651), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n693), .A2(G176gat), .ZN(new_n904));
  OAI22_X1  g703(.A1(new_n903), .A2(G176gat), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT123), .Z(G1349gat));
  OAI21_X1  g705(.A(G183gat), .B1(new_n900), .B2(new_n691), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n611), .A2(new_n210), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n896), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n911));
  OAI21_X1  g710(.A(G190gat), .B1(new_n900), .B2(new_n635), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n913), .B2(KEYINPUT124), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(KEYINPUT124), .B2(new_n913), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n895), .A2(new_n211), .A3(new_n810), .A4(new_n634), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n913), .A2(KEYINPUT124), .A3(KEYINPUT61), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G1351gat));
  NOR2_X1   g717(.A1(new_n668), .A2(new_n894), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n832), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n921), .A2(KEYINPUT125), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(KEYINPUT125), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n922), .A2(new_n550), .A3(new_n564), .A4(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(KEYINPUT126), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(KEYINPUT126), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n878), .A2(new_n880), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n694), .A3(new_n920), .ZN(new_n928));
  OAI22_X1  g727(.A1(new_n925), .A2(new_n926), .B1(new_n550), .B2(new_n928), .ZN(G1352gat));
  INV_X1    g728(.A(G204gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n921), .A2(new_n930), .A3(new_n674), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT62), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n927), .A2(new_n920), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n693), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n932), .A2(new_n934), .ZN(G1353gat));
  NAND4_X1  g734(.A1(new_n922), .A2(new_n297), .A3(new_n611), .A4(new_n923), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n611), .B(new_n919), .C1(new_n878), .C2(new_n880), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n937), .B2(G211gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g741(.A(KEYINPUT127), .B(new_n936), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1354gat));
  NAND3_X1  g743(.A1(new_n922), .A2(new_n634), .A3(new_n923), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n635), .A2(new_n298), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n945), .A2(new_n298), .B1(new_n933), .B2(new_n946), .ZN(G1355gat));
endmodule


