//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G101), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT66), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G137), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(KEYINPUT66), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(G137), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n201), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n200), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n204), .A2(G134), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n208), .B1(new_n196), .B2(new_n198), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n202), .A2(KEYINPUT11), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n203), .B1(new_n211), .B2(new_n205), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT65), .B1(new_n215), .B2(G143), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G146), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n215), .A2(KEYINPUT64), .A3(G143), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT64), .B1(new_n215), .B2(G143), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n216), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n222), .A2(new_n225), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n214), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(G131), .B1(new_n198), .B2(new_n208), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n215), .A2(G143), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n216), .A2(new_n219), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n215), .A2(KEYINPUT64), .A3(G143), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n232), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n218), .A2(G146), .ZN(new_n240));
  AND4_X1   g054(.A1(new_n239), .A2(new_n231), .A3(new_n240), .A4(G128), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n213), .B(new_n229), .C1(new_n238), .C2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT68), .B1(new_n243), .B2(G119), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G116), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(G119), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G113), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT2), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G113), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n253), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n256), .A2(new_n244), .A3(new_n247), .A4(new_n248), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n228), .A2(new_n242), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n228), .A2(new_n242), .A3(KEYINPUT28), .A4(new_n259), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n213), .A2(new_n229), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n213), .A2(new_n267), .A3(new_n229), .ZN(new_n268));
  INV_X1    g082(.A(new_n232), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n222), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n231), .A2(new_n240), .A3(new_n239), .A4(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n228), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n258), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n194), .B1(new_n264), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n194), .A2(KEYINPUT70), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n228), .B2(new_n242), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n241), .B1(new_n222), .B2(new_n269), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n265), .B2(KEYINPUT67), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n281), .A2(new_n268), .B1(new_n214), .B2(new_n227), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(new_n282), .B2(new_n278), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n260), .B(new_n277), .C1(new_n283), .C2(new_n259), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n260), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n273), .A2(new_n278), .A3(new_n228), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n228), .A2(new_n242), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT30), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n291), .B2(new_n258), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT31), .A3(new_n277), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n276), .B1(new_n286), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n187), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT71), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n294), .A2(new_n296), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT32), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n194), .A2(KEYINPUT29), .ZN(new_n302));
  INV_X1    g116(.A(new_n262), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n260), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n228), .A2(new_n242), .A3(KEYINPUT73), .A4(new_n259), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n289), .A2(new_n258), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n302), .B(new_n303), .C1(new_n308), .C2(KEYINPUT28), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n301), .B1(new_n309), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n262), .B1(new_n312), .B2(new_n261), .ZN(new_n313));
  OAI211_X1 g127(.A(KEYINPUT74), .B(new_n311), .C1(new_n313), .C2(new_n302), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n275), .A2(new_n263), .A3(new_n194), .A4(new_n262), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT29), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n260), .B1(new_n283), .B2(new_n259), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n193), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n264), .A2(KEYINPUT72), .A3(new_n194), .A4(new_n275), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n310), .A2(new_n314), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G472), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n324), .B(new_n187), .C1(new_n294), .C2(new_n296), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n298), .A2(new_n300), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G478), .ZN(new_n329));
  NOR2_X1   g143(.A1(KEYINPUT100), .A2(KEYINPUT15), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(KEYINPUT100), .A2(KEYINPUT15), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT9), .B(G234), .ZN(new_n335));
  INV_X1    g149(.A(G217), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n335), .A2(new_n336), .A3(G953), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT13), .B1(new_n218), .B2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n218), .A2(G128), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n340), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n341), .A2(KEYINPUT98), .B1(KEYINPUT13), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT98), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n339), .A2(new_n344), .A3(new_n340), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n197), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n230), .A2(G143), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n347), .A3(new_n197), .ZN(new_n348));
  INV_X1    g162(.A(G122), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G116), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n243), .A2(G122), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(G107), .ZN(new_n353));
  INV_X1    g167(.A(G107), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n350), .B2(new_n351), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n348), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT99), .B1(new_n346), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n348), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n197), .B1(new_n340), .B2(new_n347), .ZN(new_n359));
  OAI22_X1  g173(.A1(new_n358), .A2(new_n359), .B1(G107), .B2(new_n352), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT14), .ZN(new_n361));
  OAI21_X1  g175(.A(G107), .B1(new_n351), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n352), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(new_n361), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n357), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n356), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n341), .A2(KEYINPUT98), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n342), .A2(KEYINPUT13), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n345), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G134), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT99), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n368), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n338), .B1(new_n367), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n368), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n365), .B1(new_n377), .B2(KEYINPUT99), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n374), .A3(new_n337), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n334), .B1(new_n380), .B2(new_n311), .ZN(new_n381));
  AOI211_X1 g195(.A(G902), .B(new_n333), .C1(new_n376), .C2(new_n379), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G237), .ZN(new_n384));
  INV_X1    g198(.A(G953), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G214), .ZN(new_n386));
  NOR2_X1   g200(.A1(KEYINPUT94), .A2(G143), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n189), .B(G214), .C1(KEYINPUT94), .C2(G143), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT18), .A3(G131), .ZN(new_n391));
  XNOR2_X1  g205(.A(G125), .B(G140), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(new_n215), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT18), .A2(G131), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  XOR2_X1   g210(.A(G113), .B(G122), .Z(new_n397));
  INV_X1    g211(.A(G104), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G104), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT95), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT95), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n399), .B2(new_n401), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT96), .ZN(new_n407));
  AND4_X1   g221(.A1(new_n407), .A2(new_n390), .A3(KEYINPUT17), .A4(G131), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n210), .B1(new_n388), .B2(new_n389), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n409), .B2(KEYINPUT17), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n390), .A2(G131), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n388), .A2(new_n389), .A3(new_n210), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G125), .ZN(new_n417));
  INV_X1    g231(.A(G125), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G140), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT16), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n418), .A2(KEYINPUT16), .A3(G140), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n420), .A2(G146), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(G146), .B1(new_n420), .B2(new_n421), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n396), .B(new_n406), .C1(new_n411), .C2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n421), .A3(G146), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT19), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n392), .B(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n427), .B1(new_n429), .B2(G146), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n388), .A2(new_n389), .A3(new_n210), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(new_n409), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n396), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n402), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n436));
  NOR2_X1   g250(.A1(G475), .A2(G902), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT97), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n426), .A2(new_n434), .ZN(new_n440));
  INV_X1    g254(.A(new_n437), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT20), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT97), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n435), .A2(new_n443), .A3(new_n436), .A4(new_n437), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n396), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n420), .A2(new_n421), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n215), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n427), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n413), .B2(new_n432), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT96), .B1(new_n412), .B2(new_n413), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n409), .A2(new_n407), .A3(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n446), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n402), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n426), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n311), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G475), .ZN(new_n458));
  INV_X1    g272(.A(G952), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(G953), .ZN(new_n460));
  INV_X1    g274(.A(G234), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(new_n384), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(G898), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(G902), .B(G953), .C1(new_n461), .C2(new_n384), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT101), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n383), .A2(new_n445), .A3(new_n458), .A4(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G210), .B1(G237), .B2(G902), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT3), .B1(new_n398), .B2(G107), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT3), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n354), .A3(G104), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n398), .A2(G107), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G101), .ZN(new_n476));
  INV_X1    g290(.A(G101), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n471), .A2(new_n473), .A3(new_n477), .A4(new_n474), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(KEYINPUT4), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT4), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n475), .A2(new_n480), .A3(G101), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n258), .A3(new_n481), .ZN(new_n482));
  OR2_X1    g296(.A1(KEYINPUT87), .A2(KEYINPUT5), .ZN(new_n483));
  NAND2_X1  g297(.A1(KEYINPUT87), .A2(KEYINPUT5), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(G116), .A3(new_n246), .A4(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT87), .B(KEYINPUT5), .Z(new_n486));
  OAI211_X1 g300(.A(G113), .B(new_n485), .C1(new_n249), .C2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G104), .B(G107), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT82), .B1(new_n488), .B2(new_n477), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n354), .A2(G104), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n474), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT82), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(G101), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n487), .A2(new_n494), .A3(new_n257), .A4(new_n478), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n482), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G110), .B(G122), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n272), .A2(new_n418), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n227), .A2(G125), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G224), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(G953), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n503), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n482), .A2(new_n495), .A3(new_n497), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n482), .A2(new_n495), .A3(KEYINPUT89), .A4(new_n497), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n499), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n497), .B1(new_n482), .B2(new_n495), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(KEYINPUT88), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT90), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n513), .A2(new_n518), .A3(new_n515), .A4(new_n521), .ZN(new_n522));
  AOI211_X1 g336(.A(new_n500), .B(new_n508), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n506), .A2(KEYINPUT93), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n501), .A2(new_n502), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n506), .A2(KEYINPUT7), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n513), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT91), .B(KEYINPUT8), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n497), .B(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n487), .A2(new_n257), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n494), .A2(new_n478), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n489), .A2(new_n493), .B1(new_n538), .B2(new_n477), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT5), .ZN(new_n540));
  OAI211_X1 g354(.A(G113), .B(new_n485), .C1(new_n249), .C2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n257), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n532), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n311), .B1(new_n529), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n470), .B1(new_n523), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n500), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n517), .A2(KEYINPUT88), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n514), .B(new_n497), .C1(new_n482), .C2(new_n495), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n547), .A2(new_n548), .A3(new_n516), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n521), .B1(new_n549), .B2(new_n513), .ZN(new_n550));
  INV_X1    g364(.A(new_n522), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n546), .B(new_n507), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n544), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n469), .ZN(new_n554));
  AOI211_X1 g368(.A(new_n328), .B(new_n468), .C1(new_n545), .C2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT23), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n246), .B2(G128), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n246), .A2(G128), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n230), .A2(KEYINPUT23), .A3(G119), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G119), .B(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n556), .A2(KEYINPUT24), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT24), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G110), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n562), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n449), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n558), .A2(new_n561), .A3(new_n556), .A4(new_n559), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n230), .A2(G119), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n559), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT24), .B(G110), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n571), .B2(new_n572), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n570), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n571), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT75), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n582), .A2(new_n573), .A3(KEYINPUT76), .A4(new_n578), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n392), .A2(new_n215), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n427), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT77), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT77), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n589), .B(new_n586), .C1(new_n580), .C2(new_n583), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n569), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT22), .B(G137), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n385), .A2(G221), .A3(G234), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n594), .B(KEYINPUT78), .Z(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n336), .B1(G234), .B2(new_n311), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(G902), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(KEYINPUT79), .Z(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n569), .B(new_n594), .C1(new_n588), .C2(new_n590), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n569), .ZN(new_n604));
  INV_X1    g418(.A(new_n579), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT76), .B1(new_n605), .B2(new_n573), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n574), .A2(new_n579), .A3(new_n570), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n587), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n589), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n584), .A2(KEYINPUT77), .A3(new_n587), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n311), .B(new_n602), .C1(new_n611), .C2(new_n595), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT25), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n597), .A2(KEYINPUT25), .A3(new_n311), .A4(new_n602), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n603), .B1(new_n616), .B2(new_n598), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT85), .ZN(new_n618));
  XNOR2_X1  g432(.A(G110), .B(G140), .ZN(new_n619));
  INV_X1    g433(.A(G227), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(G953), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n619), .B(new_n621), .Z(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(KEYINPUT81), .Z(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n271), .B1(new_n232), .B2(new_n226), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n492), .B1(new_n491), .B2(G101), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT82), .B(new_n477), .C1(new_n490), .C2(new_n474), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n625), .B(new_n478), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n272), .B2(new_n539), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT12), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT84), .B1(new_n207), .B2(new_n213), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n629), .B2(new_n631), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n272), .A2(new_n539), .A3(KEYINPUT10), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n214), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n227), .A2(new_n479), .A3(new_n481), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n635), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n624), .B1(new_n634), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n622), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n635), .A2(new_n637), .A3(new_n639), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n214), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n618), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n629), .A2(new_n631), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT12), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n640), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n640), .A2(new_n622), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n643), .A2(new_n214), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n649), .A2(new_n623), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT85), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n645), .A2(new_n653), .A3(G469), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n642), .A2(KEYINPUT86), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT86), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n640), .A2(new_n656), .A3(new_n622), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n655), .A2(new_n634), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n651), .A2(new_n640), .ZN(new_n659));
  INV_X1    g473(.A(new_n622), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(G469), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n311), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n311), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n654), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(G221), .B1(new_n335), .B2(G902), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT80), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n326), .A2(new_n555), .A3(new_n617), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT102), .B(G101), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G3));
  INV_X1    g489(.A(new_n467), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n328), .B(new_n676), .C1(new_n545), .C2(new_n554), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n329), .A2(new_n311), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n337), .B1(new_n378), .B2(new_n374), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n374), .A2(new_n357), .A3(new_n366), .A4(new_n337), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n311), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n679), .B1(new_n682), .B2(G478), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n367), .B2(new_n375), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(KEYINPUT33), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n380), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n376), .A2(new_n685), .A3(new_n379), .A4(KEYINPUT33), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n683), .B1(G478), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n445), .A2(new_n458), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n677), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n617), .A2(new_n670), .A3(new_n667), .ZN(new_n695));
  INV_X1    g509(.A(new_n299), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n294), .B2(G902), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT34), .B(G104), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G6));
  AOI21_X1  g516(.A(new_n328), .B1(new_n545), .B2(new_n554), .ZN(new_n703));
  INV_X1    g517(.A(new_n438), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n436), .B1(new_n435), .B2(new_n437), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n458), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n383), .A2(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n703), .A2(new_n467), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n699), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT104), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT35), .B(G107), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G9));
  NOR2_X1   g526(.A1(new_n596), .A2(KEYINPUT36), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n591), .B(new_n713), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n616), .A2(new_n598), .B1(new_n601), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n671), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n555), .A2(new_n716), .A3(new_n698), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT37), .B(G110), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G12));
  OAI21_X1  g533(.A(new_n462), .B1(new_n465), .B2(G900), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n458), .B(new_n720), .C1(new_n704), .C2(new_n705), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n383), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n500), .B1(new_n520), .B2(new_n522), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n544), .B(new_n470), .C1(new_n723), .C2(new_n507), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n469), .B1(new_n552), .B2(new_n553), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n327), .B(new_n722), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT105), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n545), .A2(new_n554), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n327), .A4(new_n722), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n727), .A2(new_n326), .A3(new_n730), .A4(new_n716), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G128), .ZN(G30));
  XNOR2_X1  g546(.A(new_n720), .B(KEYINPUT39), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n672), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT40), .Z(new_n735));
  INV_X1    g549(.A(new_n691), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n383), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n715), .A3(new_n327), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n318), .A2(new_n194), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n740), .B(new_n311), .C1(new_n194), .C2(new_n308), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G472), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n298), .A2(new_n300), .A3(new_n325), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n728), .B(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n735), .A2(new_n739), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G143), .ZN(G45));
  NAND3_X1  g561(.A1(new_n690), .A2(new_n691), .A3(new_n720), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n326), .A2(new_n716), .A3(new_n703), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G146), .ZN(G48));
  AOI21_X1  g565(.A(new_n663), .B1(new_n662), .B2(new_n311), .ZN(new_n752));
  AOI211_X1 g566(.A(G469), .B(G902), .C1(new_n658), .C2(new_n661), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n752), .A2(new_n753), .A3(new_n669), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n326), .A2(new_n617), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n677), .A2(new_n693), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT41), .B(G113), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  NAND2_X1  g573(.A1(new_n677), .A2(new_n707), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n243), .ZN(G18));
  OAI211_X1 g576(.A(new_n754), .B(new_n327), .C1(new_n724), .C2(new_n725), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n703), .A2(KEYINPUT108), .A3(new_n754), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n715), .A2(new_n468), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n326), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G119), .ZN(G21));
  NAND2_X1  g583(.A1(new_n682), .A2(new_n333), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n380), .A2(new_n311), .A3(new_n334), .ZN(new_n771));
  AOI221_X4 g585(.A(new_n676), .B1(new_n770), .B2(new_n771), .C1(new_n445), .C2(new_n458), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n286), .A2(new_n293), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n313), .A2(new_n193), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n295), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n617), .A2(new_n772), .A3(new_n776), .A4(new_n697), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(KEYINPUT109), .A3(new_n703), .A4(new_n754), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n617), .A2(new_n772), .A3(new_n776), .A4(new_n697), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n779), .B1(new_n763), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G122), .ZN(G24));
  NAND2_X1  g597(.A1(new_n776), .A2(new_n697), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n715), .A3(new_n748), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n765), .A2(new_n785), .A3(new_n766), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G125), .ZN(G27));
  NOR2_X1   g601(.A1(new_n724), .A2(new_n725), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n665), .B1(new_n652), .B2(G469), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n669), .B1(new_n664), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n788), .A2(new_n789), .A3(new_n327), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n545), .A2(new_n327), .A3(new_n791), .A4(new_n554), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT110), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n300), .A2(new_n323), .A3(new_n297), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(new_n617), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT42), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n748), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n326), .A2(new_n617), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n749), .A3(new_n795), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n801), .A2(new_n795), .A3(KEYINPUT111), .A4(new_n749), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n798), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n800), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G131), .ZN(G33));
  NAND3_X1  g623(.A1(new_n801), .A2(new_n722), .A3(new_n795), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G134), .ZN(G36));
  NAND2_X1  g625(.A1(new_n736), .A2(new_n690), .ZN(new_n812));
  OR2_X1    g626(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n813));
  NAND2_X1  g627(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n812), .A2(new_n814), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n698), .ZN(new_n818));
  INV_X1    g632(.A(new_n715), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT44), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n788), .A2(new_n327), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n820), .B2(new_n821), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT45), .B1(new_n645), .B2(new_n653), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n652), .A2(KEYINPUT45), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(G469), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n665), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT112), .B1(new_n829), .B2(KEYINPUT46), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n753), .B1(new_n829), .B2(KEYINPUT46), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT46), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n832), .B(new_n833), .C1(new_n828), .C2(new_n665), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n670), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n822), .A2(new_n824), .A3(new_n733), .A4(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(KEYINPUT114), .B(G137), .Z(new_n838));
  XNOR2_X1  g652(.A(new_n837), .B(new_n838), .ZN(G39));
  NAND2_X1  g653(.A1(new_n836), .A2(KEYINPUT47), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n835), .A2(new_n670), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT47), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n326), .A2(new_n823), .A3(new_n617), .A4(new_n748), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(G140), .ZN(G42));
  NOR3_X1   g661(.A1(new_n812), .A2(new_n328), .A3(new_n669), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n752), .A2(new_n753), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(KEYINPUT49), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n851), .B(new_n745), .C1(KEYINPUT49), .C2(new_n850), .ZN(new_n852));
  INV_X1    g666(.A(new_n617), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n743), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n728), .A2(new_n327), .A3(new_n737), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n715), .A2(new_n720), .A3(new_n791), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n743), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n731), .A2(new_n786), .A3(new_n858), .A4(new_n750), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n763), .A2(new_n764), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT108), .B1(new_n703), .B2(new_n754), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n326), .A2(new_n767), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n863), .A2(new_n864), .B1(new_n781), .B2(new_n778), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n692), .B1(new_n691), .B2(new_n383), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n677), .A2(new_n695), .A3(new_n698), .A4(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n673), .A2(new_n717), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n801), .B(new_n754), .C1(new_n694), .C2(new_n708), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n721), .A2(new_n381), .A3(new_n382), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n327), .A2(new_n545), .A3(new_n871), .A4(new_n554), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n326), .A2(new_n716), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n326), .A2(new_n872), .A3(new_n716), .A4(KEYINPUT115), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n795), .A2(new_n785), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n810), .A3(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n860), .A2(new_n870), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n731), .A2(new_n786), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n750), .A4(new_n858), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n859), .A2(new_n881), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n880), .A2(new_n808), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n870), .A2(new_n879), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n808), .A3(new_n883), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT116), .B1(new_n890), .B2(new_n886), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n877), .A2(new_n810), .A3(new_n878), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n782), .A2(new_n768), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n755), .B1(new_n756), .B2(new_n760), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n673), .A2(new_n867), .A3(new_n717), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AND4_X1   g710(.A1(new_n883), .A2(new_n892), .A3(new_n896), .A4(new_n889), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT53), .A4(new_n808), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n887), .A2(new_n891), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT54), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n897), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n904));
  AOI22_X1  g718(.A1(KEYINPUT116), .A2(new_n904), .B1(new_n885), .B2(new_n886), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n905), .B2(new_n899), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n892), .A2(new_n896), .A3(new_n883), .A4(new_n889), .ZN(new_n907));
  INV_X1    g721(.A(new_n800), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n806), .A2(new_n798), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n804), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n907), .A2(KEYINPUT53), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(KEYINPUT53), .B2(new_n885), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT117), .B1(new_n912), .B2(KEYINPUT54), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n902), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n754), .A2(new_n328), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT118), .B1(new_n745), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n462), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n815), .B2(new_n816), .ZN(new_n919));
  INV_X1    g733(.A(new_n784), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n617), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n745), .A2(KEYINPUT118), .A3(new_n916), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT119), .B(KEYINPUT50), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OR3_X1    g740(.A1(new_n745), .A2(KEYINPUT118), .A3(new_n916), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n922), .A3(new_n917), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT50), .B1(new_n928), .B2(KEYINPUT119), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n915), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NOR4_X1   g744(.A1(new_n823), .A2(new_n462), .A3(new_n669), .A4(new_n850), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n690), .A2(new_n691), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n854), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n817), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n920), .A2(new_n819), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n840), .B(new_n843), .C1(new_n670), .C2(new_n850), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n921), .A2(new_n919), .A3(new_n823), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT119), .B1(new_n923), .B2(new_n924), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT50), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(KEYINPUT120), .A3(new_n925), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n930), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT51), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n931), .A2(new_n797), .A3(new_n817), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT48), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n931), .A2(new_n693), .A3(new_n854), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n922), .A2(new_n863), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n948), .A2(new_n460), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  AOI211_X1 g765(.A(new_n945), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n926), .A2(new_n929), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT121), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n946), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n946), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n914), .A2(KEYINPUT122), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n459), .A2(new_n385), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT122), .B1(new_n914), .B2(new_n958), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n855), .B1(new_n961), .B2(new_n962), .ZN(G75));
  XNOR2_X1  g777(.A(new_n723), .B(new_n507), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT55), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n912), .A2(G902), .ZN(new_n966));
  INV_X1    g780(.A(G210), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n965), .B1(new_n968), .B2(KEYINPUT56), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n385), .A2(G952), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT123), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n912), .A2(KEYINPUT123), .A3(G902), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n470), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n965), .A2(KEYINPUT56), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(G51));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n828), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n665), .B(KEYINPUT57), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n912), .A2(KEYINPUT54), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n912), .A2(KEYINPUT54), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n662), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n970), .B1(new_n980), .B2(new_n986), .ZN(G54));
  AND2_X1   g801(.A1(KEYINPUT58), .A2(G475), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n974), .A2(new_n975), .A3(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n989), .A2(KEYINPUT124), .A3(new_n440), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n971), .B1(new_n989), .B2(new_n440), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT124), .B1(new_n989), .B2(new_n440), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(G60));
  XNOR2_X1  g807(.A(new_n678), .B(KEYINPUT59), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n689), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n983), .B2(new_n984), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n971), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n914), .A2(new_n994), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n998), .B2(new_n689), .ZN(G63));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT60), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n912), .A2(new_n714), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n912), .A2(new_n1002), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n597), .A2(new_n602), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n971), .B(new_n1003), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g822(.A(G953), .B1(new_n463), .B2(new_n504), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(new_n896), .B2(G953), .ZN(new_n1010));
  INV_X1    g824(.A(new_n723), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(G898), .B2(new_n385), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1010), .B(new_n1012), .ZN(G69));
  XNOR2_X1  g827(.A(new_n291), .B(new_n429), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(G900), .B(G953), .C1(new_n1015), .C2(G227), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(G227), .B2(new_n1015), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n846), .A2(new_n837), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n881), .A2(new_n750), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n1019), .A2(new_n746), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT62), .ZN(new_n1021));
  OR2_X1    g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  INV_X1    g837(.A(new_n734), .ZN(new_n1024));
  INV_X1    g838(.A(new_n823), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n801), .A2(new_n1024), .A3(new_n1025), .A4(new_n866), .ZN(new_n1026));
  AND4_X1   g840(.A1(new_n1018), .A2(new_n1022), .A3(new_n1023), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(G953), .B1(new_n1028), .B2(new_n1014), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n836), .A2(new_n733), .A3(new_n797), .A4(new_n856), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1019), .A2(new_n1030), .A3(new_n810), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1018), .A2(new_n808), .A3(new_n1031), .ZN(new_n1032));
  OR2_X1    g846(.A1(new_n1032), .A2(KEYINPUT125), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(KEYINPUT125), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1033), .A2(new_n1015), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1017), .B1(new_n1029), .B2(new_n1035), .ZN(G72));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT63), .Z(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1039), .B1(new_n1027), .B2(new_n896), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n971), .B1(new_n1040), .B2(new_n740), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n292), .A2(new_n193), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1033), .A2(new_n896), .A3(new_n1034), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1042), .B1(new_n1043), .B2(new_n1038), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1038), .B1(new_n319), .B2(KEYINPUT126), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n740), .A2(new_n1042), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1045), .B1(KEYINPUT126), .B2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT127), .Z(new_n1048));
  AOI211_X1 g862(.A(new_n1041), .B(new_n1044), .C1(new_n900), .C2(new_n1048), .ZN(G57));
endmodule


