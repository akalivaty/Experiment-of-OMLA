//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  OAI211_X1 g001(.A(new_n187), .B(G119), .C1(KEYINPUT72), .C2(KEYINPUT23), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G128), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT72), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n192), .B1(new_n190), .B2(G128), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n188), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G119), .B(G128), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT24), .B(G110), .Z(new_n196));
  AOI22_X1  g010(.A1(new_n194), .A2(G110), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n198), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G140), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT73), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G146), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n199), .B1(new_n208), .B2(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT73), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n197), .A2(new_n207), .A3(new_n213), .ZN(new_n214));
  OAI22_X1  g028(.A1(new_n194), .A2(G110), .B1(new_n195), .B2(new_n196), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n208), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n209), .A2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n215), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G137), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(G221), .A3(G234), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n223), .B(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n214), .A2(new_n222), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n214), .A2(new_n222), .A3(KEYINPUT75), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n214), .A2(new_n222), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT74), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT74), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n214), .A2(new_n222), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n226), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G217), .ZN(new_n238));
  INV_X1    g052(.A(G902), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n238), .B1(G234), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(G902), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n231), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT78), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n231), .A2(new_n237), .A3(new_n239), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT76), .B(KEYINPUT25), .Z(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT77), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n231), .A2(new_n237), .A3(KEYINPUT25), .A4(new_n239), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT77), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n245), .A2(new_n250), .A3(new_n246), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n244), .B1(new_n252), .B2(new_n240), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  AOI21_X1  g071(.A(G131), .B1(new_n256), .B2(G137), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT67), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n256), .A2(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n257), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NAND3_X1  g087(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT65), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G143), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n210), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n276), .B1(new_n217), .B2(new_n218), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n275), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n216), .A2(G146), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(G143), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n277), .A2(new_n279), .A3(G146), .ZN(new_n287));
  INV_X1    g101(.A(new_n270), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n269), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n286), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(G146), .B1(new_n277), .B2(new_n279), .ZN(new_n294));
  AOI21_X1  g108(.A(G143), .B1(new_n284), .B2(new_n285), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n187), .B1(new_n286), .B2(KEYINPUT1), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G131), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n259), .A2(G134), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n266), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n263), .B2(new_n264), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n291), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(KEYINPUT2), .B(G113), .Z(new_n305));
  XNOR2_X1  g119(.A(G116), .B(G119), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n307), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n291), .A2(new_n309), .A3(new_n303), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(KEYINPUT71), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n304), .A2(new_n312), .A3(new_n307), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(KEYINPUT28), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G237), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n224), .A3(G210), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT27), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n314), .A2(new_n316), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n310), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n291), .A2(new_n327), .A3(new_n303), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n291), .B2(new_n303), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n307), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n298), .A2(new_n302), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n263), .A2(new_n264), .B1(G131), .B2(new_n267), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n272), .A2(new_n274), .A3(new_n273), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n294), .B2(new_n295), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT30), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n291), .A2(new_n327), .A3(new_n303), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT68), .A3(new_n307), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n326), .B1(new_n332), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(new_n321), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n326), .A2(KEYINPUT28), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n321), .B(KEYINPUT69), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(new_n316), .A3(new_n308), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n323), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n239), .B(new_n325), .C1(new_n345), .C2(new_n349), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n346), .A2(new_n316), .A3(new_n308), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(new_n347), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n332), .A2(new_n343), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n310), .A2(new_n321), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT31), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT31), .ZN(new_n358));
  AOI211_X1 g172(.A(new_n358), .B(new_n355), .C1(new_n332), .C2(new_n343), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n353), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(G472), .A2(G902), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n350), .A2(G472), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT68), .B1(new_n342), .B2(new_n307), .ZN(new_n368));
  AOI211_X1 g182(.A(new_n331), .B(new_n309), .C1(new_n340), .C2(new_n341), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n356), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n358), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n354), .A2(KEYINPUT31), .A3(new_n356), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n352), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n367), .B1(new_n373), .B2(new_n362), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n254), .B1(new_n365), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G110), .B(G140), .ZN(new_n376));
  INV_X1    g190(.A(G227), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G953), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n376), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G104), .ZN(new_n385));
  INV_X1    g199(.A(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(G107), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n381), .A2(G107), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n384), .A2(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(G101), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n293), .B(new_n392), .C1(new_n296), .C2(new_n297), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n286), .A2(new_n287), .A3(new_n292), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n286), .A2(new_n287), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT1), .ZN(new_n396));
  OAI21_X1  g210(.A(G128), .B1(new_n294), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n393), .B1(new_n398), .B2(new_n392), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n334), .A2(KEYINPUT81), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT12), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(new_n404), .A3(new_n400), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n334), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT10), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n398), .B2(new_n392), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n382), .A2(new_n385), .A3(new_n387), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G101), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n416), .A3(G101), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n415), .A2(new_n336), .A3(new_n337), .A4(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n392), .A2(new_n411), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n298), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n410), .A2(new_n412), .A3(new_n418), .A4(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n380), .B1(new_n408), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n396), .B1(new_n280), .B2(new_n210), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n395), .B1(new_n423), .B2(new_n187), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n392), .B1(new_n424), .B2(new_n293), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n418), .B(new_n420), .C1(new_n425), .C2(KEYINPUT10), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n269), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n421), .A2(new_n427), .A3(new_n380), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT82), .B1(new_n422), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n334), .B(KEYINPUT80), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n407), .B2(new_n406), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n431), .B(new_n428), .C1(new_n434), .C2(new_n380), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n430), .A2(G469), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n239), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n421), .A2(new_n427), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n379), .ZN(new_n440));
  INV_X1    g254(.A(new_n407), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n404), .B1(new_n399), .B2(new_n400), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n421), .B(new_n380), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(G902), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n438), .B1(new_n444), .B2(new_n437), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n436), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT9), .B(G234), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT79), .ZN(new_n448));
  OAI21_X1  g262(.A(G221), .B1(new_n448), .B2(G902), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G210), .B1(G237), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G125), .B1(new_n283), .B2(new_n289), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n198), .B(new_n293), .C1(new_n296), .C2(new_n297), .ZN(new_n456));
  INV_X1    g270(.A(G224), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G953), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT7), .A4(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT86), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n455), .A2(new_n456), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(new_n458), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n306), .A2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g279(.A(G116), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n466), .A2(KEYINPUT5), .A3(G119), .ZN(new_n467));
  INV_X1    g281(.A(G113), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n465), .A2(new_n469), .B1(new_n305), .B2(new_n306), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n470), .B(KEYINPUT85), .C1(new_n471), .C2(new_n392), .ZN(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G122), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT8), .ZN(new_n474));
  INV_X1    g288(.A(new_n470), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n388), .A2(new_n391), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n392), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n479), .B2(KEYINPUT84), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n472), .B(new_n474), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n307), .A2(new_n415), .A3(new_n417), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n470), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n473), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n464), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n239), .B1(new_n461), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT83), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT6), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n482), .A2(new_n483), .ZN(new_n491));
  INV_X1    g305(.A(new_n473), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n492), .A3(new_n489), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n462), .A2(new_n458), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n494), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n454), .B1(new_n486), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n464), .A2(new_n481), .A3(new_n484), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n460), .B(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n494), .A2(new_n495), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n496), .A2(new_n497), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n506), .A3(new_n453), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n452), .B1(new_n499), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(G234), .A2(G237), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n509), .A2(G952), .A3(new_n224), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n509), .A2(G902), .A3(G953), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT21), .B(G898), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G113), .B(G122), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n381), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n317), .A2(new_n224), .A3(G214), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n277), .A3(new_n279), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n317), .A2(new_n224), .A3(G143), .A4(G214), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n299), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n207), .A2(new_n213), .B1(KEYINPUT17), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G131), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n299), .A3(new_n520), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n521), .A2(KEYINPUT18), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n220), .B1(new_n210), .B2(new_n208), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n299), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n529), .B(new_n530), .C1(new_n523), .C2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n517), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT89), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n528), .A2(new_n517), .A3(new_n533), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(G902), .B1(new_n534), .B2(KEYINPUT89), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G475), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n519), .A2(new_n299), .A3(new_n520), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT87), .B1(new_n542), .B2(new_n521), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT87), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n524), .A2(new_n544), .A3(new_n526), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n202), .A2(new_n203), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT19), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n208), .A2(KEYINPUT19), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n550), .A2(new_n219), .B1(G146), .B2(new_n209), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(new_n545), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT88), .A3(new_n533), .ZN(new_n553));
  INV_X1    g367(.A(new_n517), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT88), .B1(new_n552), .B2(new_n533), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n537), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n558));
  NOR2_X1   g372(.A1(G475), .A2(G902), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n541), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n448), .A2(new_n238), .A3(G953), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G116), .B(G122), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(new_n384), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n277), .A2(new_n279), .A3(G128), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n187), .A2(G143), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n256), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT13), .A4(G128), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(KEYINPUT91), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT65), .B(G143), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n575), .A2(KEYINPUT91), .A3(KEYINPUT13), .A4(G128), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n568), .A2(KEYINPUT90), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT90), .B1(new_n568), .B2(new_n577), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n574), .B(new_n576), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n571), .B1(new_n580), .B2(G134), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n568), .A2(new_n569), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G134), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n570), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n466), .A2(G122), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n384), .B1(new_n585), .B2(KEYINPUT14), .ZN(new_n586));
  INV_X1    g400(.A(new_n566), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n565), .B1(new_n581), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n568), .A2(new_n577), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT90), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n568), .A2(KEYINPUT90), .A3(new_n577), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n574), .A2(new_n576), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n256), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n564), .B(new_n592), .C1(new_n599), .C2(new_n571), .ZN(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n591), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G478), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT92), .B1(new_n602), .B2(KEYINPUT15), .ZN(new_n603));
  OR3_X1    g417(.A1(new_n602), .A2(KEYINPUT92), .A3(KEYINPUT15), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(new_n601), .B2(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n563), .A2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n450), .A2(new_n515), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n375), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  OAI21_X1  g424(.A(G472), .B1(new_n373), .B2(G902), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n446), .A2(new_n253), .A3(new_n449), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n371), .A2(new_n372), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n362), .B1(new_n615), .B2(new_n353), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI211_X1 g431(.A(KEYINPUT93), .B(G472), .C1(new_n373), .C2(G902), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n613), .A2(new_n614), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n360), .B2(new_n239), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n616), .B1(new_n623), .B2(KEYINPUT93), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n624), .A2(KEYINPUT94), .A3(new_n613), .A4(new_n614), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n591), .A2(new_n600), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n239), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(KEYINPUT96), .A3(new_n602), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n601), .B2(G478), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n600), .B2(KEYINPUT95), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n627), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n591), .B(new_n600), .C1(KEYINPUT95), .C2(new_n633), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n602), .A2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n562), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n515), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n626), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT97), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n643), .B(new_n645), .ZN(G6));
  INV_X1    g460(.A(new_n606), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n563), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n515), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n626), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT98), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  AND2_X1   g467(.A1(new_n624), .A2(new_n613), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n251), .A2(new_n249), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n250), .B1(new_n245), .B2(new_n246), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n240), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n233), .A2(new_n235), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n658), .B(new_n659), .Z(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n241), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR4_X1   g477(.A1(new_n450), .A2(new_n663), .A3(new_n607), .A4(new_n515), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n360), .A2(new_n364), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n310), .B1(new_n368), .B2(new_n369), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n349), .B1(new_n669), .B2(new_n322), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n325), .A2(new_n239), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n668), .B(new_n672), .C1(new_n616), .C2(new_n366), .ZN(new_n673));
  INV_X1    g487(.A(new_n450), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n486), .A2(new_n498), .A3(new_n454), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n453), .B1(new_n503), .B2(new_n506), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n451), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n663), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n510), .B1(new_n511), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n648), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n673), .A2(new_n674), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XOR2_X1   g497(.A(new_n680), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n674), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n499), .A2(new_n507), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n562), .A2(new_n647), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n689), .A2(new_n452), .A3(new_n662), .A4(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n347), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n311), .A2(new_n692), .A3(new_n313), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n370), .A2(KEYINPUT100), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n239), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT100), .B1(new_n370), .B2(new_n693), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n374), .A2(new_n668), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n686), .A2(new_n691), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n280), .ZN(G45));
  INV_X1    g515(.A(new_n680), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n562), .A2(new_n640), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n673), .A2(new_n674), .A3(new_n678), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT101), .B(G146), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G48));
  OAI21_X1  g521(.A(new_n380), .B1(new_n426), .B2(new_n432), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n407), .B2(new_n406), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n380), .B1(new_n421), .B2(new_n427), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n239), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n437), .B(new_n239), .C1(new_n709), .C2(new_n710), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n449), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n254), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n673), .A2(new_n642), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND3_X1  g532(.A1(new_n673), .A2(new_n649), .A3(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  NOR3_X1   g534(.A1(new_n607), .A2(new_n513), .A3(new_n714), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n673), .A2(new_n721), .A3(new_n678), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  OAI21_X1  g537(.A(KEYINPUT103), .B1(new_n690), .B2(new_n677), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n508), .A2(new_n725), .A3(new_n562), .A4(new_n647), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n513), .B(new_n714), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n314), .A2(new_n316), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n692), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n362), .B1(new_n615), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n623), .A2(new_n254), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(KEYINPUT102), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n623), .A2(new_n730), .A3(new_n733), .A4(new_n254), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n727), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NOR3_X1   g550(.A1(new_n623), .A2(new_n663), .A3(new_n730), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n703), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n714), .A2(new_n677), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n562), .A2(new_n640), .A3(KEYINPUT104), .A4(new_n702), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n737), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n730), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n611), .A3(new_n662), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT105), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NAND4_X1  g564(.A1(new_n499), .A2(new_n507), .A3(new_n451), .A4(new_n449), .ZN(new_n751));
  INV_X1    g565(.A(new_n438), .ZN(new_n752));
  OAI211_X1 g566(.A(G469), .B(new_n428), .C1(new_n434), .C2(new_n380), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n713), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n713), .A2(new_n753), .A3(KEYINPUT106), .A4(new_n752), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n751), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n739), .A3(new_n741), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n363), .B1(new_n373), .B2(new_n362), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n254), .B1(new_n365), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n762), .A3(KEYINPUT42), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  INV_X1    g578(.A(new_n364), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n672), .B1(new_n373), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n366), .B1(new_n360), .B2(new_n361), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n253), .B(new_n758), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n739), .A2(new_n741), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  INV_X1    g586(.A(new_n681), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n256), .ZN(G36));
  INV_X1    g589(.A(new_n654), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n563), .A2(new_n640), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n780));
  OAI22_X1  g594(.A1(new_n779), .A2(KEYINPUT108), .B1(new_n780), .B2(new_n777), .ZN(new_n781));
  INV_X1    g595(.A(new_n779), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n776), .B(new_n662), .C1(new_n781), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n687), .A2(new_n452), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n786), .ZN(new_n789));
  INV_X1    g603(.A(new_n449), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n428), .B1(new_n434), .B2(new_n380), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  OAI21_X1  g606(.A(G469), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n430), .A2(new_n435), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n793), .B1(new_n794), .B2(new_n792), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(new_n438), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n796), .A2(new_n797), .B1(new_n437), .B2(new_n444), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n790), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(new_n684), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n787), .A2(new_n788), .A3(new_n789), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  INV_X1    g617(.A(new_n673), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n254), .A3(new_n704), .A4(new_n788), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n800), .A2(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n800), .A2(KEYINPUT47), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(new_n201), .ZN(G42));
  NAND2_X1  g623(.A1(new_n712), .A2(new_n713), .ZN(new_n810));
  INV_X1    g624(.A(new_n510), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n810), .A2(new_n751), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n698), .A2(new_n813), .A3(new_n254), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT117), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n562), .A2(new_n640), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n812), .B1(new_n784), .B2(new_n781), .ZN(new_n818));
  OAI22_X1  g632(.A1(new_n815), .A2(new_n817), .B1(new_n746), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n810), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n790), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n806), .A2(new_n807), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n784), .A2(new_n781), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n811), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n732), .A2(new_n734), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n826), .A2(new_n827), .A3(new_n788), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n819), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n689), .A2(new_n452), .A3(new_n449), .A4(new_n820), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT115), .Z(new_n831));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(KEYINPUT50), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(new_n835), .A3(KEYINPUT51), .ZN(new_n836));
  INV_X1    g650(.A(G952), .ZN(new_n837));
  INV_X1    g651(.A(new_n762), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n818), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n840), .A2(KEYINPUT48), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n837), .B(G953), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(KEYINPUT48), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n839), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n815), .A2(new_n641), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n826), .A2(new_n827), .A3(new_n740), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n842), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n836), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT51), .B1(new_n829), .B2(new_n835), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n716), .A2(new_n719), .A3(new_n722), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n771), .A2(new_n851), .A3(new_n735), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n606), .A2(KEYINPUT110), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT110), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n605), .B(new_n854), .C1(new_n601), .C2(new_n603), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n563), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n515), .B1(new_n857), .B2(new_n641), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n621), .A2(new_n625), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n654), .A2(new_n664), .B1(new_n375), .B2(new_n608), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n768), .A2(new_n773), .B1(new_n759), .B2(new_n746), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n673), .A2(new_n674), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n856), .A2(new_n562), .A3(new_n680), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(new_n662), .A3(new_n788), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n866), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n673), .A3(KEYINPUT111), .A4(new_n674), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n862), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n852), .A2(new_n861), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n743), .B1(new_n737), .B2(new_n742), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT105), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n657), .A2(new_n449), .A3(new_n661), .A4(new_n702), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n756), .B2(new_n757), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n724), .A2(new_n726), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n698), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n682), .A2(new_n705), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT52), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n874), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n682), .A2(new_n705), .A3(new_n878), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT52), .B1(new_n882), .B2(new_n749), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n871), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g699(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT53), .B1(new_n871), .B2(new_n884), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(KEYINPUT54), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT113), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n891), .B(new_n862), .C1(new_n867), .C2(new_n869), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n852), .A3(new_n861), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n890), .B1(new_n893), .B2(new_n884), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n886), .B1(new_n871), .B2(new_n884), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n870), .A2(KEYINPUT53), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n771), .A2(new_n735), .A3(new_n851), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n880), .B1(new_n874), .B2(new_n879), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n882), .A2(KEYINPUT52), .A3(new_n749), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(new_n901), .A3(KEYINPUT113), .A4(new_n861), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n894), .A2(new_n895), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n889), .A2(new_n904), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n850), .A2(new_n905), .B1(G952), .B2(G953), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n777), .A2(new_n452), .A3(new_n790), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n253), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT109), .Z(new_n910));
  OAI21_X1  g724(.A(new_n689), .B1(new_n810), .B2(KEYINPUT49), .ZN(new_n911));
  OR3_X1    g725(.A1(new_n910), .A2(new_n698), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT119), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n906), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(G75));
  NOR2_X1   g731(.A1(new_n224), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n894), .A2(new_n895), .A3(new_n902), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n920), .A2(G902), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT56), .B1(new_n921), .B2(G210), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n504), .B(new_n505), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT55), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n922), .B2(new_n925), .ZN(G51));
  NOR2_X1   g741(.A1(new_n709), .A2(new_n710), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n920), .A2(KEYINPUT54), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n904), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n438), .B(KEYINPUT57), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n920), .A2(G902), .A3(new_n795), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT120), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n920), .A2(new_n935), .A3(G902), .A4(new_n795), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n919), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g754(.A(KEYINPUT121), .B(new_n919), .C1(new_n932), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G54));
  AND2_X1   g756(.A1(KEYINPUT58), .A2(G475), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n921), .A2(KEYINPUT122), .A3(new_n557), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n920), .A2(G902), .A3(new_n943), .ZN(new_n945));
  INV_X1    g759(.A(new_n557), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n918), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT122), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n945), .B2(new_n946), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n944), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G60));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT59), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n930), .A2(new_n637), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n637), .B1(new_n905), .B2(new_n955), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n918), .ZN(G63));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT60), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n920), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n660), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n919), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI22_X1  g777(.A1(new_n920), .A2(new_n960), .B1(new_n237), .B2(new_n231), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n919), .C1(new_n961), .C2(new_n962), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT61), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n965), .B(new_n968), .ZN(G66));
  INV_X1    g783(.A(new_n512), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n224), .B1(new_n970), .B2(G224), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n861), .A2(new_n735), .A3(new_n851), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n224), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n494), .B(new_n495), .C1(G898), .C2(new_n224), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n973), .B(new_n974), .Z(G69));
  XOR2_X1   g789(.A(new_n342), .B(new_n550), .Z(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT125), .Z(new_n977));
  INV_X1    g791(.A(new_n788), .ZN(new_n978));
  AOI211_X1 g792(.A(new_n978), .B(new_n685), .C1(new_n641), .C2(new_n857), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n808), .B1(new_n375), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n682), .A2(new_n705), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n700), .A2(new_n981), .A3(new_n749), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n980), .A2(new_n802), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n977), .B1(new_n985), .B2(new_n224), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n224), .A2(G900), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n801), .A2(new_n877), .A3(new_n762), .ZN(new_n988));
  INV_X1    g802(.A(new_n774), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n988), .A2(new_n771), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n981), .A2(new_n749), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n808), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n990), .A2(new_n992), .A3(new_n802), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n987), .B1(new_n993), .B2(new_n224), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n976), .B1(new_n994), .B2(new_n995), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n986), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n377), .B2(new_n679), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n985), .B2(new_n972), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n321), .A3(new_n669), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n370), .B1(new_n344), .B2(new_n321), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n887), .A2(new_n888), .A3(new_n1002), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n993), .A2(new_n972), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1002), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n344), .A2(new_n322), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n919), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n1012), .A2(KEYINPUT127), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(KEYINPUT127), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1007), .B1(new_n1013), .B2(new_n1014), .ZN(G57));
endmodule


