//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n202), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n207), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT65), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n227), .A2(G1), .A3(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G20), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  OAI22_X1  g0031(.A1(new_n222), .A2(KEYINPUT1), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n210), .A2(new_n224), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n218), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND2_X1  g0049(.A1(new_n203), .A2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n250), .B1(new_n251), .B2(new_n253), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n226), .A2(new_n228), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT69), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT69), .A4(new_n258), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n202), .B1(new_n265), .B2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n202), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n270), .A2(KEYINPUT70), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT70), .B1(new_n270), .B2(new_n271), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n264), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  INV_X1    g0076(.A(new_n225), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n282), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n277), .A2(new_n278), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n286), .B2(new_n212), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT68), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT3), .ZN(new_n292));
  INV_X1    g0092(.A(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT68), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(G222), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(G223), .A3(G1698), .ZN(new_n300));
  INV_X1    g0100(.A(G77), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n299), .B(new_n300), .C1(new_n301), .C2(new_n297), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n226), .A2(new_n228), .B1(G33), .B2(G41), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n287), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G169), .B2(new_n304), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n275), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n274), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(G190), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G200), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT10), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n274), .B(KEYINPUT9), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(KEYINPUT71), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n304), .B2(new_n313), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n318), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n308), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n283), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n282), .B1(new_n277), .B2(new_n278), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(G238), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n290), .B1(new_n288), .B2(new_n289), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G226), .A2(G1698), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n218), .B2(G1698), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n294), .A2(KEYINPUT68), .A3(new_n295), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT72), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G97), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n303), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n333), .B2(new_n335), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n327), .B(new_n328), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n333), .A2(new_n335), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT72), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(new_n303), .A3(new_n336), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n328), .B1(new_n343), .B2(new_n327), .ZN(new_n344));
  OAI21_X1  g0144(.A(G169), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT14), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n327), .B1(new_n337), .B2(new_n338), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(G179), .A3(new_n339), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(G169), .C1(new_n340), .C2(new_n344), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n346), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G68), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n301), .B2(new_n255), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n263), .A2(KEYINPUT11), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n267), .A2(new_n353), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT12), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n226), .A2(new_n228), .A3(new_n266), .A4(new_n258), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n265), .A2(G20), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G68), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n356), .B(new_n358), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT11), .B1(new_n263), .B2(new_n355), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n352), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(G200), .B1(new_n340), .B2(new_n344), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n348), .A2(G190), .A3(new_n339), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n372));
  INV_X1    g0172(.A(new_n303), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n293), .A2(new_n213), .ZN(new_n374));
  OAI211_X1 g0174(.A(G223), .B(new_n298), .C1(new_n288), .C2(new_n289), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G226), .A2(G1698), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n298), .A2(KEYINPUT74), .A3(G223), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n378), .A2(new_n379), .B1(new_n294), .B2(new_n295), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n373), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n283), .B1(new_n286), .B2(new_n218), .ZN(new_n383));
  OAI21_X1  g0183(.A(G169), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n326), .A2(G232), .B1(new_n279), .B2(new_n282), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n294), .A2(new_n295), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n298), .A2(G223), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT74), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n388), .A2(new_n380), .A3(new_n374), .ZN(new_n389));
  OAI211_X1 g0189(.A(G179), .B(new_n385), .C1(new_n389), .C2(new_n373), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT75), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n384), .A2(new_n390), .A3(KEYINPUT75), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n256), .B1(new_n265), .B2(G20), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n268), .A2(new_n395), .B1(new_n267), .B2(new_n256), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n386), .B2(G20), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n294), .A2(KEYINPUT7), .A3(new_n254), .A4(new_n295), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n353), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n217), .A2(new_n353), .ZN(new_n402));
  OAI21_X1  g0202(.A(G20), .B1(new_n402), .B2(new_n201), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n252), .A2(G159), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT16), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n398), .B1(new_n297), .B2(G20), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n288), .A2(new_n289), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT73), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT7), .A4(new_n254), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n353), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n403), .A2(new_n404), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n406), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n397), .B1(new_n417), .B2(new_n259), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n372), .B1(new_n394), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(G20), .B1(new_n329), .B2(new_n332), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n408), .B(new_n411), .C1(new_n420), .C2(KEYINPUT7), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n416), .B1(new_n421), .B2(G68), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT7), .B1(new_n409), .B2(new_n254), .ZN(new_n423));
  INV_X1    g0223(.A(new_n400), .ZN(new_n424));
  OAI21_X1  g0224(.A(G68), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n415), .B1(new_n425), .B2(new_n414), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n259), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n377), .A2(new_n381), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n303), .ZN(new_n429));
  INV_X1    g0229(.A(G190), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n385), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n313), .B1(new_n382), .B2(new_n383), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n427), .A2(new_n396), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n384), .A2(new_n390), .A3(KEYINPUT75), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(new_n391), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n427), .A2(new_n396), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT76), .B(KEYINPUT18), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n433), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n419), .A2(new_n436), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n256), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n444), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n445));
  XOR2_X1   g0245(.A(KEYINPUT15), .B(G87), .Z(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n255), .B2(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n448), .A2(new_n259), .B1(new_n301), .B2(new_n267), .ZN(new_n449));
  INV_X1    g0249(.A(new_n359), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G77), .A3(new_n360), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n329), .A2(new_n332), .ZN(new_n453));
  INV_X1    g0253(.A(G107), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n373), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  MUX2_X1   g0255(.A(G232), .B(G238), .S(G1698), .Z(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n325), .B1(G244), .B2(new_n326), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n452), .B1(new_n460), .B2(G190), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n313), .B2(new_n460), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n305), .ZN(new_n463));
  INV_X1    g0263(.A(G169), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n459), .A2(new_n464), .B1(new_n449), .B2(new_n451), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n443), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n324), .A2(new_n370), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n386), .A2(new_n254), .A3(G68), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT19), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n255), .B2(new_n219), .ZN(new_n473));
  NAND3_X1  g0273(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT80), .A3(new_n254), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G97), .A2(G107), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n213), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT80), .B1(new_n474), .B2(new_n254), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n471), .B(new_n473), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT81), .ZN(new_n481));
  INV_X1    g0281(.A(new_n479), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n477), .A3(new_n475), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT81), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n471), .A4(new_n473), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n259), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n447), .A2(new_n267), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n265), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n261), .A2(new_n262), .A3(new_n266), .A4(new_n488), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n489), .A2(new_n213), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n486), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G116), .ZN(new_n492));
  INV_X1    g0292(.A(G244), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G1698), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(G238), .B2(G1698), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n495), .B2(new_n409), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n303), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n281), .A2(G1), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n214), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n279), .A2(new_n498), .B1(new_n499), .B2(new_n285), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n313), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G190), .B2(new_n501), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n486), .B(new_n487), .C1(new_n447), .C2(new_n489), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n497), .A2(new_n500), .A3(new_n305), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n464), .B2(new_n501), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n491), .A2(new_n503), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n265), .A2(G45), .ZN(new_n509));
  OR2_X1    g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  NAND2_X1  g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n279), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT5), .B(G41), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n498), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n285), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n513), .B1(new_n516), .B2(new_n220), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n493), .A2(G1698), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n288), .B2(new_n289), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n493), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n329), .A2(new_n332), .A3(new_n298), .A4(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n297), .A2(KEYINPUT78), .A3(G250), .A4(G1698), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n329), .A2(new_n332), .A3(G250), .A4(G1698), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT78), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n517), .B1(new_n531), .B2(new_n303), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n305), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT77), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n489), .A2(G97), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n267), .A2(G97), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n534), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AOI211_X1 g0338(.A(KEYINPUT77), .B(new_n536), .C1(new_n489), .C2(G97), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT6), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n540), .A2(new_n219), .A3(G107), .ZN(new_n541));
  XNOR2_X1  g0341(.A(G97), .B(G107), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n543), .A2(new_n254), .B1(new_n301), .B2(new_n253), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n421), .B2(G107), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n226), .A2(new_n228), .A3(new_n258), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n538), .A2(new_n539), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n533), .B(new_n547), .C1(G169), .C2(new_n532), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n530), .A2(new_n525), .A3(new_n523), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n528), .A2(new_n529), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n303), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n517), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT79), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(G200), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT79), .B1(new_n532), .B2(new_n313), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n551), .A2(G190), .A3(new_n552), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n545), .A2(new_n546), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n539), .C2(new_n538), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n508), .B(new_n548), .C1(new_n557), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT82), .ZN(new_n562));
  INV_X1    g0362(.A(new_n547), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n555), .A3(new_n556), .A4(new_n558), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(new_n508), .A4(new_n548), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n220), .A2(G1698), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G250), .B2(G1698), .ZN(new_n569));
  INV_X1    g0369(.A(G294), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n569), .A2(new_n409), .B1(new_n293), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n303), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n514), .A2(new_n498), .B1(new_n277), .B2(new_n278), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G264), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n513), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(G179), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n464), .B2(new_n575), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n254), .B(G87), .C1(new_n288), .C2(new_n289), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  OR3_X1    g0379(.A1(new_n213), .A2(KEYINPUT22), .A3(G20), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n579), .B1(new_n453), .B2(new_n580), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n254), .A2(KEYINPUT23), .A3(G107), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT88), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT23), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n454), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n454), .A3(G20), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n586), .A2(KEYINPUT88), .B1(new_n587), .B2(G20), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n585), .A2(new_n588), .A3(KEYINPUT89), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT89), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n492), .A2(new_n584), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n582), .A2(new_n583), .B1(new_n591), .B2(new_n254), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n586), .A2(KEYINPUT88), .B1(KEYINPUT23), .B2(G107), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n581), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  XOR2_X1   g0395(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT89), .B1(new_n585), .B2(new_n588), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n592), .A2(new_n590), .A3(new_n593), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n596), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n581), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n546), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n489), .A2(new_n454), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n267), .A2(new_n454), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n605), .B(KEYINPUT25), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n577), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n600), .A2(new_n581), .A3(new_n601), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n601), .B1(new_n600), .B2(new_n581), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n259), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n575), .A2(G200), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n575), .A2(new_n430), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n615), .A3(new_n607), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  INV_X1    g0418(.A(G303), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n329), .B2(new_n332), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n220), .A2(new_n298), .ZN(new_n621));
  INV_X1    g0421(.A(G264), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G1698), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n621), .B(new_n623), .C1(new_n288), .C2(new_n289), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n303), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n573), .A2(G270), .B1(new_n279), .B2(new_n512), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n464), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT20), .ZN(new_n629));
  INV_X1    g0429(.A(G116), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(G20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n518), .A2(new_n254), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n219), .A2(G33), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n629), .B1(new_n546), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT85), .ZN(new_n636));
  AOI21_X1  g0436(.A(G20), .B1(G33), .B2(G283), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n293), .A2(G97), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n637), .A2(new_n638), .B1(G20), .B2(new_n630), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n259), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT85), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n629), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n639), .A2(new_n259), .A3(KEYINPUT20), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT84), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT84), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n639), .A2(new_n259), .A3(new_n645), .A4(KEYINPUT20), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n636), .A2(new_n642), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n488), .A2(G116), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT83), .B1(new_n359), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n359), .A2(KEYINPUT83), .A3(new_n648), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n650), .A2(new_n651), .B1(G116), .B2(new_n266), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n628), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(G303), .B1(new_n291), .B2(new_n296), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n373), .B1(new_n654), .B2(new_n624), .ZN(new_n655));
  INV_X1    g0455(.A(G270), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n513), .B1(new_n516), .B2(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(KEYINPUT21), .B(G169), .C1(new_n655), .C2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n626), .A2(G179), .A3(new_n627), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n644), .A2(new_n646), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n641), .B1(new_n640), .B2(new_n629), .ZN(new_n662));
  AOI211_X1 g0462(.A(KEYINPUT85), .B(KEYINPUT20), .C1(new_n639), .C2(new_n259), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n651), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n665), .A2(new_n649), .B1(new_n630), .B2(new_n267), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n618), .A2(new_n653), .B1(new_n660), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n313), .B1(new_n626), .B2(new_n627), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n626), .A2(G190), .A3(new_n627), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n672), .A2(new_n667), .A3(KEYINPUT86), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT86), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n626), .A2(G190), .A3(new_n627), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n669), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n647), .A2(new_n652), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n668), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  NOR4_X1   g0479(.A1(new_n470), .A2(new_n567), .A3(new_n617), .A4(new_n679), .ZN(G372));
  NAND2_X1  g0480(.A1(new_n384), .A2(new_n390), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n439), .A2(new_n371), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n371), .B1(new_n439), .B2(new_n681), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n466), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n352), .A2(new_n365), .B1(new_n369), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT90), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n434), .B(KEYINPUT17), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n686), .B2(new_n687), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n684), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n317), .A2(new_n323), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n308), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n504), .A2(new_n507), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT26), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n491), .A2(new_n503), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n694), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n698), .B2(new_n548), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n553), .A2(G179), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n532), .A2(G169), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(new_n508), .A3(KEYINPUT26), .A4(new_n547), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n695), .B1(new_n699), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n668), .A2(new_n609), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n564), .A2(new_n508), .A3(new_n548), .A4(new_n616), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n693), .B1(new_n470), .B2(new_n709), .ZN(G369));
  INV_X1    g0510(.A(new_n668), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n265), .A2(new_n254), .A3(G13), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n714), .A3(G213), .ZN(new_n715));
  INV_X1    g0515(.A(G343), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n677), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n679), .B2(new_n719), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n609), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n717), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n612), .A2(new_n607), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n717), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n609), .A3(new_n616), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n711), .A2(new_n718), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n617), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n609), .A2(new_n717), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(G399));
  INV_X1    g0535(.A(new_n208), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n476), .A2(new_n213), .A3(new_n630), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n737), .A2(new_n265), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n231), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n737), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT28), .Z(new_n742));
  OR2_X1    g0542(.A1(new_n707), .A2(new_n706), .ZN(new_n743));
  AOI211_X1 g0543(.A(KEYINPUT29), .B(new_n717), .C1(new_n743), .C2(new_n704), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n705), .A2(KEYINPUT92), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT92), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n668), .A2(new_n609), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n704), .B1(new_n707), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n745), .B1(new_n750), .B2(new_n718), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n744), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G330), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n572), .A2(new_n497), .A3(new_n500), .A4(new_n574), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n659), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(new_n551), .A3(new_n552), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT30), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n626), .A2(new_n627), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n575), .A2(new_n305), .A3(new_n501), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n553), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n532), .A2(KEYINPUT30), .A3(new_n755), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n758), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT31), .B1(new_n763), .B2(new_n717), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n717), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n764), .B1(KEYINPUT91), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT91), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n767), .B(KEYINPUT31), .C1(new_n763), .C2(new_n717), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n679), .A2(new_n617), .A3(new_n717), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n562), .A2(new_n770), .A3(new_n566), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n753), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n752), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n742), .B1(new_n775), .B2(G1), .ZN(G364));
  INV_X1    g0576(.A(G13), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n265), .B1(new_n778), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n737), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n721), .A2(G330), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n723), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n229), .B1(new_n254), .B2(G169), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT94), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT94), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n736), .A2(new_n386), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n231), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G45), .B2(new_n248), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n208), .A2(new_n297), .A3(G355), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G116), .B2(new_n208), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n792), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n781), .ZN(new_n799));
  INV_X1    g0599(.A(new_n791), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n721), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n254), .A2(new_n305), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT95), .ZN(new_n804));
  AOI21_X1  g0604(.A(G200), .B1(new_n803), .B2(KEYINPUT95), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(new_n430), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(G190), .A3(new_n805), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G311), .A2(new_n807), .B1(new_n809), .B2(G322), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n313), .A2(G179), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(G20), .A3(G190), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n453), .B1(new_n619), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT98), .Z(new_n815));
  NAND2_X1  g0615(.A1(new_n802), .A2(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n430), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G179), .A2(G200), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n254), .B1(new_n818), .B2(G190), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n817), .A2(G326), .B1(G294), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n816), .A2(G190), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(KEYINPUT33), .B(G317), .Z(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n430), .A2(G20), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT96), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n828), .A2(G179), .A3(G200), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G329), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n828), .A2(G179), .A3(new_n313), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G283), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n811), .A2(new_n815), .A3(new_n825), .A4(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT99), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(KEYINPUT99), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n829), .A2(G159), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT32), .Z(new_n840));
  AOI22_X1  g0640(.A1(G58), .A2(new_n809), .B1(new_n807), .B2(G77), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n822), .A2(G68), .B1(G97), .B2(new_n820), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT97), .Z(new_n843));
  INV_X1    g0643(.A(new_n813), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G87), .ZN(new_n845));
  INV_X1    g0645(.A(new_n817), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n297), .B(new_n845), .C1(new_n846), .C2(new_n202), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G107), .B2(new_n831), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n840), .A2(new_n841), .A3(new_n843), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n837), .A2(new_n838), .A3(new_n849), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n799), .B(new_n801), .C1(new_n788), .C2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n784), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G396));
  INV_X1    g0653(.A(new_n781), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n788), .A2(new_n789), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n301), .ZN(new_n856));
  INV_X1    g0656(.A(new_n788), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n453), .B1(new_n454), .B2(new_n813), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT101), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n831), .A2(G87), .ZN(new_n860));
  INV_X1    g0660(.A(new_n829), .ZN(new_n861));
  INV_X1    g0661(.A(G311), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n860), .B1(new_n219), .B2(new_n819), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n859), .B(new_n863), .C1(G294), .C2(new_n809), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G283), .A2(new_n822), .B1(new_n817), .B2(G303), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n630), .B2(new_n806), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT100), .Z(new_n867));
  AOI22_X1  g0667(.A1(G137), .A2(new_n817), .B1(new_n822), .B2(G150), .ZN(new_n868));
  INV_X1    g0668(.A(G159), .ZN(new_n869));
  INV_X1    g0669(.A(G143), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n868), .B1(new_n806), .B2(new_n869), .C1(new_n870), .C2(new_n808), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT34), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n386), .B1(new_n813), .B2(new_n202), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(G58), .B2(new_n820), .ZN(new_n875));
  INV_X1    g0675(.A(G132), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n875), .B1(new_n832), .B2(new_n353), .C1(new_n876), .C2(new_n861), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n871), .B2(new_n872), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n864), .A2(new_n867), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n452), .A2(new_n717), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n462), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n466), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n466), .A2(new_n717), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n856), .B1(new_n857), .B2(new_n879), .C1(new_n886), .C2(new_n790), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n709), .B2(new_n717), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n467), .A2(new_n717), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n743), .B2(new_n704), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(new_n773), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT102), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n773), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n854), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n887), .B1(new_n895), .B2(new_n897), .ZN(G384));
  OAI21_X1  g0698(.A(G77), .B1(new_n217), .B2(new_n353), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n899), .A2(new_n231), .B1(G50), .B2(new_n353), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(G1), .A3(new_n777), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT103), .ZN(new_n902));
  INV_X1    g0702(.A(new_n543), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n630), .B(new_n230), .C1(new_n903), .C2(KEYINPUT35), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(KEYINPUT35), .B2(new_n903), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT36), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n906), .B2(new_n905), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n469), .B1(new_n744), .B2(new_n751), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n909), .A2(new_n693), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n883), .B1(new_n708), .B2(new_n889), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n425), .B(new_n414), .C1(KEYINPUT105), .C2(KEYINPUT16), .ZN(new_n914));
  NOR2_X1   g0714(.A1(KEYINPUT105), .A2(KEYINPUT16), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n401), .B2(new_n405), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n914), .A2(new_n916), .A3(new_n263), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n917), .A2(new_n397), .ZN(new_n918));
  INV_X1    g0718(.A(new_n715), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND4_X1   g0720(.A1(new_n439), .A2(new_n392), .A3(new_n393), .A4(new_n440), .ZN(new_n921));
  INV_X1    g0721(.A(new_n372), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n438), .B2(new_n439), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n920), .B1(new_n924), .B2(new_n689), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n439), .A2(new_n392), .A3(new_n393), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n439), .A2(new_n919), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT37), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(new_n434), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n917), .A2(new_n397), .B1(new_n681), .B2(new_n919), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n434), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT37), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n913), .B1(new_n925), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n920), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n443), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(KEYINPUT38), .A3(new_n933), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n369), .A2(new_n346), .A3(new_n349), .A4(new_n351), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n364), .A2(new_n718), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT104), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n941), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n366), .A2(new_n369), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n940), .A2(KEYINPUT104), .A3(new_n941), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n912), .A2(new_n939), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT39), .ZN(new_n950));
  AOI221_X4 g0750(.A(new_n913), .B1(new_n929), .B2(new_n932), .C1(new_n443), .C2(new_n936), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n439), .A2(new_n681), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(new_n927), .A3(new_n434), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT37), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n929), .ZN(new_n955));
  INV_X1    g0755(.A(new_n681), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT18), .B1(new_n418), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n439), .A2(new_n371), .A3(new_n681), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n957), .A2(new_n442), .A3(new_n436), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n715), .B1(new_n427), .B2(new_n396), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT38), .B1(new_n955), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n950), .B1(new_n951), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n935), .A2(KEYINPUT39), .A3(new_n938), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n352), .A2(new_n365), .A3(new_n718), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n715), .B1(new_n682), .B2(new_n683), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n949), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n910), .B(new_n969), .Z(new_n970));
  INV_X1    g0770(.A(KEYINPUT106), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n765), .B1(new_n764), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n763), .A2(KEYINPUT106), .A3(KEYINPUT31), .A4(new_n717), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n771), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n948), .A2(new_n974), .A3(new_n886), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT40), .B1(new_n951), .B2(new_n962), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT107), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n972), .A2(new_n973), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n885), .B1(new_n978), .B2(new_n771), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT40), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n927), .B1(new_n684), .B2(new_n689), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n960), .B1(new_n418), .B2(new_n433), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT37), .B1(new_n438), .B2(new_n439), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n953), .A2(KEYINPUT37), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n913), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n980), .B1(new_n985), .B2(new_n938), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT107), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n979), .A2(new_n986), .A3(new_n987), .A4(new_n948), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n939), .A2(new_n886), .A3(new_n948), .A4(new_n974), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n977), .A2(new_n988), .B1(new_n980), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n469), .A2(new_n974), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n753), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n990), .B2(new_n991), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n970), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n265), .B2(new_n778), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n970), .A2(new_n993), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n908), .B1(new_n995), .B2(new_n996), .ZN(G367));
  OAI211_X1 g0797(.A(new_n564), .B(new_n548), .C1(new_n563), .C2(new_n718), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n548), .B2(new_n718), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n999), .A2(KEYINPUT109), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(KEYINPUT109), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT108), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1003), .A2(new_n1004), .A3(new_n723), .A4(new_n729), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT108), .B1(new_n1002), .B2(new_n730), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n491), .A2(new_n718), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n695), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n698), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1007), .B(new_n1011), .Z(new_n1012));
  INV_X1    g0812(.A(new_n732), .ZN(new_n1013));
  OR3_X1    g0813(.A1(new_n1002), .A2(KEYINPUT42), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(KEYINPUT42), .B1(new_n1002), .B2(new_n1013), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1003), .A2(new_n724), .B1(new_n547), .B2(new_n702), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1014), .B(new_n1015), .C1(new_n1016), .C2(new_n717), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n737), .B(KEYINPUT41), .Z(new_n1022));
  OR3_X1    g0822(.A1(new_n1000), .A2(new_n1001), .A3(new_n734), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT44), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n734), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT45), .Z(new_n1027));
  AOI21_X1  g0827(.A(new_n730), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n731), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1013), .B1(new_n729), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(new_n722), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n774), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1025), .A2(new_n1027), .A3(new_n730), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1029), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1022), .B1(new_n1035), .B2(new_n775), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1020), .B(new_n1021), .C1(new_n1036), .C2(new_n780), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n792), .B1(new_n208), .B2(new_n447), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n241), .A2(new_n736), .A3(new_n386), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n781), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n409), .B1(new_n823), .B2(new_n570), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n846), .A2(new_n862), .B1(new_n819), .B2(new_n454), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(G303), .C2(new_n809), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n833), .B2(new_n806), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n844), .A2(G116), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT46), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n831), .A2(G97), .ZN(new_n1047));
  INV_X1    g0847(.A(G317), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1046), .B(new_n1047), .C1(new_n1048), .C2(new_n861), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n819), .A2(new_n353), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n817), .B2(G143), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n808), .B2(new_n251), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT110), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(KEYINPUT110), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT111), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n807), .A2(G50), .B1(new_n822), .B2(G159), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1053), .B(new_n1054), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1055), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n831), .A2(G77), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n829), .A2(G137), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n453), .B1(G58), .B2(new_n844), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1044), .A2(new_n1049), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n857), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1040), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n800), .B2(new_n1010), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1037), .A2(new_n1068), .ZN(G387));
  INV_X1    g0869(.A(new_n1033), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n774), .A2(new_n1032), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n737), .A3(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n844), .A2(G294), .B1(new_n820), .B2(G283), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G311), .A2(new_n822), .B1(new_n817), .B2(G322), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n806), .B2(new_n619), .C1(new_n1048), .C2(new_n808), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT115), .Z(new_n1076));
  OAI21_X1  g0876(.A(new_n1073), .B1(new_n1076), .B2(KEYINPUT48), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(KEYINPUT48), .B2(new_n1076), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT49), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n386), .B1(new_n829), .B2(G326), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n630), .B2(new_n832), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n813), .A2(new_n301), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n409), .B(new_n1083), .C1(G159), .C2(new_n817), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n820), .A2(new_n446), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n256), .C2(new_n823), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1047), .B1(new_n861), .B2(new_n251), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n202), .A2(new_n808), .B1(new_n806), .B2(new_n353), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n788), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1091));
  NOR3_X1   g0891(.A1(new_n1091), .A2(G50), .A3(new_n256), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n281), .B1(new_n353), .B2(new_n301), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1092), .A2(new_n738), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(G50), .B2(new_n256), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n736), .B(new_n386), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n281), .B2(new_n237), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n208), .A2(new_n297), .A3(new_n738), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(G107), .C2(new_n208), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(KEYINPUT114), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n792), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1100), .B2(KEYINPUT114), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n854), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1090), .B(new_n1104), .C1(new_n729), .C2(new_n800), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1072), .B(new_n1105), .C1(new_n779), .C2(new_n1032), .ZN(G393));
  INV_X1    g0906(.A(new_n1034), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1070), .B1(new_n1107), .B2(new_n1028), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1035), .A2(new_n1108), .A3(new_n737), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1002), .A2(new_n791), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT116), .Z(new_n1111));
  NAND2_X1  g0911(.A1(new_n793), .A2(new_n245), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n219), .B2(new_n208), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n808), .A2(new_n869), .B1(new_n251), .B2(new_n846), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT51), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n409), .B1(new_n844), .B2(G68), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n820), .A2(G77), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n823), .C2(new_n202), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n860), .B1(new_n861), .B2(new_n870), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(new_n444), .C2(new_n807), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n822), .A2(G303), .B1(G116), .B2(new_n820), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n453), .C1(new_n833), .C2(new_n813), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n829), .A2(G322), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n832), .B2(new_n454), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(G294), .C2(new_n807), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n808), .A2(new_n862), .B1(new_n1048), .B2(new_n846), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT52), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1115), .A2(new_n1120), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n781), .B1(new_n1102), .B2(new_n1113), .C1(new_n1128), .C2(new_n857), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1111), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1107), .A2(new_n1028), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n780), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1109), .A2(new_n1132), .ZN(G390));
  AOI21_X1  g0933(.A(new_n948), .B1(new_n772), .B2(new_n886), .ZN(new_n1134));
  AND4_X1   g0934(.A1(G330), .A2(new_n948), .A3(new_n974), .A4(new_n886), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n912), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n772), .A2(new_n886), .A3(new_n948), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n974), .A2(G330), .A3(new_n886), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n948), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n750), .A2(new_n718), .A3(new_n882), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1141), .A2(new_n884), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1136), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n469), .A2(G330), .A3(new_n974), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n909), .A2(new_n1145), .A3(new_n693), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n965), .B1(new_n951), .B2(new_n962), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1142), .B2(new_n1139), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n965), .B1(new_n911), .B2(new_n1139), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n963), .A2(new_n964), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1150), .A2(new_n1153), .A3(new_n1137), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n948), .B1(new_n891), .B2(new_n883), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1155), .A2(new_n965), .B1(new_n963), .B2(new_n964), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1141), .A2(new_n884), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1148), .B1(new_n1157), .B2(new_n948), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1135), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1147), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1144), .A2(new_n1154), .A3(new_n1159), .A4(new_n1146), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n737), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1154), .A2(new_n1159), .A3(new_n780), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n855), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n781), .B1(new_n1165), .B2(new_n444), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n832), .A2(new_n202), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n844), .A2(G150), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(G125), .C2(new_n829), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n817), .A2(G128), .B1(G159), .B2(new_n820), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n453), .B1(new_n822), .B2(G137), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT54), .B(G143), .Z(new_n1173));
  NAND2_X1  g0973(.A1(new_n807), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1170), .B(new_n1175), .C1(new_n876), .C2(new_n808), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n806), .A2(new_n219), .B1(new_n454), .B2(new_n823), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT117), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n817), .A2(G283), .ZN(new_n1181));
  AND4_X1   g0981(.A1(new_n453), .A2(new_n1181), .A3(new_n845), .A4(new_n1117), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G68), .A2(new_n831), .B1(new_n829), .B2(G294), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n809), .A2(G116), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1176), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1166), .B1(new_n1186), .B2(new_n788), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1152), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n790), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1163), .A2(new_n1164), .A3(new_n1189), .ZN(G378));
  NAND2_X1  g0990(.A1(new_n977), .A2(new_n988), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n753), .B1(new_n989), .B2(new_n980), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT10), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n318), .B2(new_n315), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n322), .A2(new_n319), .A3(new_n321), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n310), .A2(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1194), .A2(new_n1196), .B1(new_n275), .B2(new_n307), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n274), .A2(new_n919), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n324), .A2(new_n1198), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1191), .A2(new_n1192), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1208), .A2(new_n1209), .A3(new_n969), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n969), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1207), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1191), .A2(new_n1192), .A3(new_n1207), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1211), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n780), .B1(new_n1210), .B2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1207), .A2(new_n790), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n844), .A2(new_n1173), .ZN(new_n1219));
  INV_X1    g1019(.A(G128), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1219), .B1(new_n1220), .B2(new_n808), .C1(new_n823), .C2(new_n876), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G137), .B2(new_n807), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n817), .A2(G125), .B1(G150), .B2(new_n820), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT118), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n829), .A2(G124), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(G33), .A2(G41), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(new_n832), .C2(new_n869), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n823), .A2(new_n219), .B1(new_n846), .B2(new_n630), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n409), .A2(new_n280), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1232), .A2(new_n1050), .A3(new_n1083), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n829), .A2(G283), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n831), .A2(G58), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G107), .A2(new_n809), .B1(new_n807), .B2(new_n446), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT58), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1229), .A2(G50), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1238), .A2(new_n1239), .B1(new_n1233), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1239), .B2(new_n1238), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n788), .B1(new_n1231), .B2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n781), .C1(G50), .C2(new_n1165), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1218), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT119), .B1(new_n1217), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n969), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1214), .A2(new_n1211), .A3(new_n1215), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n779), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT119), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n1245), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1247), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT57), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1162), .B2(new_n1146), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT120), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1162), .A2(new_n1146), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1210), .B2(new_n1216), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1255), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1254), .A2(new_n1256), .A3(KEYINPUT120), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1259), .A2(new_n1262), .A3(new_n737), .A4(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1253), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(G375));
  INV_X1    g1066(.A(new_n1144), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1146), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1022), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n1147), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1139), .A2(new_n789), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n781), .B1(new_n1165), .B2(G68), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n829), .A2(G128), .B1(G159), .B2(new_n844), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT123), .Z(new_n1275));
  AOI22_X1  g1075(.A1(G132), .A2(new_n817), .B1(new_n822), .B2(new_n1173), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n409), .B1(new_n820), .B2(G50), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1236), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(G137), .A2(new_n809), .B1(new_n807), .B2(G150), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1059), .A2(new_n453), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT121), .Z(new_n1282));
  AOI22_X1  g1082(.A1(new_n817), .A2(G294), .B1(new_n844), .B2(G97), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n630), .B2(new_n823), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(G303), .B2(new_n829), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1282), .B(new_n1285), .C1(new_n454), .C2(new_n806), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1085), .B1(new_n808), .B2(new_n833), .ZN(new_n1287));
  XOR2_X1   g1087(.A(new_n1287), .B(KEYINPUT122), .Z(new_n1288));
  OAI21_X1  g1088(.A(new_n1280), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1273), .B1(new_n1289), .B2(new_n788), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1144), .A2(new_n780), .B1(new_n1272), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1271), .A2(new_n1291), .ZN(G381));
  NOR3_X1   g1092(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1293), .B(KEYINPUT124), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1294), .A2(G390), .A3(G381), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(G387), .A2(G378), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n1265), .A3(new_n1296), .ZN(G407));
  INV_X1    g1097(.A(G378), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n716), .A2(G213), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1265), .A2(new_n1298), .A3(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(G407), .A2(G213), .A3(new_n1301), .ZN(G409));
  NAND2_X1  g1102(.A1(new_n1147), .A2(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1269), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1267), .A2(KEYINPUT60), .A3(new_n1268), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n737), .A3(new_n1305), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1306), .A2(G384), .A3(new_n1291), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G384), .B1(new_n1306), .B2(new_n1291), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1300), .A2(G2897), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1309), .B(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1253), .A2(new_n1264), .A3(G378), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1217), .B(new_n1246), .C1(new_n1261), .C2(new_n1022), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1298), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1300), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT63), .B1(new_n1315), .B2(new_n1309), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(G393), .B(new_n852), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1037), .A2(new_n1068), .A3(G390), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G390), .B1(new_n1037), .B2(new_n1068), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1319), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(G390), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G387), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1037), .A2(new_n1068), .A3(G390), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1318), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1322), .A2(new_n1326), .ZN(new_n1327));
  NOR4_X1   g1127(.A1(new_n1316), .A2(new_n1317), .A3(new_n1327), .A4(KEYINPUT61), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT125), .B1(new_n1329), .B2(new_n1299), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT125), .ZN(new_n1331));
  AOI211_X1 g1131(.A(new_n1331), .B(new_n1300), .C1(new_n1312), .C2(new_n1314), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1333), .A2(KEYINPUT63), .A3(new_n1309), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1328), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1311), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1330), .B2(new_n1332), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1333), .A2(KEYINPUT62), .A3(new_n1309), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT126), .ZN(new_n1341));
  AOI211_X1 g1141(.A(new_n1341), .B(KEYINPUT62), .C1(new_n1315), .C2(new_n1309), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1329), .A2(new_n1299), .A3(new_n1309), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT62), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT126), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1339), .B1(new_n1340), .B2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1327), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1335), .B1(new_n1347), .B2(new_n1348), .ZN(G405));
  NOR2_X1   g1149(.A1(new_n1265), .A2(G378), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1312), .ZN(new_n1351));
  OR3_X1    g1151(.A1(new_n1350), .A2(new_n1351), .A3(new_n1309), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1309), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT127), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1352), .B(new_n1353), .C1(new_n1354), .C2(new_n1327), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1348), .A2(KEYINPUT127), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1355), .B(new_n1356), .ZN(G402));
endmodule


