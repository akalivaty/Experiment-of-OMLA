//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n191));
  INV_X1    g005(.A(G110), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n190), .A2(new_n191), .A3(new_n192), .A4(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n188), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT24), .B(G110), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n195), .A2(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(G125), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(G146), .B(new_n204), .C1(new_n208), .C2(new_n202), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT73), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n200), .A2(KEYINPUT16), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G146), .A4(new_n204), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n201), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT74), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n201), .A2(new_n210), .A3(KEYINPUT74), .A4(new_n213), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n204), .B1(new_n208), .B2(new_n202), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n199), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT72), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(new_n209), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(KEYINPUT72), .A3(new_n199), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n196), .A2(new_n197), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n190), .A2(new_n191), .A3(new_n194), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(G110), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n216), .A2(new_n217), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G953), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  XOR2_X1   g043(.A(new_n229), .B(KEYINPUT75), .Z(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G137), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n216), .A2(new_n234), .A3(new_n226), .A4(new_n217), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n236), .A2(new_n237), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(G217), .A2(G902), .ZN(new_n241));
  INV_X1    g055(.A(G217), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G234), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(KEYINPUT71), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT25), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n236), .A2(new_n239), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n244), .A2(G902), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n245), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n252), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  INV_X1    g073(.A(G137), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .A4(G134), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  OAI22_X1  g076(.A1(new_n262), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n260), .B2(G134), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G131), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n260), .A2(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n262), .A2(G137), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n266), .B1(new_n263), .B2(new_n261), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n272), .B1(new_n277), .B2(new_n268), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n199), .A2(G143), .ZN(new_n280));
  INV_X1    g094(.A(G143), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n199), .A2(G143), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n283), .A2(new_n187), .B1(KEYINPUT1), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G143), .B(G146), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT66), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AND4_X1   g102(.A1(KEYINPUT66), .A2(new_n287), .A3(new_n280), .A4(new_n282), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n276), .A2(new_n279), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT0), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n286), .B1(new_n292), .B2(new_n187), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT0), .B(G128), .Z(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n286), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n264), .A2(new_n268), .A3(new_n267), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n268), .B1(new_n264), .B2(new_n267), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n193), .A2(G116), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G119), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT2), .B(G113), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n304), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT67), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n290), .A2(new_n311), .A3(new_n278), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(new_n290), .B2(new_n278), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n308), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n298), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n310), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n281), .A2(KEYINPUT1), .A3(G146), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n318), .B1(new_n286), .B2(G128), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n287), .A2(new_n280), .A3(new_n282), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n286), .A2(KEYINPUT66), .A3(new_n287), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n319), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT67), .B1(new_n324), .B2(new_n274), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n290), .A2(new_n311), .A3(new_n278), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n298), .A2(new_n315), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n327), .A2(KEYINPUT68), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n309), .B1(new_n317), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT28), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n290), .A2(new_n278), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT28), .B1(new_n316), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n257), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT31), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT70), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n337), .B(new_n257), .C1(new_n317), .C2(new_n329), .ZN(new_n338));
  AND4_X1   g152(.A1(KEYINPUT30), .A2(new_n325), .A3(new_n298), .A4(new_n326), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT30), .B1(new_n291), .B2(new_n298), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n308), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n325), .A2(new_n298), .A3(new_n326), .A4(new_n315), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT68), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n316), .A2(new_n310), .A3(new_n325), .A4(new_n326), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n337), .B1(new_n347), .B2(new_n257), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n336), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n257), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n345), .B2(new_n346), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n351), .A2(new_n337), .B1(new_n341), .B2(new_n308), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n257), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT70), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n354), .A3(KEYINPUT31), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n335), .B1(new_n349), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G472), .A2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT32), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n331), .A2(new_n334), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n350), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n343), .A2(new_n336), .A3(new_n348), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT31), .B1(new_n352), .B2(new_n354), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT32), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n357), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n342), .A2(new_n347), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n350), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n369), .B(new_n370), .C1(new_n360), .C2(new_n350), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n325), .A2(new_n298), .A3(new_n326), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n308), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n347), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n333), .B1(new_n374), .B2(KEYINPUT28), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n350), .A2(new_n370), .ZN(new_n376));
  AOI21_X1  g190(.A(G902), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G472), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n251), .B1(new_n367), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT9), .B(G234), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT76), .ZN(new_n382));
  OAI21_X1  g196(.A(G221), .B1(new_n382), .B2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n385), .B2(G107), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G101), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT77), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n394), .A3(G101), .ZN(new_n395));
  INV_X1    g209(.A(G101), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n386), .A2(new_n389), .A3(new_n396), .A4(new_n390), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(KEYINPUT4), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n391), .B2(G101), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n295), .B(new_n393), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT10), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n385), .A2(G107), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n388), .A2(G104), .ZN(new_n403));
  OAI21_X1  g217(.A(G101), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n401), .B1(new_n324), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n296), .A2(new_n297), .ZN(new_n407));
  INV_X1    g221(.A(new_n405), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n290), .A2(KEYINPUT10), .A3(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n400), .A2(new_n406), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n296), .A2(new_n297), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n290), .A2(new_n408), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n322), .A2(new_n323), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n405), .B1(new_n414), .B2(new_n285), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n411), .B(new_n412), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT12), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT79), .B(new_n412), .C1(new_n413), .C2(new_n415), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n418), .B1(new_n416), .B2(new_n417), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n410), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  INV_X1    g238(.A(G227), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G953), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n424), .B(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n400), .A2(new_n406), .A3(new_n409), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n407), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n400), .A2(new_n406), .A3(KEYINPUT81), .A4(new_n409), .ZN(new_n431));
  INV_X1    g245(.A(new_n427), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n410), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n430), .A2(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n410), .A2(KEYINPUT80), .A3(new_n432), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n423), .A2(new_n427), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G469), .B1(new_n437), .B2(G902), .ZN(new_n438));
  XOR2_X1   g252(.A(KEYINPUT82), .B(G469), .Z(new_n439));
  INV_X1    g253(.A(new_n421), .ZN(new_n440));
  INV_X1    g254(.A(new_n422), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n433), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n430), .A2(new_n431), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n432), .B1(new_n443), .B2(new_n410), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n238), .B(new_n439), .C1(new_n442), .C2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n384), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n290), .A2(new_n206), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n295), .A2(G125), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n228), .A2(G224), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n454), .B(KEYINPUT84), .Z(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n453), .B(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT5), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G113), .B1(new_n300), .B2(KEYINPUT5), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n305), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n408), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G122), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n398), .A2(new_n399), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n308), .A2(new_n393), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n463), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT6), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  INV_X1    g283(.A(new_n464), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n470), .A2(KEYINPUT83), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(KEYINPUT6), .A3(new_n471), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n457), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT87), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT7), .B(new_n454), .C1(new_n453), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n470), .A2(KEYINPUT85), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n464), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n478), .A2(KEYINPUT8), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT8), .B1(new_n478), .B2(new_n480), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n462), .A2(new_n405), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n460), .B1(new_n458), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n459), .A2(KEYINPUT86), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n305), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n483), .B(new_n484), .C1(new_n405), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n454), .A2(new_n476), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n454), .A2(KEYINPUT7), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n451), .A2(new_n452), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n477), .A2(new_n467), .A3(new_n489), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n238), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n450), .B1(new_n475), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n493), .A2(new_n238), .ZN(new_n496));
  INV_X1    g310(.A(new_n457), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n467), .A2(KEYINPUT6), .B1(new_n469), .B2(new_n471), .ZN(new_n498));
  INV_X1    g312(.A(new_n474), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n496), .A2(new_n500), .A3(new_n449), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n448), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n200), .B(KEYINPUT19), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n199), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n507), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n268), .A3(new_n505), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n504), .A2(new_n511), .A3(new_n210), .A4(new_n213), .ZN(new_n512));
  XNOR2_X1  g326(.A(G113), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(G104), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n509), .A2(new_n505), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(KEYINPUT18), .A3(G131), .ZN(new_n516));
  NAND2_X1  g330(.A1(KEYINPUT18), .A2(G131), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(new_n505), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n200), .B(new_n199), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n512), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(G475), .A2(G902), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n508), .A2(new_n510), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n515), .A2(KEYINPUT17), .A3(G131), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n221), .A2(new_n222), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n523), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n521), .B(new_n522), .C1(new_n530), .C2(new_n514), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT20), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n221), .A2(new_n222), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n520), .B1(new_n533), .B2(new_n527), .ZN(new_n534));
  INV_X1    g348(.A(new_n514), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n521), .A4(new_n522), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n534), .B1(KEYINPUT88), .B2(new_n535), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n530), .A2(new_n541), .A3(new_n514), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n542), .A3(new_n238), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G475), .ZN(new_n544));
  NAND2_X1  g358(.A1(G234), .A2(G237), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n545), .A2(G952), .A3(new_n228), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n545), .A2(G902), .A3(G953), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT21), .B(G898), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n539), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  XOR2_X1   g365(.A(G116), .B(G122), .Z(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n388), .ZN(new_n553));
  XNOR2_X1  g367(.A(G116), .B(G122), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G107), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n281), .A2(G128), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n187), .A2(G143), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n262), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT13), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n187), .B2(G143), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n281), .A2(KEYINPUT13), .A3(G128), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n557), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G134), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT89), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n555), .A2(new_n558), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT89), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n564), .A4(new_n553), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n228), .A2(G217), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n382), .A2(new_n571), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n301), .A2(G122), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n388), .B1(new_n573), .B2(KEYINPUT14), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(new_n554), .ZN(new_n575));
  INV_X1    g389(.A(new_n558), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n262), .B1(new_n556), .B2(new_n557), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT90), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OR3_X1    g392(.A1(new_n576), .A2(KEYINPUT90), .A3(new_n577), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n570), .A2(new_n572), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n572), .B1(new_n570), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n238), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT91), .ZN(new_n584));
  INV_X1    g398(.A(G478), .ZN(new_n585));
  OR2_X1    g399(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n586));
  NAND2_X1  g400(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT91), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n589), .B(new_n238), .C1(new_n581), .C2(new_n582), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n584), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n583), .A2(new_n588), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT93), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT93), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n595), .A3(new_n592), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n551), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n446), .A2(new_n502), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n380), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  OAI21_X1  g415(.A(G472), .B1(new_n356), .B2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n364), .A2(new_n357), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n495), .A2(new_n501), .ZN(new_n604));
  AND4_X1   g418(.A1(new_n250), .A2(new_n604), .A3(new_n447), .A4(new_n550), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n602), .A2(new_n603), .A3(new_n446), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n585), .A2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n582), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n570), .A2(new_n572), .A3(new_n580), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT33), .B1(new_n610), .B2(KEYINPUT94), .ZN(new_n611));
  OAI211_X1 g425(.A(KEYINPUT94), .B(KEYINPUT33), .C1(new_n581), .C2(new_n582), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n607), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n584), .A2(new_n585), .A3(new_n590), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n539), .A2(new_n544), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n606), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n385), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n539), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n532), .A2(new_n538), .A3(KEYINPUT96), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n624), .A2(new_n625), .B1(G475), .B2(new_n543), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n594), .A3(new_n596), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n606), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G107), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NOR3_X1   g444(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT36), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n227), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n631), .A2(new_n217), .A3(new_n216), .A4(new_n226), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n249), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT97), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n247), .A2(new_n244), .A3(new_n240), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n637), .B1(new_n636), .B2(new_n638), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n602), .A2(new_n603), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n598), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT37), .B(G110), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  AOI21_X1  g460(.A(new_n365), .B1(new_n364), .B2(new_n357), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n356), .A2(KEYINPUT32), .A3(new_n358), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n379), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n641), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n639), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n546), .B1(new_n547), .B2(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n651), .A2(new_n627), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n446), .A2(new_n502), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n649), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  XOR2_X1   g472(.A(new_n653), .B(KEYINPUT39), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n446), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n662));
  INV_X1    g476(.A(new_n596), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n595), .B1(new_n591), .B2(new_n592), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n448), .B1(new_n539), .B2(new_n544), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n604), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n636), .A2(new_n638), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n661), .A2(new_n662), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n352), .A2(new_n354), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n374), .A2(new_n350), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(KEYINPUT100), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n238), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT100), .B1(new_n674), .B2(new_n675), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n367), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n673), .B1(new_n367), .B2(new_n679), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n672), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  INV_X1    g498(.A(new_n653), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n616), .A2(new_n617), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n651), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n649), .A2(new_n656), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  OAI21_X1  g503(.A(new_n238), .B1(new_n442), .B2(new_n444), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n383), .A3(new_n445), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n502), .A2(new_n550), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n618), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n649), .A2(new_n694), .A3(new_n250), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NOR3_X1   g511(.A1(new_n627), .A2(new_n692), .A3(new_n693), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n649), .A2(new_n250), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  INV_X1    g514(.A(new_n597), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n691), .A2(new_n502), .A3(new_n383), .A4(new_n445), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n701), .A2(new_n651), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n649), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  INV_X1    g519(.A(G472), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n364), .B2(new_n238), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n374), .A2(KEYINPUT28), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n334), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n350), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n362), .B2(new_n363), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n708), .B1(new_n712), .B2(new_n357), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n708), .A3(new_n357), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n691), .A2(new_n383), .A3(new_n445), .A4(new_n550), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n594), .A2(new_n604), .A3(new_n596), .A4(new_n666), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n714), .A2(new_n250), .A3(new_n715), .A4(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT103), .B(G122), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G24));
  AOI21_X1  g535(.A(new_n257), .B1(new_n709), .B2(new_n334), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n349), .B2(new_n355), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT102), .B1(new_n723), .B2(new_n358), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n602), .A2(new_n724), .A3(new_n715), .A4(new_n670), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n702), .A2(new_n686), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n206), .ZN(G27));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  AOI221_X4 g544(.A(new_n653), .B1(new_n539), .B2(new_n544), .C1(new_n614), .C2(new_n615), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n423), .A2(new_n427), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n435), .A2(new_n436), .ZN(new_n733));
  AOI21_X1  g547(.A(G902), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(G469), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n445), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n604), .A2(new_n448), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n731), .A2(new_n736), .A3(new_n383), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT42), .B1(new_n380), .B2(new_n739), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n359), .A2(new_n366), .B1(G472), .B2(new_n378), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NOR4_X1   g556(.A1(new_n741), .A2(new_n742), .A3(new_n251), .A4(new_n738), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n730), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n649), .A2(new_n250), .A3(new_n739), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n742), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n380), .A2(KEYINPUT42), .A3(new_n739), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(KEYINPUT104), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n268), .ZN(G33));
  NAND2_X1  g564(.A1(new_n736), .A2(new_n383), .ZN(new_n751));
  INV_X1    g565(.A(new_n737), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n751), .A2(new_n627), .A3(new_n752), .A4(new_n653), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n380), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  OAI21_X1  g570(.A(G469), .B1(new_n437), .B2(KEYINPUT45), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n732), .A2(new_n733), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n437), .A2(KEYINPUT105), .A3(KEYINPUT45), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n735), .A2(new_n238), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT46), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n763), .B2(new_n764), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n445), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n383), .ZN(new_n770));
  INV_X1    g584(.A(new_n659), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n756), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(KEYINPUT106), .A3(new_n383), .A4(new_n659), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n737), .B(KEYINPUT107), .ZN(new_n774));
  INV_X1    g588(.A(new_n617), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n616), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT43), .Z(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n670), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n602), .A2(new_n603), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT44), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n772), .A2(new_n773), .A3(new_n774), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NOR4_X1   g598(.A1(new_n649), .A2(new_n250), .A3(new_n686), .A4(new_n752), .ZN(new_n785));
  XNOR2_X1  g599(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n770), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n769), .B2(new_n383), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n785), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NOR2_X1   g605(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n691), .A2(new_n445), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT109), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(new_n383), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n250), .A2(new_n724), .A3(new_n602), .A4(new_n715), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n797), .A2(new_n546), .A3(new_n777), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n774), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT116), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(KEYINPUT116), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n796), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n692), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n737), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT117), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n546), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n805), .A2(KEYINPUT117), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(KEYINPUT118), .A3(new_n777), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(new_n777), .A3(new_n808), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n725), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n804), .A2(new_n669), .A3(new_n448), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n798), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n798), .A2(new_n815), .A3(new_n816), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n814), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n681), .A2(new_n251), .A3(new_n682), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n616), .A2(new_n617), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n809), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n803), .A2(new_n819), .A3(KEYINPUT51), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n810), .A2(new_n813), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT48), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT120), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n825), .A2(KEYINPUT120), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n824), .A2(new_n380), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n824), .A2(new_n380), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n829), .B2(new_n826), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n798), .A2(new_n502), .A3(new_n804), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT119), .ZN(new_n832));
  INV_X1    g646(.A(new_n618), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n809), .A2(new_n833), .A3(new_n820), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n832), .A2(G952), .A3(new_n228), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  INV_X1    g651(.A(new_n814), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n818), .A2(new_n817), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n822), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n840), .B2(new_n802), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n823), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n642), .A2(new_n665), .A3(new_n626), .A4(new_n685), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n741), .A2(new_n844), .A3(new_n655), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT114), .B1(new_n845), .B2(new_n728), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n717), .A2(new_n670), .A3(new_n653), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n446), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n681), .B2(new_n682), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n602), .A2(new_n724), .A3(new_n715), .A4(new_n670), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n726), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n657), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n846), .A2(new_n850), .A3(new_n854), .A4(new_n688), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n856));
  OR3_X1    g670(.A1(new_n725), .A2(KEYINPUT113), .A3(new_n738), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT113), .B1(new_n725), .B2(new_n738), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n642), .A2(new_n446), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n593), .A2(new_n653), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n737), .A2(new_n626), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n737), .A2(KEYINPUT112), .A3(new_n626), .A4(new_n861), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n380), .A2(new_n753), .B1(new_n866), .B2(new_n649), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n606), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n380), .A2(new_n599), .B1(new_n869), .B2(new_n833), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n775), .A2(new_n593), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n606), .A2(new_n871), .B1(new_n643), .B2(new_n598), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT111), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n874));
  OAI221_X1 g688(.A(new_n874), .B1(new_n643), .B2(new_n598), .C1(new_n606), .C2(new_n871), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n868), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n655), .B1(new_n367), .B2(new_n379), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n878), .A2(new_n654), .B1(new_n851), .B2(new_n726), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT52), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n850), .A2(new_n879), .A3(new_n880), .A4(new_n688), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT53), .B1(new_n740), .B2(new_n743), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n695), .A2(new_n699), .A3(new_n719), .A4(new_n704), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n856), .A2(new_n877), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n380), .A2(new_n698), .B1(new_n797), .B2(new_n718), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(KEYINPUT110), .A3(new_n695), .A4(new_n704), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT110), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n852), .A2(new_n657), .A3(new_n688), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n679), .B1(new_n647), .B2(new_n648), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT101), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n848), .B1(new_n894), .B2(new_n680), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT52), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n881), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n744), .A2(new_n748), .A3(new_n859), .A4(new_n867), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n891), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n843), .B(new_n885), .C1(new_n899), .C2(KEYINPUT53), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT115), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n891), .A2(new_n898), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n881), .A4(new_n856), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(KEYINPUT54), .C1(new_n904), .C2(new_n899), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n886), .A2(new_n888), .A3(new_n890), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n896), .A2(new_n881), .ZN(new_n908));
  AND4_X1   g722(.A1(new_n744), .A2(new_n748), .A3(new_n859), .A4(new_n867), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n904), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(KEYINPUT115), .A3(new_n843), .A4(new_n885), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n902), .A2(new_n906), .A3(new_n912), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n842), .A2(new_n913), .B1(G952), .B2(G953), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n794), .A2(KEYINPUT49), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n794), .A2(KEYINPUT49), .ZN(new_n916));
  INV_X1    g730(.A(new_n776), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n383), .A2(new_n669), .A3(new_n447), .A4(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n820), .A2(new_n915), .A3(new_n916), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n914), .A2(new_n919), .ZN(G75));
  NAND2_X1  g734(.A1(new_n911), .A2(new_n885), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(G210), .A3(G902), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n498), .A2(new_n499), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n497), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT55), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n922), .B2(new_n923), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n228), .A2(G952), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G51));
  XNOR2_X1  g744(.A(new_n764), .B(KEYINPUT57), .ZN(new_n931));
  INV_X1    g745(.A(new_n900), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n843), .B1(new_n911), .B2(new_n885), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n444), .B2(new_n442), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n921), .A2(G902), .A3(new_n763), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(G54));
  NAND2_X1  g751(.A1(new_n536), .A2(new_n521), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n921), .A2(G902), .ZN(new_n939));
  NAND2_X1  g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n929), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n939), .A2(new_n938), .A3(new_n940), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(G60));
  NOR2_X1   g759(.A1(new_n611), .A2(new_n613), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT121), .Z(new_n947));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT59), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n913), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n949), .B(new_n947), .C1(new_n932), .C2(new_n933), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n942), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n950), .A2(new_n952), .ZN(G63));
  XNOR2_X1  g767(.A(new_n241), .B(KEYINPUT60), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n911), .B2(new_n885), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n633), .A2(new_n634), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n929), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n248), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT53), .B1(new_n903), .B2(new_n908), .ZN(new_n959));
  INV_X1    g773(.A(new_n885), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n958), .B1(new_n961), .B2(new_n954), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n957), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n954), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n956), .B(new_n966), .C1(new_n959), .C2(new_n960), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n967), .B(new_n942), .C1(new_n955), .C2(new_n248), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n963), .A3(new_n942), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(KEYINPUT61), .A3(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n965), .A2(new_n970), .ZN(G66));
  INV_X1    g785(.A(new_n548), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n228), .B1(new_n972), .B2(G224), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n891), .B2(new_n228), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n924), .B1(G898), .B2(new_n228), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n974), .B(new_n975), .Z(G69));
  AOI211_X1 g790(.A(new_n752), .B(new_n660), .C1(new_n618), .C2(new_n871), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n380), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n783), .A2(new_n790), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n852), .A2(new_n657), .ZN(new_n981));
  AOI22_X1  g795(.A1(new_n981), .A2(KEYINPUT114), .B1(new_n878), .B2(new_n687), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(new_n683), .A3(new_n854), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n982), .A2(KEYINPUT62), .A3(new_n683), .A4(new_n854), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(G953), .B1(new_n980), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n341), .B(new_n503), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT123), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n989), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(G900), .B2(G953), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n982), .A2(new_n854), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n749), .B(new_n993), .C1(new_n380), .C2(new_n753), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n741), .A2(new_n251), .A3(new_n717), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n772), .A2(new_n773), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT124), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n783), .A2(new_n790), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n994), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n992), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT123), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n979), .B1(new_n985), .B2(new_n986), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n1001), .B(new_n991), .C1(new_n1002), .C2(G953), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n990), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n425), .B2(new_n652), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT125), .Z(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n990), .A2(new_n1000), .A3(new_n1003), .A4(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(new_n368), .A2(new_n257), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n980), .A2(new_n907), .A3(new_n987), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT63), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT126), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1011), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1014), .B1(new_n674), .B2(new_n369), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n905), .B(new_n1017), .C1(new_n904), .C2(new_n899), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n942), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1015), .B1(new_n999), .B2(new_n891), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n368), .A2(new_n257), .ZN(new_n1021));
  AOI211_X1 g835(.A(new_n1016), .B(new_n1019), .C1(new_n1020), .C2(new_n1021), .ZN(G57));
endmodule


