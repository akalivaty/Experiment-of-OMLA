//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT85), .ZN(new_n210));
  INV_X1    g009(.A(G1gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(KEYINPUT85), .A3(G1gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n216), .A2(G8gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(G8gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT14), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT14), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT84), .B(G36gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n226), .B(KEYINPUT15), .C1(new_n220), .C2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT15), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n227), .A2(new_n220), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(new_n225), .ZN(new_n231));
  XNOR2_X1  g030(.A(G43gat), .B(G50gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n230), .A2(new_n225), .ZN(new_n235));
  INV_X1    g034(.A(new_n232), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(KEYINPUT15), .A3(new_n236), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n234), .B1(new_n233), .B2(new_n237), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n219), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT86), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT87), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n217), .B2(new_n218), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n216), .A2(G8gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n216), .A2(G8gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(KEYINPUT87), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n237), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n219), .B(KEYINPUT86), .C1(new_n238), .C2(new_n239), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n242), .A2(new_n243), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n243), .B(KEYINPUT13), .Z(new_n256));
  INV_X1    g055(.A(new_n250), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n249), .B1(new_n245), .B2(new_n248), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n252), .B2(new_n253), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n208), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n252), .A2(KEYINPUT88), .A3(new_n253), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n259), .B(new_n207), .C1(new_n252), .C2(new_n253), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n261), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G15gat), .B(G43gat), .Z(new_n269));
  XNOR2_X1  g068(.A(G71gat), .B(G99gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G227gat), .ZN(new_n272));
  INV_X1    g071(.A(G233gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT25), .ZN(new_n276));
  NAND3_X1  g075(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT66), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(G183gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n276), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT23), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n291), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n285), .A2(new_n281), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(new_n277), .C1(new_n279), .C2(KEYINPUT64), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n279), .A2(KEYINPUT64), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n293), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n295), .B1(new_n301), .B2(KEYINPUT25), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT27), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT67), .B1(new_n304), .B2(G183gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(new_n282), .A3(new_n284), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n285), .A2(KEYINPUT27), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(G183gat), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT67), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n303), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n282), .A2(new_n284), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n311), .A2(KEYINPUT28), .A3(new_n307), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(G169gat), .ZN(new_n315));
  INV_X1    g114(.A(G176gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT26), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n290), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n314), .B(new_n317), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n313), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G134gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G127gat), .ZN(new_n325));
  INV_X1    g124(.A(G127gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G134gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(KEYINPUT1), .ZN(new_n330));
  INV_X1    g129(.A(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G113gat), .ZN(new_n332));
  INV_X1    g131(.A(G113gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G120gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G127gat), .B(G134gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n302), .A2(new_n323), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n330), .A2(new_n338), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n320), .B1(KEYINPUT23), .B2(new_n288), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n342), .B(new_n292), .C1(new_n297), .C2(new_n299), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n343), .A2(new_n276), .B1(new_n287), .B2(new_n294), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n321), .B1(new_n310), .B2(new_n312), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n275), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n271), .B1(new_n347), .B2(KEYINPUT33), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT32), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n340), .A2(new_n346), .ZN(new_n352));
  AOI221_X4 g151(.A(new_n349), .B1(KEYINPUT33), .B2(new_n271), .C1(new_n352), .C2(new_n274), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n352), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n274), .A2(KEYINPUT34), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT70), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n274), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n340), .A2(new_n346), .A3(KEYINPUT69), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n362), .B2(KEYINPUT34), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT34), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT70), .B(new_n364), .C1(new_n360), .C2(new_n361), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n354), .B(new_n357), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n357), .B1(new_n363), .B2(new_n365), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT68), .B1(new_n351), .B2(new_n353), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n274), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n372), .A3(new_n271), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT68), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n350), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n367), .A2(new_n368), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G228gat), .A2(G233gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT2), .ZN(new_n380));
  OR2_X1    g179(.A1(G141gat), .A2(G148gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n384), .A3(new_n382), .ZN(new_n385));
  XNOR2_X1  g184(.A(G155gat), .B(G162gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(G141gat), .A2(G148gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n380), .B(new_n390), .C1(new_n393), .C2(new_n384), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G211gat), .B(G218gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(G197gat), .A2(G204gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n406));
  OAI21_X1  g205(.A(G218gat), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT22), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n401), .B1(new_n409), .B2(KEYINPUT73), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT73), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT72), .B(G211gat), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT22), .B1(new_n412), .B2(G218gat), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n411), .B(new_n400), .C1(new_n413), .C2(new_n404), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n378), .B1(new_n399), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(new_n414), .A3(new_n398), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n395), .B1(new_n417), .B2(new_n396), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(KEYINPUT79), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n420));
  AOI211_X1 g219(.A(new_n420), .B(new_n395), .C1(new_n417), .C2(new_n396), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT80), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(new_n396), .ZN(new_n423));
  INV_X1    g222(.A(new_n395), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n420), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n418), .A2(KEYINPUT79), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .A4(new_n416), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n422), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  INV_X1    g230(.A(G218gat), .ZN(new_n432));
  OR2_X1    g231(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n435), .A2(KEYINPUT22), .B1(new_n403), .B2(new_n402), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT29), .B1(new_n436), .B2(new_n400), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n409), .A2(new_n401), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(KEYINPUT78), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n396), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT78), .B1(new_n437), .B2(new_n438), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n424), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n400), .B1(new_n436), .B2(new_n411), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n409), .A2(KEYINPUT73), .A3(new_n401), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT3), .B1(new_n387), .B2(new_n394), .ZN(new_n445));
  OAI22_X1  g244(.A1(new_n443), .A2(new_n444), .B1(new_n445), .B2(KEYINPUT29), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n378), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n430), .A2(new_n431), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n431), .B1(new_n430), .B2(new_n448), .ZN(new_n450));
  XNOR2_X1  g249(.A(G78gat), .B(G106gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT31), .B(G50gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n449), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n378), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n446), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n425), .B2(new_n420), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n427), .B1(new_n458), .B2(new_n428), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n419), .A2(KEYINPUT80), .A3(new_n421), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n448), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G22gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n430), .A2(new_n431), .A3(new_n448), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n453), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n366), .B(new_n377), .C1(new_n455), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n387), .A2(new_n394), .A3(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n397), .A2(new_n341), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n339), .A2(new_n395), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT4), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n339), .A2(new_n395), .A3(KEYINPUT4), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n467), .A2(new_n470), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n341), .A2(new_n394), .A3(new_n387), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n471), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT77), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n470), .A2(new_n472), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n482), .A2(new_n474), .A3(new_n471), .A4(new_n467), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT77), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n473), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G1gat), .B(G29gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT0), .ZN(new_n488));
  XNOR2_X1  g287(.A(G57gat), .B(G85gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT6), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n490), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n480), .A2(new_n492), .A3(new_n483), .A4(new_n485), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n483), .A2(new_n485), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n484), .B1(new_n473), .B2(new_n478), .ZN(new_n496));
  OAI211_X1 g295(.A(KEYINPUT6), .B(new_n490), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT75), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n500));
  NAND2_X1  g299(.A1(G226gat), .A2(G233gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n344), .B2(new_n345), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(new_n302), .B2(new_n323), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(new_n502), .ZN(new_n505));
  INV_X1    g304(.A(new_n415), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n398), .B1(new_n344), .B2(new_n345), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT74), .B1(new_n508), .B2(new_n501), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n501), .B1(new_n302), .B2(new_n323), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n501), .B2(new_n508), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT74), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n507), .B1(new_n514), .B2(new_n506), .ZN(new_n515));
  XNOR2_X1  g314(.A(G8gat), .B(G36gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(G64gat), .B(G92gat), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n516), .B(new_n517), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n499), .B(new_n500), .C1(new_n515), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n512), .A2(new_n415), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n509), .B1(new_n505), .B2(KEYINPUT74), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n521), .B(new_n519), .C1(new_n522), .C2(new_n415), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n501), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n513), .B1(new_n524), .B2(new_n503), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n506), .B1(new_n525), .B2(new_n509), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n519), .B1(new_n526), .B2(new_n521), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT30), .B1(new_n527), .B2(KEYINPUT75), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n498), .A2(new_n520), .A3(new_n523), .A4(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT35), .B1(new_n465), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n520), .A3(new_n523), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT82), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n486), .A2(new_n533), .A3(KEYINPUT6), .A4(new_n490), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n532), .A2(new_n534), .B1(new_n491), .B2(new_n493), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n531), .A2(new_n535), .A3(KEYINPUT35), .ZN(new_n536));
  INV_X1    g335(.A(new_n366), .ZN(new_n537));
  INV_X1    g336(.A(new_n361), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT69), .B1(new_n340), .B2(new_n346), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n538), .A2(new_n539), .A3(new_n274), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT70), .B1(new_n540), .B2(new_n364), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n362), .A2(new_n358), .A3(KEYINPUT34), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n354), .B1(new_n543), .B2(new_n357), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n454), .B1(new_n449), .B2(new_n450), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n462), .A2(new_n463), .A3(new_n453), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n536), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT36), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n537), .B2(new_n544), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n541), .A2(new_n542), .B1(new_n355), .B2(new_n356), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n368), .A2(new_n376), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n366), .B(KEYINPUT36), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n515), .A2(KEYINPUT37), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n519), .A2(KEYINPUT37), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n523), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT38), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n522), .A2(new_n415), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n564), .B1(new_n505), .B2(new_n506), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT38), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n527), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(new_n535), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n486), .A2(new_n490), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT40), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT39), .B1(new_n476), .B2(new_n477), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n482), .A2(new_n467), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(new_n477), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT39), .ZN(new_n574));
  INV_X1    g373(.A(new_n467), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n574), .B(new_n477), .C1(new_n481), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n492), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n570), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n573), .ZN(new_n580));
  INV_X1    g379(.A(new_n577), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(KEYINPUT40), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT81), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT81), .A4(KEYINPUT40), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n579), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n531), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n587), .A3(new_n548), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n377), .A2(KEYINPUT71), .A3(KEYINPUT36), .A4(new_n366), .ZN(new_n589));
  INV_X1    g388(.A(new_n498), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n547), .B(new_n546), .C1(new_n590), .C2(new_n531), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n557), .A2(new_n588), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n268), .B1(new_n550), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT9), .ZN(new_n596));
  OR2_X1    g395(.A1(G57gat), .A2(G64gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(G57gat), .A2(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n600), .B2(new_n599), .ZN(new_n602));
  OR2_X1    g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n603), .B2(new_n596), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n597), .A2(KEYINPUT91), .A3(new_n598), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT91), .B1(new_n597), .B2(new_n598), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n608), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT92), .B1(new_n615), .B2(new_n607), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n606), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(new_n326), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n611), .A2(new_n612), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n615), .A2(KEYINPUT92), .A3(new_n607), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n623), .A2(new_n624), .B1(new_n602), .B2(new_n605), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n245), .A2(new_n248), .B1(KEYINPUT21), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n622), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT94), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n630));
  INV_X1    g429(.A(G155gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n627), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n642));
  INV_X1    g441(.A(new_n249), .ZN(new_n643));
  XOR2_X1   g442(.A(G99gat), .B(G106gat), .Z(new_n644));
  NAND2_X1  g443(.A1(G99gat), .A2(G106gat), .ZN(new_n645));
  INV_X1    g444(.A(G85gat), .ZN(new_n646));
  INV_X1    g445(.A(G92gat), .ZN(new_n647));
  AOI22_X1  g446(.A1(KEYINPUT8), .A2(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(G85gat), .A3(G92gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT7), .Z(new_n653));
  OAI21_X1  g452(.A(new_n644), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n648), .B(KEYINPUT98), .ZN(new_n655));
  INV_X1    g454(.A(new_n644), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n652), .B(KEYINPUT7), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n642), .B1(new_n643), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n659), .B1(new_n238), .B2(new_n239), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n654), .A2(new_n658), .ZN(new_n665));
  INV_X1    g464(.A(new_n239), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT99), .B1(new_n668), .B2(new_n660), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT95), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT96), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n664), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n664), .B2(new_n669), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n639), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n664), .A2(new_n669), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n672), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n638), .A3(new_n674), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n606), .B(KEYINPUT10), .C1(new_n613), .C2(new_n616), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n683), .B2(new_n659), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n665), .A2(KEYINPUT101), .A3(KEYINPUT10), .A4(new_n625), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n644), .A2(KEYINPUT100), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n665), .A2(new_n625), .A3(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n606), .B(new_n687), .C1(new_n613), .C2(new_n616), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n659), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT10), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(G230gat), .A2(G233gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n688), .B2(new_n690), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(G120gat), .B(G148gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n696), .B2(new_n697), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n695), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n694), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n705), .B1(new_n686), .B2(new_n692), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n702), .B1(new_n706), .B2(new_n696), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n635), .A2(new_n681), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n595), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n590), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g512(.A1(new_n711), .A2(KEYINPUT104), .A3(new_n531), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  INV_X1    g514(.A(new_n531), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n710), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(G8gat), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT16), .B(G8gat), .Z(new_n719));
  NAND4_X1  g518(.A1(new_n711), .A2(KEYINPUT42), .A3(new_n531), .A4(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n719), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n714), .B2(new_n717), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n723));
  OAI211_X1 g522(.A(new_n718), .B(new_n720), .C1(new_n722), .C2(new_n723), .ZN(G1325gat));
  INV_X1    g523(.A(G15gat), .ZN(new_n725));
  INV_X1    g524(.A(new_n545), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n710), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n556), .A2(new_n553), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n367), .B1(new_n351), .B2(new_n353), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT36), .B1(new_n729), .B2(new_n366), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n589), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n557), .A2(KEYINPUT105), .A3(new_n589), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G15gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT106), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n727), .B1(new_n710), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT107), .Z(G1326gat));
  INV_X1    g538(.A(new_n548), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n711), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT43), .B(G22gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1327gat));
  INV_X1    g542(.A(new_n708), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n635), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n681), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n595), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n220), .A3(new_n590), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n677), .A2(new_n680), .A3(KEYINPUT108), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT108), .B1(new_n677), .B2(new_n680), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n588), .A2(new_n591), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n733), .A2(new_n758), .A3(new_n734), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n759), .B2(new_n550), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n550), .A2(new_n592), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n756), .B1(new_n761), .B2(new_n681), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n268), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G29gat), .B1(new_n765), .B2(new_n498), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n766), .A3(new_n767), .ZN(G1328gat));
  INV_X1    g567(.A(new_n227), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n765), .B2(new_n716), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n749), .A2(new_n531), .A3(new_n227), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n771), .A2(KEYINPUT109), .A3(KEYINPUT46), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT109), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n773));
  OAI221_X1 g572(.A(new_n770), .B1(KEYINPUT46), .B2(new_n771), .C1(new_n772), .C2(new_n773), .ZN(G1329gat));
  INV_X1    g573(.A(new_n765), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n735), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G43gat), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n726), .A2(G43gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n748), .B2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n780), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n777), .B(new_n782), .C1(new_n748), .C2(new_n778), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1330gat));
  INV_X1    g583(.A(G50gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n748), .B2(new_n548), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n740), .A2(G50gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n765), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g588(.A1(new_n759), .A2(new_n550), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n634), .A2(new_n268), .A3(new_n746), .A4(new_n708), .ZN(new_n792));
  OR3_X1    g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n790), .B2(new_n792), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n590), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n531), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT49), .B(G64gat), .Z(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n798), .B2(new_n800), .ZN(G1333gat));
  NAND2_X1  g600(.A1(new_n795), .A2(new_n735), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G71gat), .ZN(new_n803));
  INV_X1    g602(.A(G71gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n795), .A2(new_n804), .A3(new_n545), .ZN(new_n805));
  XNOR2_X1  g604(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n803), .B2(new_n805), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(G1334gat));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n740), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g611(.A1(new_n635), .A2(new_n268), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n744), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n760), .B2(new_n762), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT113), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n817), .B(new_n814), .C1(new_n760), .C2(new_n762), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n590), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT114), .B1(new_n790), .B2(new_n746), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n746), .B1(new_n759), .B2(new_n550), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n813), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n821), .A2(new_n824), .A3(KEYINPUT51), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT51), .B1(new_n821), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n590), .A2(new_n646), .A3(new_n708), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n820), .A2(new_n646), .B1(new_n827), .B2(new_n828), .ZN(G1336gat));
  NOR3_X1   g628(.A1(new_n716), .A2(G92gat), .A3(new_n744), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n825), .B2(new_n826), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832));
  OAI21_X1  g631(.A(G92gat), .B1(new_n815), .B2(new_n716), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n531), .A3(new_n818), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G92gat), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT115), .B1(new_n837), .B2(KEYINPUT52), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n839), .B(new_n832), .C1(new_n831), .C2(new_n836), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n834), .B1(new_n838), .B2(new_n840), .ZN(G1337gat));
  AND2_X1   g640(.A1(new_n819), .A2(new_n735), .ZN(new_n842));
  INV_X1    g641(.A(G99gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n545), .A2(new_n843), .A3(new_n708), .ZN(new_n844));
  OAI22_X1  g643(.A1(new_n842), .A2(new_n843), .B1(new_n827), .B2(new_n844), .ZN(G1338gat));
  OR2_X1    g644(.A1(new_n825), .A2(new_n826), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n548), .A2(G106gat), .A3(new_n744), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(KEYINPUT117), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n763), .A2(new_n740), .A3(new_n814), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT116), .B(G106gat), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT117), .B1(new_n846), .B2(new_n847), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n816), .A2(new_n740), .A3(new_n818), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n846), .A2(new_n847), .B1(new_n855), .B2(new_n850), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n852), .A2(new_n853), .B1(new_n854), .B2(new_n856), .ZN(G1339gat));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n252), .A2(KEYINPUT88), .A3(new_n253), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT88), .B1(new_n252), .B2(new_n253), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n859), .A2(new_n266), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n242), .A2(new_n250), .A3(new_n251), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(G229gat), .A3(G233gat), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n257), .A2(new_n258), .A3(new_n256), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n206), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n708), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n686), .A2(new_n692), .A3(new_n705), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n695), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n701), .B1(new_n706), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(KEYINPUT55), .A3(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n704), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n686), .A2(new_n692), .A3(new_n705), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n706), .A3(new_n870), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n693), .A2(new_n870), .A3(new_n694), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n702), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n874), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n873), .A2(new_n267), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n755), .B1(new_n867), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n753), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n879), .A2(new_n704), .A3(new_n872), .ZN(new_n883));
  INV_X1    g682(.A(new_n754), .ZN(new_n884));
  AND4_X1   g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .A4(new_n866), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n858), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n755), .A2(new_n866), .A3(new_n883), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n861), .A2(new_n744), .A3(new_n865), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n267), .B2(new_n883), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n887), .B(KEYINPUT118), .C1(new_n889), .C2(new_n755), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n886), .A2(new_n890), .A3(new_n635), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n709), .A2(new_n268), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n726), .A2(new_n740), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n590), .A3(new_n716), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n896), .A2(new_n333), .A3(new_n268), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n498), .B1(new_n891), .B2(new_n892), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n465), .A2(new_n531), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(G113gat), .B1(new_n901), .B2(new_n267), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n897), .A2(new_n902), .ZN(G1340gat));
  OAI21_X1  g702(.A(G120gat), .B1(new_n896), .B2(new_n744), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n708), .A2(new_n331), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT119), .Z(new_n906));
  OAI21_X1  g705(.A(new_n904), .B1(new_n900), .B2(new_n906), .ZN(G1341gat));
  OAI21_X1  g706(.A(G127gat), .B1(new_n896), .B2(new_n635), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n901), .A2(new_n326), .A3(new_n634), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1342gat));
  OAI21_X1  g709(.A(G134gat), .B1(new_n896), .B2(new_n746), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n901), .A2(new_n324), .A3(new_n681), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT56), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n912), .B2(KEYINPUT56), .ZN(new_n915));
  OAI221_X1 g714(.A(new_n911), .B1(KEYINPUT56), .B2(new_n912), .C1(new_n914), .C2(new_n915), .ZN(G1343gat));
  NOR3_X1   g715(.A1(new_n735), .A2(new_n498), .A3(new_n531), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT57), .B1(new_n893), .B2(new_n740), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n740), .A2(KEYINPUT57), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n869), .A2(new_n871), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT121), .B1(new_n920), .B2(new_n874), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  AOI211_X1 g721(.A(new_n922), .B(KEYINPUT55), .C1(new_n869), .C2(new_n871), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n873), .B(new_n267), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n681), .B1(new_n924), .B2(new_n867), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n635), .B1(new_n925), .B2(new_n885), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n919), .B1(new_n892), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n917), .B1(new_n918), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G141gat), .B1(new_n928), .B2(new_n268), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n735), .A2(new_n531), .A3(new_n548), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n898), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(G141gat), .A3(new_n268), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(KEYINPUT58), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g735(.A(KEYINPUT122), .B(new_n917), .C1(new_n918), .C2(new_n927), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n267), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n932), .B1(new_n938), .B2(G141gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(G1344gat));
  AND2_X1   g740(.A1(new_n891), .A2(new_n892), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n883), .A2(new_n866), .A3(new_n681), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n943), .B1(new_n925), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n872), .A2(new_n704), .ZN(new_n947));
  INV_X1    g746(.A(new_n266), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n263), .A3(new_n264), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n261), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n879), .A2(new_n922), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n920), .A2(KEYINPUT121), .A3(new_n874), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n888), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g753(.A(KEYINPUT123), .B(new_n944), .C1(new_n954), .C2(new_n681), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n946), .A2(new_n955), .A3(new_n635), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n548), .B1(new_n956), .B2(new_n892), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n942), .A2(new_n919), .B1(new_n957), .B2(KEYINPUT57), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(new_n708), .A3(new_n917), .ZN(new_n959));
  INV_X1    g758(.A(G148gat), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT59), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n936), .A2(new_n708), .A3(new_n937), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n960), .A2(KEYINPUT59), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n931), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n960), .A3(new_n708), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1345gat));
  NAND3_X1  g766(.A1(new_n965), .A2(new_n631), .A3(new_n634), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n936), .A2(new_n634), .A3(new_n937), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(new_n631), .ZN(G1346gat));
  AOI21_X1  g769(.A(G162gat), .B1(new_n965), .B2(new_n681), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n936), .A2(new_n937), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n755), .A2(G162gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G1347gat));
  AOI21_X1  g773(.A(new_n590), .B1(new_n891), .B2(new_n892), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n465), .A2(new_n716), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(G169gat), .B1(new_n978), .B2(new_n267), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n716), .A2(new_n590), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n893), .A2(new_n894), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n268), .A2(new_n315), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1348gat));
  AOI21_X1  g782(.A(new_n316), .B1(new_n981), .B2(new_n708), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n977), .A2(G176gat), .A3(new_n744), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(new_n985), .ZN(G1349gat));
  AOI21_X1  g785(.A(new_n285), .B1(new_n981), .B2(new_n634), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n307), .A2(new_n308), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n977), .A2(new_n988), .A3(new_n635), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g789(.A(new_n990), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g790(.A1(new_n978), .A2(new_n311), .A3(new_n755), .ZN(new_n992));
  INV_X1    g791(.A(new_n981), .ZN(new_n993));
  OAI21_X1  g792(.A(G190gat), .B1(new_n993), .B2(new_n746), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G1351gat));
  NOR3_X1   g796(.A1(new_n735), .A2(new_n716), .A3(new_n548), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n975), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n999), .A2(G197gat), .A3(new_n268), .ZN(new_n1000));
  XOR2_X1   g799(.A(new_n1000), .B(KEYINPUT124), .Z(new_n1001));
  NOR3_X1   g800(.A1(new_n735), .A2(new_n590), .A3(new_n716), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n958), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(new_n267), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(G197gat), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1001), .A2(new_n1005), .ZN(G1352gat));
  NAND2_X1  g805(.A1(new_n956), .A2(new_n892), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT57), .B1(new_n1007), .B2(new_n740), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n919), .B1(new_n891), .B2(new_n892), .ZN(new_n1009));
  OAI211_X1 g808(.A(new_n708), .B(new_n1002), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g811(.A1(new_n958), .A2(KEYINPUT125), .A3(new_n708), .A4(new_n1002), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1012), .A2(G204gat), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n744), .A2(G204gat), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n975), .A2(new_n998), .A3(new_n1015), .ZN(new_n1016));
  XOR2_X1   g815(.A(new_n1016), .B(KEYINPUT62), .Z(new_n1017));
  NAND2_X1  g816(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(KEYINPUT126), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1014), .A2(new_n1020), .A3(new_n1017), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1019), .A2(new_n1021), .ZN(G1353gat));
  OR3_X1    g821(.A1(new_n999), .A2(new_n412), .A3(new_n635), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1003), .A2(new_n634), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n1024), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1025));
  AOI21_X1  g824(.A(KEYINPUT63), .B1(new_n1024), .B2(G211gat), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(G1354gat));
  INV_X1    g826(.A(new_n755), .ZN(new_n1028));
  OAI21_X1  g827(.A(new_n432), .B1(new_n999), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g828(.A1(new_n1029), .A2(KEYINPUT127), .ZN(new_n1030));
  AND2_X1   g829(.A1(new_n1029), .A2(KEYINPUT127), .ZN(new_n1031));
  NOR2_X1   g830(.A1(new_n746), .A2(new_n432), .ZN(new_n1032));
  AOI211_X1 g831(.A(new_n1030), .B(new_n1031), .C1(new_n1003), .C2(new_n1032), .ZN(G1355gat));
endmodule


