//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(KEYINPUT3), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(G137), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n460), .A2(new_n461), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(new_n463), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT67), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n471), .A3(new_n468), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(KEYINPUT65), .A3(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n473), .A2(new_n483), .ZN(G160));
  AND3_X1   g059(.A1(new_n462), .A2(G2105), .A3(new_n465), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n463), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n462), .A2(new_n465), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n463), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n489), .B1(G136), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT68), .ZN(G162));
  NAND2_X1  g069(.A1(new_n485), .A2(G126), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n463), .A2(G138), .ZN(new_n499));
  OR2_X1    g074(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n479), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n462), .A2(new_n465), .A3(new_n499), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n503), .B1(new_n505), .B2(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n498), .B1(new_n506), .B2(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT72), .A3(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(new_n514), .B1(KEYINPUT5), .B2(new_n511), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT71), .A3(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n518), .A2(new_n520), .B1(KEYINPUT6), .B2(new_n517), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n517), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n526), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  INV_X1    g105(.A(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  INV_X1    g107(.A(new_n524), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n515), .A2(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n532), .A2(new_n534), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  AOI22_X1  g116(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(G651), .A3(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(G90), .A2(new_n531), .B1(new_n533), .B2(G52), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n522), .A2(new_n550), .B1(new_n524), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n512), .A2(new_n514), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g141(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n567));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  NAND2_X1  g145(.A1(new_n531), .A2(G91), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n533), .A2(G53), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT78), .Z(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n558), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n573), .A2(new_n575), .A3(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n531), .A2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n533), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n522), .A2(new_n586), .B1(new_n524), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n517), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n589), .A2(new_n592), .ZN(G305));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n522), .A2(new_n594), .B1(new_n524), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n517), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n596), .A2(new_n598), .ZN(G290));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(G301), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n558), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n533), .B2(G54), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n606));
  NAND3_X1  g181(.A1(new_n531), .A2(G92), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n606), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n522), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n605), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT80), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n601), .B1(new_n613), .B2(new_n600), .ZN(G284));
  AOI21_X1  g189(.A(new_n601), .B1(new_n613), .B2(new_n600), .ZN(G321));
  NAND2_X1  g190(.A1(G299), .A2(new_n600), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n600), .B2(G168), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(new_n600), .B2(G168), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(new_n619), .B2(G860), .ZN(G148));
  NOR2_X1   g195(.A1(new_n564), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n619), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n485), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n463), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(G135), .ZN(new_n629));
  OAI221_X1 g204(.A(new_n626), .B1(new_n627), .B2(new_n628), .C1(new_n491), .C2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT82), .Z(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT83), .B(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n467), .A2(new_n463), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(new_n479), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n651), .B(new_n652), .Z(new_n653));
  OR2_X1    g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n662), .B2(new_n658), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n673), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n673), .B2(new_n679), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  MUX2_X1   g266(.A(G24), .B(G290), .S(G16), .Z(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT87), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G25), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n492), .A2(G131), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n485), .A2(G119), .ZN(new_n698));
  OR2_X1    g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n696), .B1(new_n702), .B2(new_n695), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  XOR2_X1   g279(.A(new_n703), .B(new_n704), .Z(new_n705));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n706));
  AOI211_X1 g281(.A(new_n694), .B(new_n705), .C1(new_n706), .C2(KEYINPUT36), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n708), .A2(G22), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G166), .B2(new_n708), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1971), .ZN(new_n716));
  MUX2_X1   g291(.A(G6), .B(G305), .S(G16), .Z(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT89), .Z(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT32), .B(G1981), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n713), .B(new_n716), .C1(new_n718), .C2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n720), .B2(new_n718), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n707), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n723), .B2(new_n722), .ZN(new_n725));
  OR3_X1    g300(.A1(new_n725), .A2(new_n706), .A3(KEYINPUT36), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n706), .B2(KEYINPUT36), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n613), .A2(new_n708), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G4), .B2(new_n708), .ZN(new_n729));
  INV_X1    g304(.A(G1348), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G19), .ZN(new_n732));
  OR3_X1    g307(.A1(new_n732), .A2(KEYINPUT91), .A3(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(KEYINPUT91), .B1(new_n732), .B2(G16), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n733), .B(new_n734), .C1(new_n564), .C2(new_n708), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n708), .A2(G20), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT23), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G299), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1956), .ZN(new_n740));
  INV_X1    g315(.A(G34), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(KEYINPUT24), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(KEYINPUT24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n695), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G160), .B2(new_n695), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(G2084), .Z(new_n746));
  NAND4_X1  g321(.A1(new_n731), .A2(new_n736), .A3(new_n740), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n695), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n695), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(G2078), .ZN(new_n750));
  NAND2_X1  g325(.A1(G171), .A2(G16), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G5), .B2(G16), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G35), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G162), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT29), .B(G2090), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n750), .B1(new_n752), .B2(new_n753), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G21), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G168), .B2(G16), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT94), .B(G1966), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT30), .B(G28), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n762), .B1(new_n695), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n631), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n761), .B(new_n764), .C1(new_n695), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G2078), .B2(new_n749), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n729), .A2(new_n730), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n755), .A2(new_n756), .B1(new_n752), .B2(new_n753), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n695), .A2(G32), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n492), .A2(G141), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n485), .A2(G129), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT26), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n635), .A2(G105), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n771), .A2(new_n772), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n770), .B1(new_n779), .B2(new_n695), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT27), .B(G1996), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n492), .A2(G139), .ZN(new_n783));
  NAND2_X1  g358(.A1(G115), .A2(G2104), .ZN(new_n784));
  INV_X1    g359(.A(G127), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n476), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n463), .B1(new_n786), .B2(KEYINPUT93), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(KEYINPUT93), .B2(new_n786), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT25), .Z(new_n790));
  NAND3_X1  g365(.A1(new_n783), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G33), .B(new_n791), .S(G29), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2072), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n695), .A2(G26), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT28), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n492), .A2(G140), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n485), .A2(G128), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT92), .B1(G104), .B2(G2105), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(KEYINPUT92), .A2(G104), .A3(G2105), .ZN(new_n800));
  OAI221_X1 g375(.A(G2104), .B1(G116), .B2(new_n463), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n796), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n795), .B1(new_n803), .B2(new_n695), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2067), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n782), .A2(new_n793), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n747), .A2(new_n757), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n726), .A2(new_n727), .A3(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  INV_X1    g386(.A(G55), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n522), .A2(new_n811), .B1(new_n524), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n517), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G860), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT37), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n613), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  INV_X1    g396(.A(new_n816), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n563), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n554), .A2(new_n562), .A3(new_n816), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n821), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT39), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT95), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n817), .B1(new_n827), .B2(KEYINPUT39), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n819), .B1(new_n829), .B2(new_n830), .ZN(G145));
  AND2_X1   g406(.A1(new_n495), .A2(new_n497), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n834));
  AND4_X1   g409(.A1(new_n833), .A2(new_n834), .A3(new_n508), .A4(new_n502), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n833), .B1(new_n506), .B2(new_n508), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n803), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n791), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n778), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n791), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n791), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n779), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n485), .A2(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n463), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  INV_X1    g421(.A(G142), .ZN(new_n847));
  OAI221_X1 g422(.A(new_n844), .B1(new_n845), .B2(new_n846), .C1(new_n491), .C2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n637), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n701), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n840), .A2(new_n843), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n840), .A2(KEYINPUT98), .A3(new_n843), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n840), .A2(new_n843), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n850), .B(KEYINPUT97), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(G162), .B(G160), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n765), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n765), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(KEYINPUT99), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n855), .A2(new_n859), .A3(new_n864), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n840), .A2(new_n857), .A3(new_n843), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(G37), .B1(new_n870), .B2(new_n865), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(KEYINPUT100), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT100), .B1(new_n868), .B2(new_n871), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n868), .A2(new_n871), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT40), .B1(new_n879), .B2(new_n872), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n876), .A2(new_n880), .ZN(G395));
  NAND2_X1  g456(.A1(new_n822), .A2(new_n600), .ZN(new_n882));
  XNOR2_X1  g457(.A(G290), .B(G288), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(G303), .B(G305), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n883), .B2(new_n884), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n622), .B(new_n825), .ZN(new_n894));
  OR2_X1    g469(.A1(G299), .A2(new_n611), .ZN(new_n895));
  NAND2_X1  g470(.A1(G299), .A2(new_n611), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(KEYINPUT41), .A3(new_n896), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n898), .B1(new_n894), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n893), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n882), .B1(new_n904), .B2(new_n600), .ZN(G295));
  OAI21_X1  g480(.A(new_n882), .B1(new_n904), .B2(new_n600), .ZN(G331));
  XNOR2_X1  g481(.A(G301), .B(G168), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n897), .B1(new_n825), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(G171), .A2(G168), .ZN(new_n910));
  NAND2_X1  g485(.A1(G301), .A2(G286), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n823), .A2(new_n910), .A3(new_n824), .A4(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(KEYINPUT104), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n907), .A2(new_n915), .A3(new_n823), .A4(new_n824), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n908), .A2(new_n825), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n902), .A2(new_n919), .A3(KEYINPUT105), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n914), .A2(new_n916), .B1(new_n825), .B2(new_n908), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n900), .A2(new_n901), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI211_X1 g499(.A(new_n891), .B(new_n913), .C1(new_n920), .C2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n918), .B2(new_n912), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n909), .A2(new_n917), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n891), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n913), .B1(new_n920), .B2(new_n924), .ZN(new_n932));
  INV_X1    g507(.A(new_n891), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n931), .B(KEYINPUT44), .C1(new_n934), .C2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  INV_X1    g514(.A(new_n936), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n934), .B2(new_n925), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n935), .A2(new_n929), .A3(new_n928), .A4(new_n936), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI211_X1 g520(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n941), .C2(new_n942), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n938), .B1(new_n945), .B2(new_n946), .ZN(G397));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT45), .B1(new_n837), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT107), .B(G40), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n466), .A2(new_n471), .A3(new_n468), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n471), .B1(new_n466), .B2(new_n468), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n483), .B(new_n950), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT108), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n473), .A2(new_n955), .A3(new_n483), .A4(new_n950), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n949), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1996), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT46), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT123), .Z(new_n962));
  XNOR2_X1  g537(.A(new_n958), .B(KEYINPUT109), .ZN(new_n963));
  INV_X1    g538(.A(G2067), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n802), .B(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n963), .B1(new_n778), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n959), .A2(new_n960), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n971));
  OR3_X1    g546(.A1(new_n962), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n962), .B2(new_n970), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n972), .A2(KEYINPUT124), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT124), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n965), .B1(new_n960), .B2(new_n779), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n963), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n778), .B2(new_n969), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n701), .B(new_n704), .Z(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n979), .B2(new_n963), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n958), .A2(G1986), .A3(G290), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT48), .Z(new_n982));
  AND2_X1   g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n702), .A2(new_n704), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n978), .A2(new_n984), .B1(G2067), .B2(new_n802), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n985), .A2(new_n963), .ZN(new_n986));
  NOR4_X1   g561(.A1(new_n974), .A2(new_n975), .A3(new_n983), .A4(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n954), .A2(new_n956), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT114), .B1(new_n949), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n834), .A2(new_n508), .A3(new_n502), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT96), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n506), .A2(new_n833), .A3(new_n508), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n994), .B2(new_n832), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n990), .B(new_n957), .C1(new_n995), .C2(KEYINPUT45), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(G1384), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(G164), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n989), .A2(new_n996), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1966), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n837), .A2(new_n1005), .A3(new_n948), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n991), .A2(new_n832), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n948), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1008), .A2(KEYINPUT50), .B1(new_n954), .B2(new_n956), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT115), .B(G2084), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1006), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1004), .A2(G168), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(G8), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1011), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(G168), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT51), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  AOI211_X1 g593(.A(KEYINPUT51), .B(new_n1018), .C1(new_n1015), .C2(G168), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT62), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1018), .B1(new_n1015), .B2(G168), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n837), .A2(new_n948), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n988), .B1(new_n1025), .B2(new_n997), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1000), .B1(new_n1026), .B2(new_n990), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1966), .B1(new_n1027), .B2(new_n989), .ZN(new_n1028));
  OAI21_X1  g603(.A(G286), .B1(new_n1028), .B2(new_n1011), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1023), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT62), .B1(new_n1030), .B2(new_n1019), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n957), .A2(new_n837), .A3(new_n948), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n710), .A2(G1976), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(G8), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n589), .B2(new_n592), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n588), .A2(new_n591), .A3(G1981), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1037), .A2(new_n1038), .B1(KEYINPUT113), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(KEYINPUT49), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT113), .B(new_n1039), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1032), .A3(G8), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1035), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1032), .A2(G8), .A3(new_n1033), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1045), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G303), .A2(G8), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT55), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n997), .B1(G164), .B2(G1384), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n957), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n498), .B1(new_n992), .B2(new_n993), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n999), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT110), .B1(new_n837), .B2(new_n998), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1971), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1005), .B1(new_n837), .B2(new_n948), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1384), .B1(new_n991), .B2(new_n832), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1005), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n957), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT111), .B(G2090), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1061), .A2(new_n1062), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1054), .B1(new_n1069), .B2(new_n1018), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1054), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n957), .A2(new_n1055), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1058), .B1(new_n1057), .B2(new_n999), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n837), .A2(KEYINPUT110), .A3(new_n998), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(G1971), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1068), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(G8), .B(new_n1071), .C1(new_n1076), .C2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1052), .A2(new_n1070), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1061), .B2(G2078), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1077), .A2(new_n753), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(G2078), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n989), .A2(new_n996), .A3(new_n1001), .A4(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G171), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1081), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1022), .A2(new_n1031), .A3(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1044), .A2(new_n1046), .A3(new_n710), .ZN(new_n1091));
  OAI211_X1 g666(.A(G8), .B(new_n1032), .C1(new_n1091), .C2(new_n1038), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1052), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(new_n1080), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT63), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1015), .A2(new_n1018), .A3(G286), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1095), .B1(new_n1097), .B2(new_n1081), .ZN(new_n1098));
  OAI21_X1  g673(.A(G8), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1095), .B1(new_n1099), .B2(new_n1054), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1096), .A2(new_n1100), .A3(new_n1080), .A4(new_n1052), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1094), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1090), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1105));
  INV_X1    g680(.A(new_n949), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1085), .A2(G40), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(G160), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1083), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT120), .B1(new_n1077), .B2(new_n753), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1111), .B(G1961), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT121), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1084), .A2(new_n1111), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1077), .A2(KEYINPUT120), .A3(new_n753), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n1083), .A4(new_n1108), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1114), .A2(G171), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1087), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(G301), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1117), .A2(G301), .A3(new_n1083), .A4(new_n1108), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1088), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1081), .B1(new_n1126), .B2(new_n1121), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1104), .A2(KEYINPUT122), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT118), .B(G1996), .Z(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1056), .B(new_n1130), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT58), .B(G1341), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n1032), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1032), .A2(KEYINPUT119), .A3(new_n1132), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1131), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n564), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT59), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1140), .A3(new_n564), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT56), .B(G2072), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1061), .A2(new_n1145), .B1(new_n1067), .B2(G1956), .ZN(new_n1146));
  OR2_X1    g721(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n573), .A2(new_n575), .A3(new_n580), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n956), .A2(new_n954), .B1(new_n1064), .B2(new_n1005), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n995), .B2(new_n1005), .ZN(new_n1154));
  INV_X1    g729(.A(G1956), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1075), .A2(new_n1144), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(new_n1150), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1143), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n1156), .B2(new_n1150), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1143), .B1(new_n1156), .B2(new_n1150), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1146), .A2(new_n1151), .A3(KEYINPUT117), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n995), .A2(new_n964), .A3(new_n957), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(G1348), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n612), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1077), .A2(new_n730), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1168), .A2(new_n611), .A3(new_n1164), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n611), .A2(KEYINPUT60), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1170), .A2(KEYINPUT60), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1142), .A2(new_n1158), .A3(new_n1163), .A4(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1160), .A2(new_n1162), .A3(new_n1167), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n1151), .B2(new_n1146), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1127), .B(new_n1124), .C1(new_n1030), .C2(new_n1019), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1103), .B1(new_n1128), .B2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(G290), .B(G1986), .Z(new_n1182));
  OAI21_X1  g757(.A(new_n980), .B1(new_n958), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n987), .B1(new_n1181), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g759(.A1(new_n879), .A2(new_n872), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n670), .A2(G319), .ZN(new_n1187));
  XNOR2_X1  g761(.A(new_n1187), .B(KEYINPUT125), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1188), .A2(new_n656), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n1190));
  XNOR2_X1  g764(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  AND2_X1   g765(.A1(new_n688), .A2(new_n689), .ZN(new_n1192));
  NOR2_X1   g766(.A1(new_n688), .A2(new_n689), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n690), .A2(KEYINPUT127), .A3(new_n1191), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AND3_X1   g772(.A1(new_n1186), .A2(new_n943), .A3(new_n1198), .ZN(G308));
  NAND3_X1  g773(.A1(new_n1186), .A2(new_n1198), .A3(new_n943), .ZN(G225));
endmodule


