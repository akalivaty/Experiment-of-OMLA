

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U552 ( .A(KEYINPUT15), .B(n608), .Z(n1000) );
  XNOR2_X2 U553 ( .A(n611), .B(n610), .ZN(n743) );
  NOR2_X1 U554 ( .A1(n538), .A2(n537), .ZN(n609) );
  AND2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n541) );
  NOR2_X2 U556 ( .A1(n609), .A2(G1384), .ZN(n611) );
  BUF_X2 U557 ( .A(n541), .Z(n896) );
  NOR2_X1 U558 ( .A1(n533), .A2(G2104), .ZN(n528) );
  XNOR2_X1 U559 ( .A(n700), .B(KEYINPUT64), .ZN(n702) );
  NAND2_X1 U560 ( .A1(n541), .A2(G113), .ZN(n542) );
  AND2_X1 U561 ( .A1(n646), .A2(n619), .ZN(n620) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n652) );
  INV_X1 U563 ( .A(KEYINPUT103), .ZN(n659) );
  XOR2_X1 U564 ( .A(KEYINPUT107), .B(n714), .Z(n715) );
  NOR2_X2 U565 ( .A1(n582), .A2(n522), .ZN(n803) );
  BUF_X1 U566 ( .A(n730), .Z(n904) );
  INV_X1 U567 ( .A(KEYINPUT68), .ZN(n545) );
  BUF_X1 U568 ( .A(n612), .Z(G160) );
  OR2_X1 U569 ( .A1(G301), .A2(n668), .ZN(n517) );
  XOR2_X1 U570 ( .A(KEYINPUT27), .B(KEYINPUT99), .Z(n616) );
  NOR2_X1 U571 ( .A1(n639), .A2(n638), .ZN(n642) );
  INV_X1 U572 ( .A(n661), .ZN(n654) );
  INV_X1 U573 ( .A(G168), .ZN(n666) );
  INV_X1 U574 ( .A(KEYINPUT31), .ZN(n671) );
  AND2_X1 U575 ( .A1(n683), .A2(n676), .ZN(n677) );
  INV_X1 U576 ( .A(KEYINPUT32), .ZN(n691) );
  XNOR2_X1 U577 ( .A(n692), .B(n691), .ZN(n693) );
  INV_X1 U578 ( .A(n986), .ZN(n705) );
  INV_X1 U579 ( .A(n720), .ZN(n698) );
  NOR2_X1 U580 ( .A1(n703), .A2(n695), .ZN(n990) );
  INV_X1 U581 ( .A(KEYINPUT33), .ZN(n701) );
  INV_X1 U582 ( .A(KEYINPUT65), .ZN(n610) );
  NAND2_X1 U583 ( .A1(n811), .A2(G66), .ZN(n603) );
  INV_X1 U584 ( .A(G2105), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n532), .A2(n533), .ZN(n534) );
  INV_X1 U586 ( .A(KEYINPUT1), .ZN(n518) );
  NOR2_X1 U587 ( .A1(G651), .A2(G543), .ZN(n804) );
  NOR2_X2 U588 ( .A1(G2105), .A2(n532), .ZN(n901) );
  NOR2_X2 U589 ( .A1(n630), .A2(n629), .ZN(n998) );
  NOR2_X1 U590 ( .A1(n551), .A2(n550), .ZN(n612) );
  XOR2_X1 U591 ( .A(G543), .B(KEYINPUT0), .Z(n582) );
  NOR2_X2 U592 ( .A1(G651), .A2(n582), .ZN(n807) );
  NAND2_X1 U593 ( .A1(G52), .A2(n807), .ZN(n521) );
  INV_X1 U594 ( .A(G651), .ZN(n522) );
  NOR2_X1 U595 ( .A1(G543), .A2(n522), .ZN(n519) );
  XNOR2_X2 U596 ( .A(n519), .B(n518), .ZN(n811) );
  NAND2_X1 U597 ( .A1(G64), .A2(n811), .ZN(n520) );
  NAND2_X1 U598 ( .A1(n521), .A2(n520), .ZN(n527) );
  NAND2_X1 U599 ( .A1(G77), .A2(n803), .ZN(n524) );
  NAND2_X1 U600 ( .A1(G90), .A2(n804), .ZN(n523) );
  NAND2_X1 U601 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U602 ( .A(KEYINPUT9), .B(n525), .Z(n526) );
  NOR2_X1 U603 ( .A1(n527), .A2(n526), .ZN(G171) );
  INV_X1 U604 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U605 ( .A(n528), .B(KEYINPUT66), .ZN(n540) );
  NAND2_X1 U606 ( .A1(n540), .A2(G126), .ZN(n530) );
  NAND2_X1 U607 ( .A1(n896), .A2(G114), .ZN(n529) );
  NAND2_X1 U608 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U609 ( .A(n531), .B(KEYINPUT88), .ZN(n538) );
  INV_X1 U610 ( .A(G2104), .ZN(n532) );
  NAND2_X1 U611 ( .A1(G102), .A2(n901), .ZN(n536) );
  XNOR2_X2 U612 ( .A(n534), .B(KEYINPUT17), .ZN(n730) );
  NAND2_X1 U613 ( .A1(G138), .A2(n730), .ZN(n535) );
  NAND2_X1 U614 ( .A1(n536), .A2(n535), .ZN(n537) );
  BUF_X1 U615 ( .A(n609), .Z(G164) );
  BUF_X1 U616 ( .A(n540), .Z(n897) );
  NAND2_X1 U617 ( .A1(G125), .A2(n897), .ZN(n548) );
  NAND2_X1 U618 ( .A1(n730), .A2(G137), .ZN(n544) );
  XOR2_X1 U619 ( .A(KEYINPUT67), .B(n542), .Z(n543) );
  NAND2_X1 U620 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U621 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U622 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U623 ( .A1(G101), .A2(n901), .ZN(n549) );
  XNOR2_X1 U624 ( .A(KEYINPUT23), .B(n549), .ZN(n550) );
  NAND2_X1 U625 ( .A1(G91), .A2(n804), .ZN(n553) );
  NAND2_X1 U626 ( .A1(G65), .A2(n811), .ZN(n552) );
  NAND2_X1 U627 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U628 ( .A1(G78), .A2(n803), .ZN(n555) );
  NAND2_X1 U629 ( .A1(G53), .A2(n807), .ZN(n554) );
  NAND2_X1 U630 ( .A1(n555), .A2(n554), .ZN(n556) );
  OR2_X1 U631 ( .A1(n557), .A2(n556), .ZN(G299) );
  XOR2_X1 U632 ( .A(KEYINPUT4), .B(KEYINPUT74), .Z(n559) );
  NAND2_X1 U633 ( .A1(G89), .A2(n804), .ZN(n558) );
  XNOR2_X1 U634 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U635 ( .A(KEYINPUT73), .B(n560), .ZN(n562) );
  NAND2_X1 U636 ( .A1(n803), .A2(G76), .ZN(n561) );
  NAND2_X1 U637 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U638 ( .A(n563), .B(KEYINPUT5), .ZN(n569) );
  XNOR2_X1 U639 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n567) );
  NAND2_X1 U640 ( .A1(G51), .A2(n807), .ZN(n565) );
  NAND2_X1 U641 ( .A1(G63), .A2(n811), .ZN(n564) );
  NAND2_X1 U642 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U643 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U644 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U645 ( .A(KEYINPUT7), .B(n570), .ZN(G168) );
  XOR2_X1 U646 ( .A(G168), .B(KEYINPUT8), .Z(n571) );
  XNOR2_X1 U647 ( .A(KEYINPUT76), .B(n571), .ZN(G286) );
  NAND2_X1 U648 ( .A1(G75), .A2(n803), .ZN(n573) );
  NAND2_X1 U649 ( .A1(G88), .A2(n804), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U651 ( .A1(G50), .A2(n807), .ZN(n575) );
  NAND2_X1 U652 ( .A1(G62), .A2(n811), .ZN(n574) );
  NAND2_X1 U653 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U654 ( .A1(n577), .A2(n576), .ZN(G166) );
  INV_X1 U655 ( .A(G166), .ZN(G303) );
  NAND2_X1 U656 ( .A1(G49), .A2(n807), .ZN(n579) );
  NAND2_X1 U657 ( .A1(G74), .A2(G651), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U659 ( .A(KEYINPUT81), .B(n580), .Z(n581) );
  NOR2_X1 U660 ( .A1(n811), .A2(n581), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n582), .A2(G87), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(G288) );
  XOR2_X1 U663 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n586) );
  NAND2_X1 U664 ( .A1(G73), .A2(n803), .ZN(n585) );
  XNOR2_X1 U665 ( .A(n586), .B(n585), .ZN(n590) );
  NAND2_X1 U666 ( .A1(G86), .A2(n804), .ZN(n588) );
  NAND2_X1 U667 ( .A1(G61), .A2(n811), .ZN(n587) );
  NAND2_X1 U668 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U669 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n807), .A2(G48), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n592), .A2(n591), .ZN(G305) );
  NAND2_X1 U672 ( .A1(G72), .A2(n803), .ZN(n594) );
  NAND2_X1 U673 ( .A1(G85), .A2(n804), .ZN(n593) );
  NAND2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U675 ( .A1(G60), .A2(n811), .ZN(n595) );
  XNOR2_X1 U676 ( .A(KEYINPUT69), .B(n595), .ZN(n596) );
  NOR2_X1 U677 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n807), .A2(G47), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(G290) );
  NAND2_X1 U680 ( .A1(G92), .A2(n804), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n600), .B(KEYINPUT72), .ZN(n607) );
  NAND2_X1 U682 ( .A1(G79), .A2(n803), .ZN(n602) );
  NAND2_X1 U683 ( .A1(G54), .A2(n807), .ZN(n601) );
  NAND2_X1 U684 ( .A1(n602), .A2(n601), .ZN(n605) );
  XNOR2_X1 U685 ( .A(KEYINPUT71), .B(n603), .ZN(n604) );
  NOR2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n612), .A2(G40), .ZN(n744) );
  INV_X1 U689 ( .A(n744), .ZN(n613) );
  NAND2_X2 U690 ( .A1(n743), .A2(n613), .ZN(n661) );
  BUF_X2 U691 ( .A(n661), .Z(n663) );
  NAND2_X1 U692 ( .A1(G1348), .A2(n663), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G2067), .A2(n654), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n640) );
  NOR2_X1 U695 ( .A1(n1000), .A2(n640), .ZN(n621) );
  INV_X1 U696 ( .A(G2072), .ZN(n932) );
  NOR2_X2 U697 ( .A1(n661), .A2(n932), .ZN(n617) );
  XNOR2_X1 U698 ( .A(n617), .B(n616), .ZN(n646) );
  NAND2_X1 U699 ( .A1(n661), .A2(G1956), .ZN(n647) );
  INV_X1 U700 ( .A(G299), .ZN(n618) );
  AND2_X1 U701 ( .A1(n647), .A2(n618), .ZN(n619) );
  NOR2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n644) );
  NAND2_X1 U703 ( .A1(n804), .A2(G81), .ZN(n622) );
  XNOR2_X1 U704 ( .A(n622), .B(KEYINPUT12), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G68), .A2(n803), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U707 ( .A(n625), .B(KEYINPUT13), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G43), .A2(n807), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n811), .A2(G56), .ZN(n628) );
  XOR2_X1 U711 ( .A(KEYINPUT14), .B(n628), .Z(n629) );
  XOR2_X1 U712 ( .A(G1996), .B(KEYINPUT100), .Z(n972) );
  XNOR2_X1 U713 ( .A(KEYINPUT26), .B(KEYINPUT101), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n972), .A2(n632), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n998), .A2(n631), .ZN(n639) );
  INV_X1 U716 ( .A(G1341), .ZN(n1017) );
  INV_X1 U717 ( .A(n632), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n1017), .A2(n634), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n633), .A2(n663), .ZN(n637) );
  NOR2_X1 U720 ( .A1(n972), .A2(n661), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n640), .A2(n1000), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n645), .B(KEYINPUT102), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n646), .A2(n647), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n648), .A2(G299), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n649), .B(KEYINPUT28), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n658) );
  XNOR2_X1 U732 ( .A(G1961), .B(KEYINPUT97), .ZN(n1026) );
  NAND2_X1 U733 ( .A1(n663), .A2(n1026), .ZN(n656) );
  XNOR2_X1 U734 ( .A(KEYINPUT25), .B(G2078), .ZN(n963) );
  NAND2_X1 U735 ( .A1(n654), .A2(n963), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U737 ( .A(n657), .B(KEYINPUT98), .Z(n668) );
  NAND2_X1 U738 ( .A1(n658), .A2(n517), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n660), .B(n659), .ZN(n674) );
  NOR2_X2 U740 ( .A1(G2084), .A2(n661), .ZN(n678) );
  XOR2_X1 U741 ( .A(KEYINPUT96), .B(n678), .Z(n662) );
  NAND2_X1 U742 ( .A1(G8), .A2(n662), .ZN(n664) );
  NAND2_X1 U743 ( .A1(G8), .A2(n663), .ZN(n720) );
  NOR2_X1 U744 ( .A1(G1966), .A2(n720), .ZN(n675) );
  NOR2_X1 U745 ( .A1(n664), .A2(n675), .ZN(n665) );
  XNOR2_X1 U746 ( .A(n665), .B(KEYINPUT30), .ZN(n667) );
  AND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(n670) );
  AND2_X1 U748 ( .A1(G301), .A2(n668), .ZN(n669) );
  NOR2_X1 U749 ( .A1(n670), .A2(n669), .ZN(n672) );
  XNOR2_X1 U750 ( .A(n672), .B(n671), .ZN(n673) );
  NAND2_X1 U751 ( .A1(n674), .A2(n673), .ZN(n683) );
  INV_X1 U752 ( .A(n675), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n677), .B(KEYINPUT104), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n678), .B(KEYINPUT96), .ZN(n679) );
  NAND2_X1 U755 ( .A1(G8), .A2(n679), .ZN(n680) );
  NAND2_X1 U756 ( .A1(n681), .A2(n680), .ZN(n694) );
  AND2_X1 U757 ( .A1(G286), .A2(G8), .ZN(n682) );
  NAND2_X1 U758 ( .A1(n683), .A2(n682), .ZN(n690) );
  INV_X1 U759 ( .A(G8), .ZN(n688) );
  NOR2_X1 U760 ( .A1(G2090), .A2(n663), .ZN(n685) );
  NOR2_X1 U761 ( .A1(G1971), .A2(n720), .ZN(n684) );
  NOR2_X1 U762 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U763 ( .A1(n686), .A2(G303), .ZN(n687) );
  OR2_X1 U764 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U765 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n711) );
  NOR2_X1 U767 ( .A1(G1976), .A2(G288), .ZN(n703) );
  NOR2_X1 U768 ( .A1(G1971), .A2(G303), .ZN(n695) );
  NAND2_X1 U769 ( .A1(n711), .A2(n990), .ZN(n696) );
  NAND2_X1 U770 ( .A1(G1976), .A2(G288), .ZN(n989) );
  NAND2_X1 U771 ( .A1(n696), .A2(n989), .ZN(n697) );
  XNOR2_X1 U772 ( .A(n697), .B(KEYINPUT105), .ZN(n699) );
  NAND2_X1 U773 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U774 ( .A1(n702), .A2(n701), .ZN(n708) );
  NAND2_X1 U775 ( .A1(n703), .A2(KEYINPUT33), .ZN(n704) );
  NOR2_X1 U776 ( .A1(n720), .A2(n704), .ZN(n706) );
  XOR2_X1 U777 ( .A(G1981), .B(G305), .Z(n986) );
  NOR2_X1 U778 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n716) );
  NOR2_X1 U780 ( .A1(G2090), .A2(G303), .ZN(n709) );
  NAND2_X1 U781 ( .A1(G8), .A2(n709), .ZN(n710) );
  XNOR2_X1 U782 ( .A(n710), .B(KEYINPUT106), .ZN(n712) );
  NAND2_X1 U783 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n713), .A2(n720), .ZN(n714) );
  NAND2_X1 U785 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U786 ( .A(n717), .B(KEYINPUT108), .ZN(n722) );
  NOR2_X1 U787 ( .A1(G1981), .A2(G305), .ZN(n718) );
  XOR2_X1 U788 ( .A(n718), .B(KEYINPUT24), .Z(n719) );
  NOR2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X2 U790 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U791 ( .A(n723), .B(KEYINPUT109), .ZN(n761) );
  NAND2_X1 U792 ( .A1(n896), .A2(G117), .ZN(n725) );
  NAND2_X1 U793 ( .A1(G129), .A2(n897), .ZN(n724) );
  NAND2_X1 U794 ( .A1(n725), .A2(n724), .ZN(n729) );
  NAND2_X1 U795 ( .A1(G105), .A2(n901), .ZN(n726) );
  XNOR2_X1 U796 ( .A(n726), .B(KEYINPUT95), .ZN(n727) );
  XNOR2_X1 U797 ( .A(n727), .B(KEYINPUT38), .ZN(n728) );
  NOR2_X1 U798 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U799 ( .A1(n904), .A2(G141), .ZN(n731) );
  NAND2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n878) );
  NAND2_X1 U801 ( .A1(n878), .A2(G1996), .ZN(n742) );
  NAND2_X1 U802 ( .A1(G95), .A2(n901), .ZN(n734) );
  NAND2_X1 U803 ( .A1(G131), .A2(n904), .ZN(n733) );
  NAND2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U805 ( .A(KEYINPUT94), .B(n735), .ZN(n738) );
  NAND2_X1 U806 ( .A1(G107), .A2(n896), .ZN(n736) );
  XNOR2_X1 U807 ( .A(KEYINPUT93), .B(n736), .ZN(n737) );
  NOR2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U809 ( .A1(G119), .A2(n897), .ZN(n739) );
  NAND2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n879) );
  NAND2_X1 U811 ( .A1(n879), .A2(G1991), .ZN(n741) );
  NAND2_X1 U812 ( .A1(n742), .A2(n741), .ZN(n943) );
  NOR2_X1 U813 ( .A1(n743), .A2(n744), .ZN(n773) );
  AND2_X1 U814 ( .A1(n943), .A2(n773), .ZN(n764) );
  XNOR2_X1 U815 ( .A(G1986), .B(G290), .ZN(n997) );
  NAND2_X1 U816 ( .A1(n773), .A2(n997), .ZN(n745) );
  XNOR2_X1 U817 ( .A(KEYINPUT89), .B(n745), .ZN(n746) );
  NOR2_X1 U818 ( .A1(n764), .A2(n746), .ZN(n759) );
  XNOR2_X1 U819 ( .A(KEYINPUT34), .B(KEYINPUT90), .ZN(n750) );
  NAND2_X1 U820 ( .A1(G104), .A2(n901), .ZN(n748) );
  NAND2_X1 U821 ( .A1(G140), .A2(n904), .ZN(n747) );
  NAND2_X1 U822 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U823 ( .A(n750), .B(n749), .ZN(n756) );
  XNOR2_X1 U824 ( .A(KEYINPUT35), .B(KEYINPUT91), .ZN(n754) );
  NAND2_X1 U825 ( .A1(n896), .A2(G116), .ZN(n752) );
  NAND2_X1 U826 ( .A1(G128), .A2(n897), .ZN(n751) );
  NAND2_X1 U827 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U828 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U830 ( .A(n757), .B(KEYINPUT36), .ZN(n758) );
  XNOR2_X1 U831 ( .A(n758), .B(KEYINPUT92), .ZN(n893) );
  XNOR2_X1 U832 ( .A(G2067), .B(KEYINPUT37), .ZN(n769) );
  NOR2_X1 U833 ( .A1(n893), .A2(n769), .ZN(n951) );
  NAND2_X1 U834 ( .A1(n773), .A2(n951), .ZN(n767) );
  AND2_X1 U835 ( .A1(n759), .A2(n767), .ZN(n760) );
  NAND2_X1 U836 ( .A1(n761), .A2(n760), .ZN(n775) );
  NOR2_X1 U837 ( .A1(G1996), .A2(n878), .ZN(n940) );
  NOR2_X1 U838 ( .A1(G1986), .A2(G290), .ZN(n762) );
  NOR2_X1 U839 ( .A1(G1991), .A2(n879), .ZN(n947) );
  NOR2_X1 U840 ( .A1(n762), .A2(n947), .ZN(n763) );
  NOR2_X1 U841 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U842 ( .A1(n940), .A2(n765), .ZN(n766) );
  XNOR2_X1 U843 ( .A(KEYINPUT39), .B(n766), .ZN(n768) );
  NAND2_X1 U844 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n769), .A2(n893), .ZN(n770) );
  XNOR2_X1 U846 ( .A(n770), .B(KEYINPUT110), .ZN(n937) );
  NAND2_X1 U847 ( .A1(n771), .A2(n937), .ZN(n772) );
  NAND2_X1 U848 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U849 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U850 ( .A(n776), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U851 ( .A1(G123), .A2(n897), .ZN(n778) );
  XNOR2_X1 U852 ( .A(KEYINPUT78), .B(KEYINPUT18), .ZN(n777) );
  XNOR2_X1 U853 ( .A(n778), .B(n777), .ZN(n785) );
  NAND2_X1 U854 ( .A1(G111), .A2(n896), .ZN(n780) );
  NAND2_X1 U855 ( .A1(G99), .A2(n901), .ZN(n779) );
  NAND2_X1 U856 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U857 ( .A1(G135), .A2(n904), .ZN(n781) );
  XNOR2_X1 U858 ( .A(KEYINPUT79), .B(n781), .ZN(n782) );
  NOR2_X1 U859 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U860 ( .A1(n785), .A2(n784), .ZN(n948) );
  XNOR2_X1 U861 ( .A(G2096), .B(n948), .ZN(n786) );
  OR2_X1 U862 ( .A1(G2100), .A2(n786), .ZN(G156) );
  INV_X1 U863 ( .A(G132), .ZN(G219) );
  INV_X1 U864 ( .A(G82), .ZN(G220) );
  INV_X1 U865 ( .A(G57), .ZN(G237) );
  NAND2_X1 U866 ( .A1(G94), .A2(G452), .ZN(n787) );
  XOR2_X1 U867 ( .A(KEYINPUT70), .B(n787), .Z(G173) );
  NAND2_X1 U868 ( .A1(G7), .A2(G661), .ZN(n788) );
  XNOR2_X1 U869 ( .A(n788), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U870 ( .A(G223), .ZN(n844) );
  NAND2_X1 U871 ( .A1(n844), .A2(G567), .ZN(n789) );
  XOR2_X1 U872 ( .A(KEYINPUT11), .B(n789), .Z(G234) );
  NAND2_X1 U873 ( .A1(n998), .A2(G860), .ZN(G153) );
  NAND2_X1 U874 ( .A1(G868), .A2(G301), .ZN(n791) );
  INV_X1 U875 ( .A(G868), .ZN(n826) );
  NAND2_X1 U876 ( .A1(n1000), .A2(n826), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(G284) );
  NOR2_X1 U878 ( .A1(G868), .A2(G299), .ZN(n792) );
  XOR2_X1 U879 ( .A(KEYINPUT77), .B(n792), .Z(n794) );
  NOR2_X1 U880 ( .A1(G286), .A2(n826), .ZN(n793) );
  NOR2_X1 U881 ( .A1(n794), .A2(n793), .ZN(G297) );
  INV_X1 U882 ( .A(G860), .ZN(n795) );
  NAND2_X1 U883 ( .A1(n795), .A2(G559), .ZN(n796) );
  INV_X1 U884 ( .A(n1000), .ZN(n801) );
  NAND2_X1 U885 ( .A1(n796), .A2(n801), .ZN(n797) );
  XNOR2_X1 U886 ( .A(n797), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U887 ( .A1(n801), .A2(G868), .ZN(n798) );
  NOR2_X1 U888 ( .A1(G559), .A2(n798), .ZN(n800) );
  AND2_X1 U889 ( .A1(n826), .A2(n998), .ZN(n799) );
  NOR2_X1 U890 ( .A1(n800), .A2(n799), .ZN(G282) );
  NAND2_X1 U891 ( .A1(n801), .A2(G559), .ZN(n823) );
  XOR2_X1 U892 ( .A(n998), .B(n823), .Z(n802) );
  NOR2_X1 U893 ( .A1(G860), .A2(n802), .ZN(n814) );
  NAND2_X1 U894 ( .A1(G80), .A2(n803), .ZN(n806) );
  NAND2_X1 U895 ( .A1(G93), .A2(n804), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n807), .A2(G55), .ZN(n808) );
  XOR2_X1 U898 ( .A(KEYINPUT80), .B(n808), .Z(n809) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n811), .A2(G67), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n825) );
  XOR2_X1 U902 ( .A(n814), .B(n825), .Z(G145) );
  XOR2_X1 U903 ( .A(G305), .B(G299), .Z(n818) );
  XOR2_X1 U904 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n816) );
  XNOR2_X1 U905 ( .A(G166), .B(KEYINPUT19), .ZN(n815) );
  XNOR2_X1 U906 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U907 ( .A(n818), .B(n817), .ZN(n820) );
  XNOR2_X1 U908 ( .A(G288), .B(n998), .ZN(n819) );
  XNOR2_X1 U909 ( .A(n820), .B(n819), .ZN(n821) );
  XNOR2_X1 U910 ( .A(n821), .B(G290), .ZN(n822) );
  XNOR2_X1 U911 ( .A(n822), .B(n825), .ZN(n912) );
  XNOR2_X1 U912 ( .A(n823), .B(n912), .ZN(n824) );
  NAND2_X1 U913 ( .A1(n824), .A2(G868), .ZN(n828) );
  NAND2_X1 U914 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U915 ( .A1(n828), .A2(n827), .ZN(G295) );
  NAND2_X1 U916 ( .A1(G2084), .A2(G2078), .ZN(n829) );
  XOR2_X1 U917 ( .A(KEYINPUT20), .B(n829), .Z(n830) );
  NAND2_X1 U918 ( .A1(G2090), .A2(n830), .ZN(n831) );
  XNOR2_X1 U919 ( .A(KEYINPUT21), .B(n831), .ZN(n832) );
  NAND2_X1 U920 ( .A1(n832), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U921 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U922 ( .A1(G120), .A2(G69), .ZN(n833) );
  NOR2_X1 U923 ( .A1(G237), .A2(n833), .ZN(n834) );
  XNOR2_X1 U924 ( .A(KEYINPUT86), .B(n834), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n835), .A2(G108), .ZN(n848) );
  NAND2_X1 U926 ( .A1(n848), .A2(G567), .ZN(n841) );
  NOR2_X1 U927 ( .A1(G220), .A2(G219), .ZN(n836) );
  XOR2_X1 U928 ( .A(KEYINPUT22), .B(n836), .Z(n837) );
  NOR2_X1 U929 ( .A1(G218), .A2(n837), .ZN(n838) );
  NAND2_X1 U930 ( .A1(G96), .A2(n838), .ZN(n849) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n849), .ZN(n839) );
  XOR2_X1 U932 ( .A(KEYINPUT85), .B(n839), .Z(n840) );
  NAND2_X1 U933 ( .A1(n841), .A2(n840), .ZN(n851) );
  NAND2_X1 U934 ( .A1(G483), .A2(G661), .ZN(n842) );
  NOR2_X1 U935 ( .A1(n851), .A2(n842), .ZN(n843) );
  XOR2_X1 U936 ( .A(KEYINPUT87), .B(n843), .Z(n847) );
  NAND2_X1 U937 ( .A1(n847), .A2(G36), .ZN(G176) );
  NAND2_X1 U938 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U940 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n847), .A2(n846), .ZN(G188) );
  XOR2_X1 U943 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  INV_X1 U945 ( .A(G120), .ZN(G236) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  INV_X1 U947 ( .A(G69), .ZN(G235) );
  NOR2_X1 U948 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n850), .B(KEYINPUT111), .ZN(G261) );
  INV_X1 U950 ( .A(G261), .ZN(G325) );
  INV_X1 U951 ( .A(n851), .ZN(G319) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT43), .Z(n853) );
  XNOR2_X1 U953 ( .A(G2090), .B(KEYINPUT112), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n854), .B(G2678), .Z(n856) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2100), .Z(n858) );
  XNOR2_X1 U959 ( .A(G2084), .B(G2078), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U962 ( .A(G1956), .B(G1966), .Z(n862) );
  XNOR2_X1 U963 ( .A(G1986), .B(G1981), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U965 ( .A(G1971), .B(G1976), .Z(n864) );
  XNOR2_X1 U966 ( .A(G1996), .B(G1991), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U969 ( .A(KEYINPUT113), .B(G2474), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(n870) );
  XOR2_X1 U971 ( .A(G1961), .B(KEYINPUT41), .Z(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(G229) );
  NAND2_X1 U973 ( .A1(G112), .A2(n896), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G100), .A2(n901), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G124), .A2(n897), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U978 ( .A1(G136), .A2(n904), .ZN(n874) );
  NAND2_X1 U979 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U980 ( .A1(n877), .A2(n876), .ZN(G162) );
  XNOR2_X1 U981 ( .A(KEYINPUT48), .B(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U983 ( .A(n881), .B(KEYINPUT46), .Z(n891) );
  NAND2_X1 U984 ( .A1(n896), .A2(G118), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G130), .A2(n897), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G106), .A2(n901), .ZN(n885) );
  NAND2_X1 U988 ( .A1(G142), .A2(n904), .ZN(n884) );
  NAND2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U990 ( .A(KEYINPUT45), .B(n886), .Z(n887) );
  NOR2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U992 ( .A(G160), .B(n889), .ZN(n890) );
  XNOR2_X1 U993 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U994 ( .A(n948), .B(n892), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n893), .B(G162), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n895), .B(n894), .ZN(n909) );
  NAND2_X1 U997 ( .A1(n896), .A2(G115), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G127), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n900), .B(KEYINPUT47), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(G103), .A2(n901), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(n904), .A2(G139), .ZN(n905) );
  XOR2_X1 U1004 ( .A(KEYINPUT114), .B(n905), .Z(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n931) );
  XNOR2_X1 U1006 ( .A(G164), .B(n931), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(n911) );
  XOR2_X1 U1009 ( .A(KEYINPUT115), .B(n911), .Z(G395) );
  XNOR2_X1 U1010 ( .A(n912), .B(n1000), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n913), .B(G286), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n914), .B(G171), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n915), .ZN(G397) );
  XOR2_X1 U1014 ( .A(G2451), .B(G2430), .Z(n917) );
  XNOR2_X1 U1015 ( .A(G2438), .B(G2443), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n923) );
  XOR2_X1 U1017 ( .A(G2435), .B(G2454), .Z(n919) );
  XNOR2_X1 U1018 ( .A(G1348), .B(G1341), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(n919), .B(n918), .ZN(n921) );
  XOR2_X1 U1020 ( .A(G2446), .B(G2427), .Z(n920) );
  XNOR2_X1 U1021 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1022 ( .A(n923), .B(n922), .Z(n924) );
  NAND2_X1 U1023 ( .A1(G14), .A2(n924), .ZN(n930) );
  NAND2_X1 U1024 ( .A1(G319), .A2(n930), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1030 ( .A(G225), .ZN(G308) );
  INV_X1 U1031 ( .A(n930), .ZN(G401) );
  XOR2_X1 U1032 ( .A(G164), .B(G2078), .Z(n934) );
  XNOR2_X1 U1033 ( .A(n932), .B(n931), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(n935), .B(KEYINPUT120), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(n936), .B(KEYINPUT50), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n957) );
  XOR2_X1 U1038 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1040 ( .A(KEYINPUT118), .B(n941), .Z(n942) );
  XNOR2_X1 U1041 ( .A(KEYINPUT51), .B(n942), .ZN(n945) );
  INV_X1 U1042 ( .A(n943), .ZN(n944) );
  NAND2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n954) );
  XOR2_X1 U1044 ( .A(G160), .B(G2084), .Z(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(n952), .B(KEYINPUT117), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(KEYINPUT119), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT52), .B(n958), .ZN(n960) );
  INV_X1 U1053 ( .A(KEYINPUT55), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n961), .A2(G29), .ZN(n962) );
  XOR2_X1 U1056 ( .A(KEYINPUT121), .B(n962), .Z(n1042) );
  XNOR2_X1 U1057 ( .A(G27), .B(n963), .ZN(n971) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G26), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(G33), .B(G2072), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(G28), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(G25), .B(G1991), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(KEYINPUT122), .B(n967), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(G32), .B(n972), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT123), .B(n973), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1069 ( .A(KEYINPUT53), .B(n976), .Z(n979) );
  XOR2_X1 U1070 ( .A(KEYINPUT54), .B(G34), .Z(n977) );
  XNOR2_X1 U1071 ( .A(G2084), .B(n977), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G35), .B(G2090), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(KEYINPUT55), .B(n982), .ZN(n984) );
  INV_X1 U1076 ( .A(G29), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n985), .A2(G11), .ZN(n1040) );
  XNOR2_X1 U1079 ( .A(G16), .B(KEYINPUT56), .ZN(n1010) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G168), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(n988), .B(KEYINPUT57), .ZN(n1008) );
  NAND2_X1 U1083 ( .A1(G303), .A2(G1971), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G299), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(n995), .B(KEYINPUT124), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(G1961), .B(G301), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1341), .B(n998), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(n999), .B(KEYINPUT125), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(G1348), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1038) );
  INV_X1 U1099 ( .A(G16), .ZN(n1036) );
  XOR2_X1 U1100 ( .A(G1976), .B(G23), .Z(n1013) );
  XNOR2_X1 U1101 ( .A(G1986), .B(KEYINPUT127), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(n1011), .B(G24), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(G22), .B(G1971), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1016), .Z(n1033) );
  XNOR2_X1 U1107 ( .A(G19), .B(n1017), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(G1981), .B(G6), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(G20), .B(G1956), .ZN(n1018) );
  NOR2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1024) );
  XOR2_X1 U1112 ( .A(KEYINPUT59), .B(G1348), .Z(n1022) );
  XNOR2_X1 U1113 ( .A(G4), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1115 ( .A(KEYINPUT60), .B(n1025), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(n1026), .B(G5), .ZN(n1027) );
  NAND2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1030) );
  XNOR2_X1 U1118 ( .A(G21), .B(G1966), .ZN(n1029) );
  NOR2_X1 U1119 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1120 ( .A(KEYINPUT126), .B(n1031), .Z(n1032) );
  NOR2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1122 ( .A(KEYINPUT61), .B(n1034), .ZN(n1035) );
  NAND2_X1 U1123 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NAND2_X1 U1126 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XOR2_X1 U1127 ( .A(KEYINPUT62), .B(n1043), .Z(G311) );
  INV_X1 U1128 ( .A(G311), .ZN(G150) );
endmodule

