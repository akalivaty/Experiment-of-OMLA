//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(G227), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(G140), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n194), .B(KEYINPUT77), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n195), .B(G110), .Z(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT78), .B1(new_n197), .B2(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G107), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n200), .B2(G107), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n197), .A3(G104), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n202), .A2(KEYINPUT79), .A3(new_n203), .A4(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n203), .A2(new_n198), .A3(new_n205), .A4(new_n201), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT79), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(G101), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n211));
  INV_X1    g025(.A(new_n207), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT0), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT0), .A3(G128), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n231));
  NAND4_X1  g045(.A1(new_n206), .A2(G101), .A3(new_n209), .A4(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n215), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n200), .A2(G107), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n197), .A2(G104), .ZN(new_n235));
  OAI21_X1  g049(.A(G101), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n207), .B2(G101), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n239), .B(KEYINPUT1), .C1(new_n218), .C2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G128), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n239), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n220), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n217), .A2(new_n219), .A3(new_n244), .A4(G128), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n243), .A2(KEYINPUT69), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n243), .B2(new_n245), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n238), .B(KEYINPUT10), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n233), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT66), .A2(G137), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT66), .A2(G137), .ZN(new_n252));
  OAI211_X1 g066(.A(KEYINPUT11), .B(G134), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G137), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT11), .B1(new_n254), .B2(G134), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G131), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n217), .A2(new_n219), .A3(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT1), .B1(new_n218), .B2(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G128), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n265), .A2(new_n244), .B1(new_n267), .B2(new_n220), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n264), .B1(new_n237), .B2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n202), .A2(new_n213), .A3(new_n203), .A4(new_n205), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n225), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n245), .B1(new_n271), .B2(new_n228), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n270), .A2(KEYINPUT81), .A3(new_n236), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n249), .A2(KEYINPUT82), .A3(new_n263), .A4(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n276), .A2(new_n233), .A3(new_n263), .A4(new_n248), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n276), .A2(new_n233), .A3(new_n248), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n262), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n196), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n196), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n243), .A2(new_n245), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n237), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n274), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n262), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n269), .A2(new_n273), .B1(new_n286), .B2(new_n237), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT12), .B1(new_n291), .B2(new_n263), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n285), .B(new_n293), .C1(new_n277), .C2(new_n280), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n191), .B(new_n189), .C1(new_n284), .C2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT83), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n293), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n281), .A2(new_n298), .A3(new_n196), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n277), .A2(new_n280), .B1(new_n262), .B2(new_n282), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n196), .B2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n301), .A2(KEYINPUT83), .A3(new_n191), .A4(new_n189), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  AOI221_X4 g117(.A(new_n285), .B1(new_n262), .B2(new_n282), .C1(new_n277), .C2(new_n280), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n196), .B1(new_n281), .B2(new_n298), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n189), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G469), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n190), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n286), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n311), .B2(new_n230), .ZN(new_n313));
  INV_X1    g127(.A(G953), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n313), .A2(G224), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n313), .B1(G224), .B2(new_n314), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(G116), .B(G119), .Z(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT2), .B(G113), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n318), .B(new_n319), .Z(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n215), .A2(new_n321), .A3(new_n232), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT84), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT5), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G116), .ZN(new_n326));
  OAI211_X1 g140(.A(G113), .B(new_n326), .C1(new_n318), .C2(new_n324), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n318), .B2(new_n319), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n328), .A2(new_n237), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n215), .A2(new_n330), .A3(new_n321), .A4(new_n232), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n323), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(G110), .B(G122), .Z(new_n333));
  OR2_X1    g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(KEYINPUT85), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT85), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n323), .A2(new_n336), .A3(new_n329), .A4(new_n331), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n333), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT6), .B(new_n334), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n335), .B2(new_n337), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n341), .A2(KEYINPUT86), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT86), .B1(new_n341), .B2(new_n342), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n317), .B(new_n340), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(G210), .B1(G237), .B2(G902), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n347), .A2(KEYINPUT7), .B1(new_n314), .B2(G224), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n347), .B2(KEYINPUT7), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n313), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n316), .A2(KEYINPUT7), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n328), .B(new_n237), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n333), .B(KEYINPUT8), .Z(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n334), .A2(new_n350), .A3(new_n351), .A4(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(new_n189), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n345), .A2(new_n346), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n346), .B1(new_n345), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n310), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n309), .A2(new_n359), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n361));
  XNOR2_X1  g175(.A(G125), .B(G140), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(KEYINPUT16), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(new_n216), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n325), .A2(G128), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n225), .A2(G119), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT24), .B(G110), .Z(new_n369));
  AOI21_X1  g183(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(KEYINPUT23), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(KEYINPUT76), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n371), .B(new_n372), .Z(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G110), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  OAI22_X1  g189(.A1(new_n373), .A2(G110), .B1(new_n368), .B2(new_n369), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n363), .A2(G146), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n362), .A2(new_n216), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n314), .A2(G221), .A3(G234), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT22), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(G137), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n380), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n189), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(KEYINPUT25), .A3(new_n189), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(G234), .B2(new_n189), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n391), .B2(new_n385), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT32), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(G101), .ZN(new_n397));
  INV_X1    g211(.A(G237), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n314), .A3(G210), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n397), .B(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(new_n400), .B(KEYINPUT71), .Z(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n251), .A2(new_n252), .A3(G134), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n256), .A2(G137), .ZN(new_n404));
  OAI21_X1  g218(.A(G131), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n261), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n246), .B2(new_n247), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n262), .A2(new_n230), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n320), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT28), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n410), .A2(KEYINPUT72), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT72), .B1(new_n410), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n227), .A2(KEYINPUT65), .A3(new_n229), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT65), .B1(new_n227), .B2(new_n229), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n243), .A2(new_n245), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n417), .A2(new_n262), .B1(new_n407), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n410), .B1(new_n320), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT28), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n402), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT31), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n417), .A2(new_n262), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n286), .A2(new_n406), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n424), .B(new_n425), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT68), .B1(new_n419), .B2(KEYINPUT30), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n408), .A2(KEYINPUT30), .A3(new_n409), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n321), .A4(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT70), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n410), .A2(new_n433), .A3(new_n400), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n410), .B2(new_n400), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n423), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n410), .A2(new_n400), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT70), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n410), .A2(new_n433), .A3(new_n400), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT31), .A3(new_n431), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n422), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G472), .A2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n395), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n414), .A2(new_n421), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n401), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n441), .A2(KEYINPUT31), .A3(new_n431), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT31), .B1(new_n441), .B2(new_n431), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT32), .A3(new_n444), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n394), .B1(new_n446), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT32), .B1(new_n451), .B2(new_n444), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT73), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n431), .A2(new_n410), .ZN(new_n457));
  INV_X1    g271(.A(new_n400), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT74), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n414), .A2(new_n421), .A3(new_n402), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT29), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n457), .A2(KEYINPUT74), .A3(new_n458), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n413), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n410), .A2(KEYINPUT72), .A3(new_n411), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(KEYINPUT75), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT75), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n412), .B2(new_n413), .ZN(new_n470));
  INV_X1    g284(.A(new_n410), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n320), .B1(new_n408), .B2(new_n409), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT28), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n400), .A2(KEYINPUT29), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n465), .A2(new_n189), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G472), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n393), .B1(new_n456), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G128), .B(G143), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(new_n256), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT88), .ZN(new_n482));
  XNOR2_X1  g296(.A(G116), .B(G122), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n197), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT89), .ZN(new_n485));
  INV_X1    g299(.A(G116), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(KEYINPUT14), .A3(G122), .ZN(new_n487));
  INV_X1    g301(.A(new_n483), .ZN(new_n488));
  OAI211_X1 g302(.A(G107), .B(new_n487), .C1(new_n488), .C2(KEYINPUT14), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n225), .A2(KEYINPUT13), .A3(G143), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n256), .B(new_n491), .C1(KEYINPUT13), .C2(new_n480), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n483), .B(new_n197), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n480), .A2(new_n256), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI22_X1  g309(.A1(new_n482), .A2(new_n490), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n188), .A2(G217), .A3(new_n314), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(KEYINPUT90), .A3(new_n499), .ZN(new_n500));
  OR3_X1    g314(.A1(new_n496), .A2(KEYINPUT90), .A3(new_n497), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n189), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G478), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n502), .B(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n398), .A2(new_n314), .A3(G214), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(G143), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(G131), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n507), .A2(new_n260), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n510), .B(new_n364), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G113), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n200), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT18), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n507), .B1(new_n515), .B2(new_n260), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n362), .B(new_n216), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n516), .B(new_n517), .C1(new_n511), .C2(new_n515), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n512), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n362), .B(KEYINPUT19), .Z(new_n520));
  OAI21_X1  g334(.A(new_n377), .B1(new_n520), .B2(G146), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n518), .B1(new_n508), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n514), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G475), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n189), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n519), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n514), .B1(new_n512), .B2(new_n518), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n189), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G475), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n525), .A2(KEYINPUT20), .A3(new_n526), .A4(new_n189), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n529), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G952), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(G953), .ZN(new_n537));
  NAND2_X1  g351(.A1(G234), .A2(G237), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT21), .B(G898), .Z(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(G902), .A3(G953), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n540), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n505), .A2(new_n535), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n546), .A2(KEYINPUT91), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(KEYINPUT91), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n360), .A2(new_n479), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(G101), .ZN(G3));
  NAND2_X1  g365(.A1(new_n345), .A2(new_n356), .ZN(new_n552));
  INV_X1    g366(.A(new_n346), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n345), .A2(new_n346), .A3(new_n356), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n545), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n500), .A2(new_n558), .A3(new_n501), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n498), .A2(KEYINPUT33), .A3(new_n499), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(G478), .A3(new_n189), .A4(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT92), .B(G478), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n502), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n535), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n556), .A2(new_n557), .A3(new_n310), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G472), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n451), .B2(new_n189), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n451), .A2(new_n444), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n309), .A2(new_n393), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT34), .B(G104), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G6));
  INV_X1    g391(.A(new_n310), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n554), .B2(new_n555), .ZN(new_n579));
  INV_X1    g393(.A(new_n535), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n580), .A2(new_n505), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n579), .A2(new_n557), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n574), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G107), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G9));
  INV_X1    g399(.A(new_n573), .ZN(new_n586));
  INV_X1    g400(.A(new_n383), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(KEYINPUT36), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n380), .B(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n391), .A2(G902), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n389), .A2(new_n391), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n360), .A2(new_n549), .A3(new_n586), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G110), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT93), .B(KEYINPUT37), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G12));
  NOR3_X1   g410(.A1(new_n443), .A2(new_n395), .A3(new_n445), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT73), .B1(new_n597), .B2(new_n454), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n446), .A2(new_n394), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n478), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n579), .A2(new_n600), .A3(new_n308), .A4(new_n592), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT94), .B(G900), .Z(new_n602));
  AOI21_X1  g416(.A(new_n540), .B1(new_n544), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n581), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n225), .ZN(G30));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n505), .A2(new_n535), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n603), .B(KEYINPUT39), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n308), .A2(new_n611), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n578), .B(new_n609), .C1(new_n612), .C2(KEYINPUT40), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n441), .A2(new_n431), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n401), .B1(new_n471), .B2(new_n472), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(G472), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(G472), .A2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT95), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n592), .B1(new_n456), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n556), .B(KEYINPUT38), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(KEYINPUT40), .B2(new_n612), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n608), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n556), .B(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n612), .A2(KEYINPUT40), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n628), .A2(KEYINPUT96), .A3(new_n620), .A4(new_n613), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n218), .ZN(G45));
  NAND3_X1  g445(.A1(new_n564), .A2(new_n535), .A3(new_n604), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT97), .B1(new_n601), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n591), .B1(new_n456), .B2(new_n478), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n635));
  INV_X1    g449(.A(new_n632), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n360), .A2(new_n634), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT98), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n216), .ZN(G48));
  INV_X1    g454(.A(new_n393), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n189), .B1(new_n284), .B2(new_n294), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n301), .A2(KEYINPUT99), .A3(new_n189), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(G469), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n190), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n303), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n600), .A2(new_n641), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n567), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT41), .B(G113), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G15));
  NAND3_X1  g466(.A1(new_n579), .A2(new_n557), .A3(new_n581), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n649), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT100), .B(G116), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G18));
  NAND3_X1  g470(.A1(new_n549), .A2(new_n600), .A3(new_n592), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n579), .A2(new_n648), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n325), .ZN(G21));
  AOI22_X1  g474(.A1(new_n437), .A2(new_n442), .B1(new_n474), .B2(new_n401), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n444), .A2(KEYINPUT101), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n444), .A2(KEYINPUT101), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NOR4_X1   g478(.A1(new_n393), .A2(new_n664), .A3(new_n570), .A4(new_n545), .ZN(new_n665));
  INV_X1    g479(.A(new_n609), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n579), .A3(new_n666), .A4(new_n648), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G122), .ZN(G24));
  NOR4_X1   g482(.A1(new_n664), .A2(new_n591), .A3(new_n632), .A4(new_n570), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n579), .A2(new_n669), .A3(new_n648), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G125), .ZN(G27));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n304), .B2(new_n305), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n300), .A2(new_n196), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n673), .A2(G469), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n303), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n673), .A2(new_n679), .A3(G469), .A4(new_n675), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n191), .A2(new_n189), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT104), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  AOI22_X1  g498(.A1(KEYINPUT103), .A2(new_n676), .B1(new_n297), .B2(new_n302), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n680), .A2(new_n682), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n190), .A2(new_n578), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n554), .A2(new_n555), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n689), .A2(new_n479), .A3(new_n636), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT106), .B1(new_n597), .B2(new_n454), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n446), .A2(new_n452), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n478), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n698), .A2(KEYINPUT42), .A3(new_n641), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n699), .A2(new_n636), .A3(new_n689), .A4(new_n691), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G131), .ZN(G33));
  INV_X1    g516(.A(new_n605), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n689), .A2(new_n479), .A3(new_n703), .A4(new_n691), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G134), .ZN(G36));
  NOR2_X1   g519(.A1(new_n556), .A2(new_n578), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n580), .A2(new_n564), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n591), .B1(new_n709), .B2(KEYINPUT108), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n710), .B(new_n573), .C1(KEYINPUT108), .C2(new_n709), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n706), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT109), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n715), .B(new_n706), .C1(new_n711), .C2(new_n712), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n711), .A2(new_n712), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n675), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n720), .B1(new_n304), .B2(new_n305), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(G469), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n682), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(KEYINPUT46), .A3(new_n682), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n303), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n727), .A2(new_n647), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT107), .B1(new_n728), .B2(new_n611), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n611), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n717), .B(new_n718), .C1(new_n729), .C2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G137), .ZN(G39));
  XNOR2_X1  g548(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n727), .A2(new_n647), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(KEYINPUT47), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n728), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n706), .A2(new_n604), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n740), .A2(new_n565), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n456), .A3(new_n478), .A4(new_n393), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G140), .ZN(G42));
  INV_X1    g558(.A(new_n688), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n687), .B1(new_n685), .B2(new_n686), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n691), .B(new_n669), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n689), .A2(KEYINPUT114), .A3(new_n669), .A4(new_n691), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n741), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n505), .A2(new_n535), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n308), .A4(new_n634), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n701), .A2(new_n704), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n567), .A2(KEYINPUT113), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n579), .A2(new_n757), .A3(new_n557), .A4(new_n566), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n574), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n550), .A3(new_n583), .A4(new_n593), .ZN(new_n760));
  INV_X1    g574(.A(new_n658), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n549), .A2(new_n600), .A3(new_n592), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n600), .A2(new_n641), .A3(new_n648), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n761), .A2(new_n762), .B1(new_n582), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n303), .A2(new_n646), .A3(new_n647), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n359), .A2(new_n609), .A3(new_n766), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n568), .A2(new_n763), .B1(new_n767), .B2(new_n665), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n764), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  OAI22_X1  g583(.A1(new_n657), .A2(new_n658), .B1(new_n653), .B2(new_n649), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n667), .B1(new_n567), .B2(new_n649), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT112), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n760), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n670), .B1(new_n601), .B2(new_n605), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n609), .A2(new_n578), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n556), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n688), .B2(new_n684), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n647), .A3(new_n604), .A4(new_n620), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n638), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT52), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n774), .B1(new_n637), .B2(new_n633), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n779), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n755), .A2(new_n773), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n783), .B1(new_n782), .B2(new_n779), .ZN(new_n788));
  AND4_X1   g602(.A1(new_n783), .A2(new_n638), .A3(new_n775), .A4(new_n779), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(KEYINPUT53), .A3(new_n773), .A4(new_n755), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT54), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n760), .A2(new_n786), .A3(new_n771), .A4(new_n770), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n790), .A2(new_n755), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n787), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n540), .A2(new_n706), .A3(new_n648), .A4(new_n709), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n698), .A2(new_n641), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT48), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n456), .A2(new_n641), .A3(new_n619), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n540), .A3(new_n648), .A4(new_n706), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n801), .B(new_n537), .C1(new_n565), .C2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n706), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n303), .A2(new_n646), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n190), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n740), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n664), .A2(new_n570), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n641), .A2(new_n709), .A3(new_n540), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n626), .A2(new_n811), .A3(new_n578), .A4(new_n648), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT50), .Z(new_n814));
  NAND3_X1  g628(.A1(new_n798), .A2(new_n592), .A3(new_n810), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n803), .A2(new_n535), .A3(new_n564), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n812), .A2(new_n814), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT51), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n816), .B1(new_n809), .B2(new_n811), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n814), .A4(new_n815), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n804), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n811), .A2(new_n761), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n793), .A2(new_n797), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n536), .A2(new_n314), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n807), .B(KEYINPUT49), .Z(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n707), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n626), .A3(new_n690), .A4(new_n802), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(KEYINPUT115), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(G75));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n787), .A2(new_n796), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(G902), .ZN(new_n838));
  INV_X1    g652(.A(G210), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n317), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT55), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n840), .A2(new_n844), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n314), .A2(G952), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G51));
  XNOR2_X1  g662(.A(new_n681), .B(KEYINPUT57), .ZN(new_n849));
  INV_X1    g663(.A(new_n797), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n794), .B1(new_n787), .B2(new_n796), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT116), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n854), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n301), .B(KEYINPUT117), .Z(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n838), .A2(new_n722), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n847), .B1(new_n857), .B2(new_n858), .ZN(G54));
  NAND4_X1  g673(.A1(new_n837), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n860));
  INV_X1    g674(.A(new_n525), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n862), .A2(new_n863), .A3(new_n847), .ZN(G60));
  INV_X1    g678(.A(new_n847), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n559), .A2(new_n560), .ZN(new_n866));
  XNOR2_X1  g680(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n503), .A2(new_n189), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n866), .B(new_n869), .C1(new_n850), .C2(new_n851), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n793), .A2(new_n797), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n871), .A2(new_n869), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n865), .B(new_n870), .C1(new_n872), .C2(new_n866), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(G63));
  NAND2_X1  g688(.A1(G217), .A2(G902), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT119), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT60), .Z(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n787), .B2(new_n796), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n847), .B1(new_n878), .B2(new_n589), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n384), .B(KEYINPUT120), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n879), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(G66));
  NOR2_X1   g698(.A1(new_n773), .A2(G953), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n314), .B1(new_n541), .B2(G224), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT122), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n841), .B1(G898), .B2(new_n314), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n890), .B(new_n891), .Z(G69));
  NAND3_X1  g706(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT123), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n520), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n624), .A2(new_n629), .A3(new_n782), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n896), .A2(new_n897), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n743), .B(new_n898), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n612), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n581), .A2(new_n566), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n479), .A2(new_n905), .A3(new_n706), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n733), .A2(new_n314), .A3(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n314), .B1(new_n192), .B2(G900), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G900), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n895), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n733), .A2(new_n743), .A3(new_n701), .A4(new_n704), .ZN(new_n913));
  INV_X1    g727(.A(new_n777), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n799), .B(new_n914), .C1(new_n732), .C2(new_n729), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n782), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n910), .B1(new_n917), .B2(new_n314), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n912), .B1(new_n895), .B2(new_n918), .ZN(G72));
  XOR2_X1   g733(.A(new_n617), .B(KEYINPUT63), .Z(new_n920));
  NAND3_X1  g734(.A1(new_n733), .A2(new_n773), .A3(new_n907), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n904), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n457), .B(KEYINPUT125), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n400), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n920), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n461), .A2(new_n464), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n614), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n792), .A2(KEYINPUT126), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT126), .B1(new_n792), .B2(new_n928), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n925), .B(new_n865), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n917), .A2(new_n773), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n400), .B(new_n924), .C1(new_n933), .C2(new_n920), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT127), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n920), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(new_n458), .A3(new_n923), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n792), .A2(new_n928), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n847), .B1(new_n940), .B2(new_n929), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n937), .A2(new_n941), .A3(new_n942), .A4(new_n925), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n935), .A2(new_n943), .ZN(G57));
endmodule


