//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n463), .B(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n468), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n472), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  OR3_X1    g051(.A1(new_n468), .A2(KEYINPUT65), .A3(new_n474), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT65), .B1(new_n468), .B2(new_n474), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(new_n469), .B2(G136), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT66), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n489), .A2(G2104), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n472), .A2(G126), .A3(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n469), .A2(G138), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT67), .B1(new_n498), .B2(G651), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n503), .A2(G50), .A3(G543), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n507));
  XNOR2_X1  g082(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT69), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(KEYINPUT69), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n503), .A2(new_n513), .A3(new_n505), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n514), .A2(new_n501), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n508), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n503), .A2(G543), .A3(new_n505), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n504), .B1(new_n499), .B2(new_n502), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(KEYINPUT70), .A3(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n519), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n526), .A2(new_n529), .A3(new_n527), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n503), .A2(new_n513), .A3(G89), .A4(new_n505), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n525), .A2(new_n536), .ZN(G168));
  AND4_X1   g112(.A1(KEYINPUT70), .A2(new_n503), .A3(G543), .A4(new_n505), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT70), .B1(new_n523), .B2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(G52), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n513), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI211_X1 g118(.A(KEYINPUT72), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n543), .B1(new_n511), .B2(new_n512), .ZN(new_n546));
  INV_X1    g121(.A(new_n541), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(G651), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n523), .A2(G90), .A3(new_n513), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n540), .A2(new_n549), .A3(new_n550), .ZN(G171));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n522), .B2(new_n524), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n511), .B2(new_n512), .ZN(new_n555));
  AND2_X1   g130(.A1(G68), .A2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n523), .A2(G81), .A3(new_n513), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT74), .Z(G188));
  NAND4_X1  g142(.A1(new_n503), .A2(G53), .A3(G543), .A4(new_n505), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n523), .A2(new_n570), .A3(G53), .A4(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n511), .B2(new_n512), .ZN(new_n574));
  AND2_X1   g149(.A1(G78), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n503), .A2(new_n513), .A3(G91), .A4(new_n505), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n572), .A2(new_n578), .A3(KEYINPUT75), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT75), .B1(new_n572), .B2(new_n578), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(G299));
  NAND3_X1  g156(.A1(new_n540), .A2(new_n549), .A3(new_n550), .ZN(G301));
  INV_X1    g157(.A(G168), .ZN(G286));
  INV_X1    g158(.A(G166), .ZN(G303));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n511), .A2(new_n585), .A3(new_n512), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT76), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n523), .A2(G49), .A3(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n523), .A2(G87), .A3(new_n513), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(G288));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n511), .B2(new_n512), .ZN(new_n594));
  AND2_X1   g169(.A1(G73), .A2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n523), .A2(G86), .A3(new_n513), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n523), .A2(G48), .A3(G543), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G305));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n522), .B2(new_n524), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n602), .A2(new_n501), .B1(new_n515), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n515), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .A4(new_n513), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n542), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n610), .A2(new_n611), .B1(G651), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(G54), .B1(new_n538), .B2(new_n539), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n607), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n607), .B1(new_n618), .B2(G868), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n572), .A2(new_n578), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n572), .A2(new_n578), .A3(KEYINPUT75), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n621), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n621), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G860), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n617), .B1(G559), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT77), .ZN(G148));
  NOR2_X1   g206(.A1(new_n560), .A2(G868), .ZN(new_n632));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n618), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n632), .B1(new_n634), .B2(G868), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT78), .ZN(G323));
  XNOR2_X1  g211(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n637));
  XNOR2_X1  g212(.A(G323), .B(new_n637), .ZN(G282));
  NAND2_X1  g213(.A1(new_n479), .A2(G123), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n474), .A2(G111), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(KEYINPUT80), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n640), .B2(KEYINPUT80), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n641), .A2(new_n643), .B1(new_n469), .B2(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n472), .A2(new_n462), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT12), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT13), .Z(new_n649));
  INV_X1    g224(.A(G2100), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n645), .A2(G2096), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n651), .B(new_n652), .C1(new_n650), .C2(new_n649), .ZN(G156));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2443), .B(G2446), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2451), .B(G2454), .Z(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n666), .A2(KEYINPUT82), .A3(new_n654), .ZN(new_n667));
  AOI21_X1  g242(.A(KEYINPUT82), .B1(new_n666), .B2(new_n654), .ZN(new_n668));
  OAI221_X1 g243(.A(G14), .B1(new_n654), .B2(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(new_n650), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(G2096), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  AND2_X1   g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT84), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n691), .A2(new_n687), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(new_n684), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n690), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT85), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  NOR2_X1   g282(.A1(G95), .A2(G2105), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT86), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n709), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT87), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n469), .A2(G131), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n479), .A2(G119), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G25), .B2(new_n719), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n605), .B2(new_n725), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1986), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n723), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(G23), .ZN(new_n730));
  INV_X1    g305(.A(G288), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n725), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT33), .B(G1976), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n725), .A2(G22), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G166), .B2(new_n725), .ZN(new_n736));
  INV_X1    g311(.A(G1971), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G6), .A2(G16), .ZN(new_n739));
  INV_X1    g314(.A(G305), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G16), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT32), .B(G1981), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n734), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT34), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(KEYINPUT34), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n729), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT36), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n725), .A2(G20), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT23), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n626), .B2(new_n725), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G1956), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n719), .A2(G35), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G162), .B2(new_n719), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT29), .Z(new_n755));
  INV_X1    g330(.A(G2090), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(KEYINPUT97), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n755), .A2(new_n756), .ZN(new_n760));
  NOR2_X1   g335(.A1(G4), .A2(G16), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT89), .Z(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n617), .B2(new_n725), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1348), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n725), .A2(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n560), .B2(new_n725), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G1341), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n719), .A2(G26), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT28), .Z(new_n769));
  NAND3_X1  g344(.A1(new_n477), .A2(G128), .A3(new_n478), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  INV_X1    g346(.A(G116), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n469), .B2(G140), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n769), .B1(new_n775), .B2(G29), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2067), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n760), .A2(new_n764), .A3(new_n767), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n758), .B2(KEYINPUT97), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n472), .A2(G127), .ZN(new_n780));
  AND2_X1   g355(.A1(G115), .A2(G2104), .ZN(new_n781));
  OAI21_X1  g356(.A(G2105), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n783));
  NAND2_X1  g358(.A1(G103), .A2(G2104), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G2105), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n474), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n469), .A2(G139), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT90), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n719), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n719), .B2(G33), .ZN(new_n792));
  INV_X1    g367(.A(G2072), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT91), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n725), .A2(G5), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G171), .B2(new_n725), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n795), .B1(G1961), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G34), .ZN(new_n799));
  AOI21_X1  g374(.A(G29), .B1(new_n799), .B2(KEYINPUT24), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(KEYINPUT24), .B2(new_n799), .ZN(new_n801));
  INV_X1    g376(.A(G160), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n719), .ZN(new_n803));
  INV_X1    g378(.A(G2084), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT94), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT93), .ZN(new_n808));
  NAND3_X1  g383(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT92), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT26), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n469), .A2(G141), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n462), .A2(G105), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n477), .A2(G129), .A3(new_n478), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n719), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n719), .B2(G32), .ZN(new_n820));
  OAI221_X1 g395(.A(new_n806), .B1(G1961), .B2(new_n797), .C1(new_n808), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT95), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(KEYINPUT95), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT30), .B(G28), .ZN(new_n824));
  OR2_X1    g399(.A1(KEYINPUT31), .A2(G11), .ZN(new_n825));
  NAND2_X1  g400(.A1(KEYINPUT31), .A2(G11), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n824), .A2(new_n719), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n827), .B1(new_n719), .B2(new_n645), .C1(new_n803), .C2(new_n804), .ZN(new_n828));
  INV_X1    g403(.A(G2078), .ZN(new_n829));
  NAND2_X1  g404(.A1(G164), .A2(G29), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G27), .B2(G29), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n828), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n829), .B2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n820), .A2(new_n808), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n792), .B2(new_n793), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n725), .A2(G21), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G168), .B2(new_n725), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1966), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n833), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n798), .A2(new_n822), .A3(new_n823), .A4(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT96), .ZN(new_n841));
  AND4_X1   g416(.A1(new_n748), .A2(new_n759), .A3(new_n779), .A4(new_n841), .ZN(G311));
  NAND4_X1  g417(.A1(new_n748), .A2(new_n759), .A3(new_n779), .A4(new_n841), .ZN(G150));
  NOR2_X1   g418(.A1(new_n617), .A2(new_n633), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G55), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n522), .B2(new_n524), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n511), .B2(new_n512), .ZN(new_n850));
  AND2_X1   g425(.A1(G80), .A2(G543), .ZN(new_n851));
  OAI21_X1  g426(.A(G651), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n523), .A2(G93), .A3(new_n513), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n553), .A2(new_n559), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(G43), .B1(new_n538), .B2(new_n539), .ZN(new_n856));
  OAI21_X1  g431(.A(G55), .B1(new_n538), .B2(new_n539), .ZN(new_n857));
  INV_X1    g432(.A(new_n559), .ZN(new_n858));
  INV_X1    g433(.A(new_n854), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n846), .B(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n629), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n848), .A2(new_n854), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(new_n629), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(G145));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n871));
  AND4_X1   g446(.A1(new_n812), .A2(new_n814), .A3(new_n813), .A4(new_n815), .ZN(new_n872));
  INV_X1    g447(.A(new_n817), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n873), .A3(new_n775), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n770), .B(new_n774), .C1(new_n816), .C2(new_n817), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n875), .A3(G164), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(G164), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n871), .B(new_n790), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(new_n875), .ZN(new_n880));
  INV_X1    g455(.A(G164), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n788), .A3(new_n876), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n876), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n871), .B1(new_n885), .B2(new_n790), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n479), .A2(G130), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  INV_X1    g464(.A(G118), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(G2105), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n469), .B2(G142), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n648), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n711), .A2(new_n712), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(new_n714), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n713), .A2(new_n648), .A3(new_n715), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n894), .A3(new_n714), .ZN(new_n899));
  INV_X1    g474(.A(new_n893), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n648), .B1(new_n713), .B2(new_n715), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n887), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n898), .A2(new_n902), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n884), .B2(new_n886), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n485), .B(new_n645), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(G160), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(G160), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n898), .A2(KEYINPUT100), .A3(new_n902), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT101), .B1(new_n910), .B2(new_n911), .ZN(new_n915));
  INV_X1    g490(.A(new_n911), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n909), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n887), .A2(new_n914), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n905), .B(KEYINPUT100), .C1(new_n886), .C2(new_n884), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT102), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n886), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n922), .A2(new_n914), .A3(new_n883), .A4(new_n879), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n915), .A2(new_n918), .ZN(new_n924));
  AND4_X1   g499(.A1(KEYINPUT102), .A2(new_n920), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n913), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g502(.A(new_n740), .B1(new_n601), .B2(new_n604), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n605), .A2(G305), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n506), .B(KEYINPUT68), .ZN(new_n930));
  INV_X1    g505(.A(new_n517), .ZN(new_n931));
  NAND3_X1  g506(.A1(G288), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n591), .B(new_n588), .C1(new_n508), .C2(new_n517), .ZN(new_n933));
  AND4_X1   g508(.A1(new_n928), .A2(new_n929), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n933), .A2(new_n932), .B1(new_n929), .B2(new_n928), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT42), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(KEYINPUT104), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(KEYINPUT104), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n634), .B(new_n861), .ZN(new_n941));
  NAND2_X1  g516(.A1(G299), .A2(new_n618), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n617), .B1(new_n579), .B2(new_n580), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(KEYINPUT103), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n617), .B(new_n947), .C1(new_n579), .C2(new_n580), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n942), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT41), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(G299), .B2(new_n618), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n949), .A2(new_n950), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n945), .B1(new_n952), .B2(new_n941), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n938), .B1(new_n940), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n940), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G868), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(G868), .B2(new_n867), .ZN(G331));
  XNOR2_X1  g532(.A(G331), .B(KEYINPUT105), .ZN(G295));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n525), .A2(new_n959), .A3(new_n536), .ZN(new_n960));
  OAI21_X1  g535(.A(G51), .B1(new_n538), .B2(new_n539), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT106), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(G171), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n959), .B1(new_n525), .B2(new_n536), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(KEYINPUT106), .A3(new_n962), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(G301), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n862), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n965), .A2(G301), .A3(new_n966), .ZN(new_n969));
  AOI21_X1  g544(.A(G301), .B1(new_n965), .B2(new_n966), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n861), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n949), .A2(new_n950), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n951), .A2(new_n943), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n969), .A2(new_n970), .A3(new_n861), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n964), .A2(new_n967), .B1(new_n855), .B2(new_n860), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n944), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n936), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT107), .B1(new_n975), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n936), .B1(new_n972), .B2(new_n944), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n982), .B(new_n983), .C1(new_n952), .C2(new_n972), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n978), .B1(new_n952), .B2(new_n972), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n986), .B2(new_n936), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n944), .A2(new_n950), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n951), .A2(new_n946), .A3(new_n948), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n978), .B(new_n991), .C1(new_n992), .C2(new_n972), .ZN(new_n993));
  AOI21_X1  g568(.A(G37), .B1(new_n993), .B2(new_n936), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n988), .B1(new_n985), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n996));
  NOR4_X1   g571(.A1(new_n990), .A2(new_n995), .A3(KEYINPUT109), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n985), .A2(new_n994), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n999), .B2(KEYINPUT43), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n1000), .B2(new_n989), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n985), .A2(new_n988), .A3(new_n994), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n988), .B1(new_n985), .B2(new_n987), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT108), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1004), .A2(KEYINPUT108), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT44), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT110), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n996), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(KEYINPUT44), .A3(new_n989), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT109), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1000), .A2(new_n998), .A3(new_n989), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1008), .A2(new_n1017), .ZN(G397));
  OR2_X1    g593(.A1(G164), .A2(G1384), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT112), .B(G40), .Z(new_n1022));
  NAND2_X1  g597(.A1(G160), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n716), .B(new_n722), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n818), .B(G1996), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n775), .B(G2067), .Z(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1986), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n605), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1031), .B(KEYINPUT113), .Z(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n1030), .B2(new_n605), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1024), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G164), .A2(G1384), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1023), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1037), .A2(KEYINPUT114), .A3(new_n1038), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n804), .B(new_n1039), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1023), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n1037), .B2(KEYINPUT45), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1036), .B1(new_n1043), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G168), .A2(new_n1036), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(KEYINPUT51), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  OR3_X1    g627(.A1(new_n1049), .A2(KEYINPUT125), .A3(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(new_n1050), .B(KEYINPUT124), .Z(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT125), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1043), .A2(new_n1048), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n1058), .A2(new_n1036), .A3(G168), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G303), .A2(G8), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT55), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT45), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1021), .B(new_n1046), .C1(new_n1063), .C2(new_n1019), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1019), .A2(KEYINPUT50), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1065), .A2(new_n1039), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n737), .A2(new_n1064), .B1(new_n1066), .B2(new_n756), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1067), .B2(new_n1036), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n737), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n756), .B(new_n1039), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1062), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(G8), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1046), .A2(new_n1037), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G8), .ZN(new_n1076));
  XNOR2_X1  g651(.A(G305), .B(G1981), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1036), .B1(new_n1046), .B2(new_n1037), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n731), .A2(G1976), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1081), .B1(KEYINPUT52), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1976), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1082), .A2(new_n1083), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1082), .A2(KEYINPUT115), .A3(new_n1083), .A4(new_n1087), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1085), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1085), .A2(KEYINPUT117), .A3(new_n1092), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1074), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1961), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1064), .B2(G2078), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1105), .A2(KEYINPUT126), .ZN(new_n1106));
  OR4_X1    g681(.A1(new_n1104), .A2(new_n1045), .A3(new_n1047), .A4(G2078), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(KEYINPUT126), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(G301), .B(KEYINPUT54), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1021), .B1(new_n1063), .B2(new_n1019), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  AND4_X1   g688(.A1(KEYINPUT53), .A2(G160), .A3(G40), .A4(new_n829), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1103), .A2(new_n1106), .A3(new_n1108), .A4(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1060), .A2(new_n1097), .A3(new_n1111), .A4(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1075), .A2(G2067), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(G1348), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT60), .B(new_n1119), .C1(new_n1120), .C2(G1348), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n618), .A3(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1064), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1066), .A2(G1956), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n622), .A2(KEYINPUT57), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n578), .B(KEYINPUT119), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1132), .A2(KEYINPUT57), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n572), .B(KEYINPUT118), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1135), .A2(KEYINPUT120), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(KEYINPUT120), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1130), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1136), .B(new_n1137), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT61), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT122), .B(G1996), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1075), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT58), .B(G1341), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1064), .A2(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AND4_X1   g721(.A1(new_n1142), .A2(new_n1146), .A3(KEYINPUT59), .A4(new_n560), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1146), .A2(new_n560), .B1(new_n1142), .B2(KEYINPUT59), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1141), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1124), .A2(new_n618), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1139), .A2(KEYINPUT61), .A3(new_n1140), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1125), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1140), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n617), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1121), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1117), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1158));
  NOR4_X1   g733(.A1(new_n1058), .A2(KEYINPUT63), .A3(new_n1036), .A4(G286), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1085), .A2(G168), .A3(new_n1049), .A4(new_n1092), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1072), .B1(new_n1071), .B2(G8), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT63), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1093), .A2(new_n1073), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n731), .A2(new_n1086), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1081), .A2(new_n1165), .B1(G1981), .B2(G305), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT116), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1076), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1164), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1160), .A2(new_n1163), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1057), .A2(new_n1172), .A3(new_n1059), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1173), .A2(G171), .A3(new_n1109), .A4(new_n1097), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1172), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1171), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1035), .B1(new_n1156), .B2(new_n1176), .ZN(new_n1177));
  OR3_X1    g752(.A1(new_n1021), .A2(G1996), .A3(new_n1023), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1178), .A2(KEYINPUT46), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(KEYINPUT46), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1027), .A2(new_n818), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1179), .A2(new_n1180), .B1(new_n1024), .B2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT47), .Z(new_n1183));
  NAND2_X1  g758(.A1(new_n1029), .A2(new_n1024), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1032), .A2(new_n1024), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1185), .A2(KEYINPUT48), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(KEYINPUT48), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n718), .A2(new_n722), .ZN(new_n1189));
  OAI22_X1  g764(.A1(new_n1189), .A2(new_n1028), .B1(G2067), .B2(new_n775), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1024), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1183), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1177), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g769(.A1(G227), .A2(new_n459), .ZN(new_n1196));
  AND4_X1   g770(.A1(new_n669), .A2(new_n926), .A3(new_n706), .A4(new_n1196), .ZN(new_n1197));
  AND3_X1   g771(.A1(new_n1197), .A2(KEYINPUT127), .A3(new_n1009), .ZN(new_n1198));
  AOI21_X1  g772(.A(KEYINPUT127), .B1(new_n1197), .B2(new_n1009), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n1199), .ZN(G308));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1009), .ZN(G225));
endmodule


