

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(n524), .A2(G2105), .ZN(n877) );
  NOR2_X2 U554 ( .A1(n538), .A2(n537), .ZN(G160) );
  INV_X1 U555 ( .A(n614), .ZN(n657) );
  NAND2_X1 U556 ( .A1(G8), .A2(n614), .ZN(n702) );
  NOR2_X2 U557 ( .A1(n591), .A2(n540), .ZN(n784) );
  OR2_X1 U558 ( .A1(n696), .A2(n702), .ZN(n520) );
  AND2_X1 U559 ( .A1(n747), .A2(n740), .ZN(n521) );
  INV_X1 U560 ( .A(KEYINPUT26), .ZN(n615) );
  XNOR2_X1 U561 ( .A(n616), .B(n615), .ZN(n618) );
  INV_X1 U562 ( .A(KEYINPUT97), .ZN(n638) );
  XNOR2_X1 U563 ( .A(n638), .B(KEYINPUT27), .ZN(n639) );
  XNOR2_X1 U564 ( .A(n640), .B(n639), .ZN(n642) );
  INV_X1 U565 ( .A(KEYINPUT30), .ZN(n661) );
  XNOR2_X1 U566 ( .A(n661), .B(KEYINPUT101), .ZN(n662) );
  XNOR2_X1 U567 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X1 U568 ( .A1(n670), .A2(n669), .ZN(n681) );
  INV_X1 U569 ( .A(KEYINPUT102), .ZN(n686) );
  XNOR2_X1 U570 ( .A(n687), .B(n686), .ZN(n688) );
  AND2_X1 U571 ( .A1(G160), .A2(G40), .ZN(n601) );
  NAND2_X1 U572 ( .A1(n520), .A2(n1004), .ZN(n697) );
  OR2_X1 U573 ( .A1(n698), .A2(n697), .ZN(n705) );
  NOR2_X1 U574 ( .A1(G164), .A2(G1384), .ZN(n709) );
  INV_X1 U575 ( .A(G2104), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n521), .A2(n736), .ZN(n737) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n527), .ZN(n874) );
  XNOR2_X1 U578 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n523) );
  NOR2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X2 U580 ( .A(n523), .B(n522), .ZN(n879) );
  NAND2_X1 U581 ( .A1(G138), .A2(n879), .ZN(n526) );
  NAND2_X1 U582 ( .A1(G102), .A2(n877), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n526), .A2(n525), .ZN(n531) );
  INV_X1 U584 ( .A(G2105), .ZN(n527) );
  NOR2_X1 U585 ( .A1(n524), .A2(n527), .ZN(n873) );
  NAND2_X1 U586 ( .A1(G114), .A2(n873), .ZN(n529) );
  NAND2_X1 U587 ( .A1(G126), .A2(n874), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n531), .A2(n530), .ZN(G164) );
  NAND2_X1 U590 ( .A1(n879), .A2(G137), .ZN(n534) );
  NAND2_X1 U591 ( .A1(G101), .A2(n877), .ZN(n532) );
  XOR2_X1 U592 ( .A(n532), .B(KEYINPUT23), .Z(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U594 ( .A1(G113), .A2(n873), .ZN(n536) );
  NAND2_X1 U595 ( .A1(G125), .A2(n874), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U597 ( .A(KEYINPUT0), .B(G543), .Z(n591) );
  INV_X1 U598 ( .A(G651), .ZN(n540) );
  NAND2_X1 U599 ( .A1(G73), .A2(n784), .ZN(n539) );
  XNOR2_X1 U600 ( .A(n539), .B(KEYINPUT2), .ZN(n549) );
  NOR2_X1 U601 ( .A1(G543), .A2(n540), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n541), .Z(n780) );
  NAND2_X1 U603 ( .A1(n780), .A2(G61), .ZN(n544) );
  NOR2_X1 U604 ( .A1(G543), .A2(G651), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n542), .B(KEYINPUT64), .ZN(n781) );
  NAND2_X1 U606 ( .A1(G86), .A2(n781), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n547) );
  NOR2_X2 U608 ( .A1(G651), .A2(n591), .ZN(n785) );
  NAND2_X1 U609 ( .A1(G48), .A2(n785), .ZN(n545) );
  XNOR2_X1 U610 ( .A(KEYINPUT85), .B(n545), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n549), .A2(n548), .ZN(G305) );
  XNOR2_X1 U613 ( .A(KEYINPUT6), .B(KEYINPUT78), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G63), .A2(n780), .ZN(n551) );
  NAND2_X1 U615 ( .A1(G51), .A2(n785), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n781), .A2(G89), .ZN(n554) );
  XOR2_X1 U619 ( .A(KEYINPUT4), .B(n554), .Z(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT77), .ZN(n557) );
  NAND2_X1 U621 ( .A1(G76), .A2(n784), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT5), .B(n558), .Z(n559) );
  NOR2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U625 ( .A(KEYINPUT79), .B(KEYINPUT7), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n562), .B(n561), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G65), .A2(n780), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT70), .ZN(n570) );
  NAND2_X1 U630 ( .A1(n784), .A2(G78), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G91), .A2(n781), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U633 ( .A1(G53), .A2(n785), .ZN(n566) );
  XNOR2_X1 U634 ( .A(KEYINPUT71), .B(n566), .ZN(n567) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(G299) );
  NAND2_X1 U637 ( .A1(G52), .A2(n785), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n780), .A2(G64), .ZN(n571) );
  XNOR2_X1 U639 ( .A(KEYINPUT67), .B(n571), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n784), .A2(G77), .ZN(n573) );
  NAND2_X1 U641 ( .A1(G90), .A2(n781), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U643 ( .A(KEYINPUT68), .B(n574), .Z(n575) );
  XNOR2_X1 U644 ( .A(KEYINPUT9), .B(n575), .ZN(n576) );
  NOR2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT69), .ZN(G171) );
  NAND2_X1 U648 ( .A1(n784), .A2(G75), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G88), .A2(n781), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n780), .A2(G62), .ZN(n583) );
  XNOR2_X1 U652 ( .A(n583), .B(KEYINPUT86), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G50), .A2(n785), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(G166) );
  INV_X1 U656 ( .A(G166), .ZN(G303) );
  NAND2_X1 U657 ( .A1(G49), .A2(n785), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G74), .A2(G651), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U660 ( .A1(n780), .A2(n590), .ZN(n593) );
  NAND2_X1 U661 ( .A1(n591), .A2(G87), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(G288) );
  NAND2_X1 U663 ( .A1(n784), .A2(G72), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G85), .A2(n781), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G47), .A2(n785), .ZN(n596) );
  XOR2_X1 U667 ( .A(KEYINPUT66), .B(n596), .Z(n597) );
  NOR2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n780), .A2(G60), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(G290) );
  NAND2_X1 U671 ( .A1(n601), .A2(n709), .ZN(n614) );
  NOR2_X1 U672 ( .A1(G1981), .A2(G305), .ZN(n602) );
  XOR2_X1 U673 ( .A(n602), .B(KEYINPUT24), .Z(n603) );
  NOR2_X1 U674 ( .A1(n702), .A2(n603), .ZN(n707) );
  INV_X1 U675 ( .A(KEYINPUT32), .ZN(n680) );
  NAND2_X1 U676 ( .A1(G56), .A2(n780), .ZN(n604) );
  XOR2_X1 U677 ( .A(KEYINPUT14), .B(n604), .Z(n611) );
  NAND2_X1 U678 ( .A1(n781), .A2(G81), .ZN(n605) );
  XNOR2_X1 U679 ( .A(n605), .B(KEYINPUT72), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT12), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G68), .A2(n784), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U683 ( .A(KEYINPUT13), .B(n609), .Z(n610) );
  NOR2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n785), .A2(G43), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n995) );
  AND2_X1 U687 ( .A1(n657), .A2(G1996), .ZN(n616) );
  INV_X1 U688 ( .A(n657), .ZN(n672) );
  NAND2_X1 U689 ( .A1(n672), .A2(G1341), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U691 ( .A1(n995), .A2(n619), .ZN(n633) );
  NAND2_X1 U692 ( .A1(G66), .A2(n780), .ZN(n628) );
  NAND2_X1 U693 ( .A1(G54), .A2(n785), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n620), .B(KEYINPUT76), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n781), .A2(G92), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n621), .B(KEYINPUT74), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G79), .A2(n784), .ZN(n624) );
  XNOR2_X1 U699 ( .A(KEYINPUT75), .B(n624), .ZN(n625) );
  NOR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X2 U702 ( .A(n629), .B(KEYINPUT15), .ZN(n999) );
  INV_X1 U703 ( .A(n999), .ZN(n759) );
  NOR2_X1 U704 ( .A1(n657), .A2(G1348), .ZN(n631) );
  NOR2_X1 U705 ( .A1(G2067), .A2(n672), .ZN(n630) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n759), .A2(n634), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n636) );
  OR2_X1 U709 ( .A1(n634), .A2(n759), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U711 ( .A(KEYINPUT99), .B(n637), .ZN(n644) );
  NAND2_X1 U712 ( .A1(G2072), .A2(n657), .ZN(n640) );
  AND2_X1 U713 ( .A1(n672), .A2(G1956), .ZN(n641) );
  NOR2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n645) );
  INV_X1 U715 ( .A(G299), .ZN(n998) );
  NAND2_X1 U716 ( .A1(n645), .A2(n998), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n649) );
  NOR2_X1 U718 ( .A1(n645), .A2(n998), .ZN(n647) );
  XOR2_X1 U719 ( .A(KEYINPUT28), .B(KEYINPUT98), .Z(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n650), .B(KEYINPUT29), .ZN(n656) );
  XOR2_X1 U723 ( .A(G1961), .B(KEYINPUT94), .Z(n951) );
  NAND2_X1 U724 ( .A1(n951), .A2(n672), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT95), .ZN(n653) );
  XOR2_X1 U726 ( .A(KEYINPUT25), .B(G2078), .Z(n915) );
  NOR2_X1 U727 ( .A1(n672), .A2(n915), .ZN(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U729 ( .A(KEYINPUT96), .B(n654), .Z(n665) );
  AND2_X1 U730 ( .A1(G171), .A2(n665), .ZN(n655) );
  NOR2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n670) );
  INV_X1 U732 ( .A(G2084), .ZN(n658) );
  AND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n683) );
  NOR2_X1 U734 ( .A1(G1966), .A2(n702), .ZN(n682) );
  NOR2_X1 U735 ( .A1(n683), .A2(n682), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n659), .B(KEYINPUT100), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n660), .A2(G8), .ZN(n663) );
  NOR2_X1 U738 ( .A1(G168), .A2(n664), .ZN(n667) );
  NOR2_X1 U739 ( .A1(G171), .A2(n665), .ZN(n666) );
  NOR2_X1 U740 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(KEYINPUT31), .ZN(n669) );
  INV_X1 U742 ( .A(n681), .ZN(n671) );
  NAND2_X1 U743 ( .A1(G286), .A2(n671), .ZN(n677) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n702), .ZN(n674) );
  NOR2_X1 U745 ( .A1(G2090), .A2(n672), .ZN(n673) );
  NOR2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U747 ( .A1(n675), .A2(G303), .ZN(n676) );
  NAND2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n678), .A2(G8), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U752 ( .A1(G8), .A2(n683), .ZN(n684) );
  NAND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n690), .B(KEYINPUT103), .ZN(n701) );
  NOR2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n691) );
  NOR2_X1 U758 ( .A1(n1012), .A2(n691), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n701), .A2(n692), .ZN(n693) );
  NAND2_X1 U760 ( .A1(G1976), .A2(G288), .ZN(n1015) );
  NAND2_X1 U761 ( .A1(n693), .A2(n1015), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n702), .A2(n694), .ZN(n695) );
  NOR2_X1 U763 ( .A1(KEYINPUT33), .A2(n695), .ZN(n698) );
  NAND2_X1 U764 ( .A1(n1012), .A2(KEYINPUT33), .ZN(n696) );
  XOR2_X1 U765 ( .A(G1981), .B(G305), .Z(n1004) );
  NOR2_X1 U766 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U767 ( .A1(G8), .A2(n699), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n738) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n708) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n751) );
  XNOR2_X1 U774 ( .A(KEYINPUT93), .B(KEYINPUT36), .ZN(n721) );
  NAND2_X1 U775 ( .A1(G116), .A2(n873), .ZN(n711) );
  NAND2_X1 U776 ( .A1(G128), .A2(n874), .ZN(n710) );
  NAND2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U778 ( .A(KEYINPUT35), .B(n712), .ZN(n719) );
  XNOR2_X1 U779 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n717) );
  NAND2_X1 U780 ( .A1(G140), .A2(n879), .ZN(n714) );
  NAND2_X1 U781 ( .A1(G104), .A2(n877), .ZN(n713) );
  NAND2_X1 U782 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U783 ( .A(n715), .B(KEYINPUT34), .ZN(n716) );
  XNOR2_X1 U784 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U786 ( .A(n721), .B(n720), .ZN(n887) );
  XNOR2_X1 U787 ( .A(G2067), .B(KEYINPUT37), .ZN(n749) );
  NOR2_X1 U788 ( .A1(n887), .A2(n749), .ZN(n979) );
  NAND2_X1 U789 ( .A1(n751), .A2(n979), .ZN(n747) );
  NAND2_X1 U790 ( .A1(G141), .A2(n879), .ZN(n723) );
  NAND2_X1 U791 ( .A1(G117), .A2(n873), .ZN(n722) );
  NAND2_X1 U792 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U793 ( .A1(n877), .A2(G105), .ZN(n724) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n724), .Z(n725) );
  NOR2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U796 ( .A1(n874), .A2(G129), .ZN(n727) );
  NAND2_X1 U797 ( .A1(n728), .A2(n727), .ZN(n861) );
  AND2_X1 U798 ( .A1(n861), .A2(G1996), .ZN(n975) );
  NAND2_X1 U799 ( .A1(G131), .A2(n879), .ZN(n730) );
  NAND2_X1 U800 ( .A1(G107), .A2(n873), .ZN(n729) );
  NAND2_X1 U801 ( .A1(n730), .A2(n729), .ZN(n734) );
  NAND2_X1 U802 ( .A1(G95), .A2(n877), .ZN(n732) );
  NAND2_X1 U803 ( .A1(G119), .A2(n874), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n733) );
  OR2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n864) );
  AND2_X1 U806 ( .A1(n864), .A2(G1991), .ZN(n969) );
  OR2_X1 U807 ( .A1(n975), .A2(n969), .ZN(n735) );
  NAND2_X1 U808 ( .A1(n751), .A2(n735), .ZN(n740) );
  XNOR2_X1 U809 ( .A(G1986), .B(G290), .ZN(n1001) );
  NAND2_X1 U810 ( .A1(n1001), .A2(n751), .ZN(n736) );
  OR2_X1 U811 ( .A1(n738), .A2(n737), .ZN(n754) );
  NOR2_X1 U812 ( .A1(n861), .A2(G1996), .ZN(n739) );
  XNOR2_X1 U813 ( .A(n739), .B(KEYINPUT104), .ZN(n965) );
  INV_X1 U814 ( .A(n740), .ZN(n743) );
  NOR2_X1 U815 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U816 ( .A1(G1991), .A2(n864), .ZN(n971) );
  NOR2_X1 U817 ( .A1(n741), .A2(n971), .ZN(n742) );
  NOR2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U819 ( .A(KEYINPUT105), .B(n744), .Z(n745) );
  NOR2_X1 U820 ( .A1(n965), .A2(n745), .ZN(n746) );
  XNOR2_X1 U821 ( .A(n746), .B(KEYINPUT39), .ZN(n748) );
  NAND2_X1 U822 ( .A1(n748), .A2(n747), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n887), .A2(n749), .ZN(n980) );
  NAND2_X1 U824 ( .A1(n750), .A2(n980), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U827 ( .A(n755), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U828 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U829 ( .A(G57), .ZN(G237) );
  INV_X1 U830 ( .A(G132), .ZN(G219) );
  INV_X1 U831 ( .A(G82), .ZN(G220) );
  NAND2_X1 U832 ( .A1(G7), .A2(G661), .ZN(n756) );
  XNOR2_X1 U833 ( .A(n756), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U834 ( .A(G223), .ZN(n818) );
  NAND2_X1 U835 ( .A1(n818), .A2(G567), .ZN(n757) );
  XOR2_X1 U836 ( .A(KEYINPUT11), .B(n757), .Z(G234) );
  INV_X1 U837 ( .A(G860), .ZN(n764) );
  OR2_X1 U838 ( .A1(n995), .A2(n764), .ZN(n758) );
  XOR2_X1 U839 ( .A(KEYINPUT73), .B(n758), .Z(G153) );
  INV_X1 U840 ( .A(G171), .ZN(G301) );
  NAND2_X1 U841 ( .A1(G868), .A2(G301), .ZN(n761) );
  INV_X1 U842 ( .A(G868), .ZN(n801) );
  NAND2_X1 U843 ( .A1(n759), .A2(n801), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n761), .A2(n760), .ZN(G284) );
  NOR2_X1 U845 ( .A1(G868), .A2(G299), .ZN(n763) );
  NOR2_X1 U846 ( .A1(G286), .A2(n801), .ZN(n762) );
  NOR2_X1 U847 ( .A1(n763), .A2(n762), .ZN(G297) );
  NAND2_X1 U848 ( .A1(n764), .A2(G559), .ZN(n765) );
  NAND2_X1 U849 ( .A1(n765), .A2(n999), .ZN(n766) );
  XNOR2_X1 U850 ( .A(n766), .B(KEYINPUT16), .ZN(n767) );
  XNOR2_X1 U851 ( .A(KEYINPUT80), .B(n767), .ZN(G148) );
  NOR2_X1 U852 ( .A1(G868), .A2(n995), .ZN(n770) );
  NAND2_X1 U853 ( .A1(G868), .A2(n999), .ZN(n768) );
  NOR2_X1 U854 ( .A1(G559), .A2(n768), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n770), .A2(n769), .ZN(G282) );
  NAND2_X1 U856 ( .A1(G123), .A2(n874), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT18), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n873), .A2(G111), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n777) );
  NAND2_X1 U860 ( .A1(G135), .A2(n879), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G99), .A2(n877), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n968) );
  XOR2_X1 U864 ( .A(G2096), .B(n968), .Z(n778) );
  NOR2_X1 U865 ( .A1(G2100), .A2(n778), .ZN(n779) );
  XNOR2_X1 U866 ( .A(KEYINPUT81), .B(n779), .ZN(G156) );
  XNOR2_X1 U867 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n792) );
  NAND2_X1 U868 ( .A1(n780), .A2(G67), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G93), .A2(n781), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n789) );
  NAND2_X1 U871 ( .A1(G80), .A2(n784), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G55), .A2(n785), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U875 ( .A(KEYINPUT83), .B(n790), .ZN(n825) );
  XOR2_X1 U876 ( .A(G288), .B(n825), .Z(n791) );
  XNOR2_X1 U877 ( .A(n792), .B(n791), .ZN(n795) );
  XNOR2_X1 U878 ( .A(n998), .B(n995), .ZN(n793) );
  XNOR2_X1 U879 ( .A(n793), .B(G305), .ZN(n794) );
  XNOR2_X1 U880 ( .A(n795), .B(n794), .ZN(n797) );
  XNOR2_X1 U881 ( .A(G290), .B(G166), .ZN(n796) );
  XNOR2_X1 U882 ( .A(n797), .B(n796), .ZN(n890) );
  NAND2_X1 U883 ( .A1(G559), .A2(n999), .ZN(n798) );
  XOR2_X1 U884 ( .A(KEYINPUT82), .B(n798), .Z(n822) );
  XNOR2_X1 U885 ( .A(n890), .B(n822), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n799), .A2(G868), .ZN(n800) );
  XNOR2_X1 U887 ( .A(n800), .B(KEYINPUT88), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n801), .A2(n825), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n803), .A2(n802), .ZN(G295) );
  XNOR2_X1 U890 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n806) );
  NAND2_X1 U891 ( .A1(G2078), .A2(G2084), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(KEYINPUT89), .ZN(n805) );
  XNOR2_X1 U893 ( .A(n806), .B(n805), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G2090), .A2(n807), .ZN(n808) );
  XNOR2_X1 U895 ( .A(KEYINPUT21), .B(n808), .ZN(n809) );
  NAND2_X1 U896 ( .A1(n809), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U897 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U898 ( .A1(G220), .A2(G219), .ZN(n810) );
  XOR2_X1 U899 ( .A(KEYINPUT22), .B(n810), .Z(n811) );
  NOR2_X1 U900 ( .A1(G218), .A2(n811), .ZN(n812) );
  NAND2_X1 U901 ( .A1(G96), .A2(n812), .ZN(n827) );
  NAND2_X1 U902 ( .A1(n827), .A2(G2106), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G69), .A2(G120), .ZN(n813) );
  NOR2_X1 U904 ( .A1(G237), .A2(n813), .ZN(n814) );
  NAND2_X1 U905 ( .A1(G108), .A2(n814), .ZN(n828) );
  NAND2_X1 U906 ( .A1(n828), .A2(G567), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n829) );
  NAND2_X1 U908 ( .A1(G661), .A2(G483), .ZN(n817) );
  NOR2_X1 U909 ( .A1(n829), .A2(n817), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n821), .A2(G36), .ZN(G176) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n818), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U913 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(G188) );
  XOR2_X1 U917 ( .A(n822), .B(n995), .Z(n823) );
  NOR2_X1 U918 ( .A1(G860), .A2(n823), .ZN(n824) );
  XOR2_X1 U919 ( .A(n825), .B(n824), .Z(n826) );
  XNOR2_X1 U920 ( .A(n826), .B(KEYINPUT84), .ZN(G145) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  INV_X1 U926 ( .A(n829), .ZN(G319) );
  XOR2_X1 U927 ( .A(G2100), .B(G2096), .Z(n831) );
  XNOR2_X1 U928 ( .A(KEYINPUT42), .B(G2678), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U930 ( .A(KEYINPUT43), .B(G2072), .Z(n833) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2090), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U933 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2084), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(G227) );
  XOR2_X1 U936 ( .A(G1976), .B(G1966), .Z(n839) );
  XNOR2_X1 U937 ( .A(G1971), .B(G1961), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(n840), .B(G2474), .Z(n842) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1956), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U942 ( .A(KEYINPUT41), .B(G1981), .Z(n844) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G124), .A2(n874), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U948 ( .A1(n873), .A2(G112), .ZN(n848) );
  NAND2_X1 U949 ( .A1(n849), .A2(n848), .ZN(n853) );
  NAND2_X1 U950 ( .A1(G136), .A2(n879), .ZN(n851) );
  NAND2_X1 U951 ( .A1(G100), .A2(n877), .ZN(n850) );
  NAND2_X1 U952 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U953 ( .A1(n853), .A2(n852), .ZN(G162) );
  NAND2_X1 U954 ( .A1(G139), .A2(n879), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G103), .A2(n877), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G115), .A2(n873), .ZN(n857) );
  NAND2_X1 U958 ( .A1(G127), .A2(n874), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(KEYINPUT47), .B(n858), .Z(n859) );
  NOR2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n983) );
  XOR2_X1 U962 ( .A(n983), .B(n968), .Z(n863) );
  XOR2_X1 U963 ( .A(G160), .B(n861), .Z(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U965 ( .A(G164), .B(n864), .Z(n865) );
  XNOR2_X1 U966 ( .A(n865), .B(G162), .ZN(n866) );
  XOR2_X1 U967 ( .A(n867), .B(n866), .Z(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT108), .B(KEYINPUT48), .Z(n869) );
  XNOR2_X1 U969 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U971 ( .A(KEYINPUT109), .B(n870), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n886) );
  NAND2_X1 U973 ( .A1(G118), .A2(n873), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G130), .A2(n874), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n884) );
  NAND2_X1 U976 ( .A1(n877), .A2(G106), .ZN(n878) );
  XOR2_X1 U977 ( .A(KEYINPUT107), .B(n878), .Z(n881) );
  NAND2_X1 U978 ( .A1(n879), .A2(G142), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(n882), .B(KEYINPUT45), .Z(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n886), .B(n885), .Z(n888) );
  XOR2_X1 U983 ( .A(n888), .B(n887), .Z(n889) );
  NOR2_X1 U984 ( .A1(G37), .A2(n889), .ZN(G395) );
  XOR2_X1 U985 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n892) );
  XNOR2_X1 U986 ( .A(n999), .B(n890), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n894) );
  XOR2_X1 U988 ( .A(G301), .B(G286), .Z(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2438), .B(KEYINPUT106), .Z(n897) );
  XNOR2_X1 U992 ( .A(G2443), .B(G2430), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(n898), .B(G2435), .Z(n900) );
  XNOR2_X1 U995 ( .A(G1348), .B(G1341), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U997 ( .A(G2451), .B(G2427), .Z(n902) );
  XNOR2_X1 U998 ( .A(G2454), .B(G2446), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n904), .B(n903), .Z(n905) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n905), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  INV_X1 U1010 ( .A(n911), .ZN(G401) );
  XOR2_X1 U1011 ( .A(G25), .B(G1991), .Z(n912) );
  NAND2_X1 U1012 ( .A1(n912), .A2(G28), .ZN(n921) );
  XNOR2_X1 U1013 ( .A(G2067), .B(G26), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(G33), .B(G2072), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(G1996), .B(G32), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G27), .B(n915), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1021 ( .A(KEYINPUT53), .B(n922), .Z(n925) );
  XOR2_X1 U1022 ( .A(KEYINPUT54), .B(G34), .Z(n923) );
  XNOR2_X1 U1023 ( .A(G2084), .B(n923), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(G35), .B(G2090), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(n928), .B(KEYINPUT55), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(G29), .B(KEYINPUT115), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(G11), .A2(n931), .ZN(n963) );
  XOR2_X1 U1031 ( .A(G1976), .B(G23), .Z(n934) );
  XNOR2_X1 U1032 ( .A(G1986), .B(KEYINPUT125), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(n932), .B(G24), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(G22), .B(G1971), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1037 ( .A(KEYINPUT58), .B(n937), .Z(n957) );
  XOR2_X1 U1038 ( .A(G1966), .B(G21), .Z(n950) );
  XNOR2_X1 U1039 ( .A(G1341), .B(G19), .ZN(n938) );
  XNOR2_X1 U1040 ( .A(n938), .B(KEYINPUT121), .ZN(n941) );
  XOR2_X1 U1041 ( .A(G1981), .B(G6), .Z(n939) );
  XNOR2_X1 U1042 ( .A(KEYINPUT122), .B(n939), .ZN(n940) );
  NAND2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(KEYINPUT123), .B(n942), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(G1348), .B(KEYINPUT59), .ZN(n943) );
  XNOR2_X1 U1046 ( .A(n943), .B(G4), .ZN(n944) );
  NAND2_X1 U1047 ( .A1(n945), .A2(n944), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(G20), .B(G1956), .ZN(n946) );
  NOR2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1050 ( .A(KEYINPUT60), .B(n948), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n954) );
  XOR2_X1 U1052 ( .A(G5), .B(n951), .Z(n952) );
  XNOR2_X1 U1053 ( .A(KEYINPUT120), .B(n952), .ZN(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1055 ( .A(KEYINPUT124), .B(n955), .Z(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1057 ( .A(n958), .B(KEYINPUT126), .Z(n959) );
  XNOR2_X1 U1058 ( .A(KEYINPUT61), .B(n959), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(G16), .A2(n960), .ZN(n961) );
  XOR2_X1 U1060 ( .A(KEYINPUT127), .B(n961), .Z(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n994) );
  XOR2_X1 U1062 ( .A(G2090), .B(G162), .Z(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(KEYINPUT51), .B(n966), .ZN(n967) );
  XNOR2_X1 U1065 ( .A(n967), .B(KEYINPUT113), .ZN(n977) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n973) );
  XOR2_X1 U1067 ( .A(G160), .B(G2084), .Z(n970) );
  NOR2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(KEYINPUT114), .B(n982), .ZN(n988) );
  XOR2_X1 U1075 ( .A(G2072), .B(n983), .Z(n985) );
  XOR2_X1 U1076 ( .A(G164), .B(G2078), .Z(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT50), .B(n986), .Z(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(KEYINPUT52), .B(n989), .ZN(n991) );
  INV_X1 U1081 ( .A(KEYINPUT55), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n992), .A2(G29), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n1024) );
  XOR2_X1 U1085 ( .A(KEYINPUT56), .B(G16), .Z(n1022) );
  XNOR2_X1 U1086 ( .A(G301), .B(G1961), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n995), .B(G1341), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1011) );
  XNOR2_X1 U1089 ( .A(n998), .B(G1956), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(G1348), .B(n999), .Z(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(G168), .B(G1966), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1006), .B(KEYINPUT116), .ZN(n1007) );
  XOR2_X1 U1096 ( .A(KEYINPUT57), .B(n1007), .Z(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1019) );
  XOR2_X1 U1099 ( .A(n1012), .B(KEYINPUT117), .Z(n1014) );
  XOR2_X1 U1100 ( .A(G166), .B(G1971), .Z(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(KEYINPUT118), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(KEYINPUT119), .B(n1020), .Z(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(n1025), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

