//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g0012(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT66), .B(G244), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G77), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G87), .A2(G250), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n209), .B1(new_n218), .B2(new_n220), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G68), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n242), .B(new_n248), .ZN(G351));
  XNOR2_X1  g0049(.A(G97), .B(G107), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT6), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G97), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n251), .A2(new_n253), .A3(G107), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n216), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT75), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT75), .ZN(new_n262));
  INV_X1    g0062(.A(new_n260), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n254), .B1(new_n251), .B2(new_n250), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n262), .B(new_n263), .C1(new_n264), .C2(new_n216), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT7), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G107), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n261), .A2(new_n265), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n212), .A2(new_n213), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G13), .A3(G20), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G97), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n282), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n284), .B1(new_n288), .B2(new_n253), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n212), .A2(new_n213), .B1(G33), .B2(G41), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT4), .A2(G244), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n270), .A2(new_n272), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n270), .A2(new_n272), .A3(G250), .A4(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G283), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT4), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT74), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n271), .B2(G33), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n269), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n272), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G244), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n300), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n292), .B1(new_n299), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT5), .B(G41), .ZN(new_n310));
  INV_X1    g0110(.A(G41), .ZN(new_n311));
  OAI211_X1 g0111(.A(G1), .B(G13), .C1(new_n269), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n281), .A2(G45), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n310), .A2(new_n312), .A3(G274), .A4(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n314), .B2(new_n310), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G257), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(G200), .B1(new_n309), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n302), .A2(new_n272), .A3(new_n303), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT4), .B1(new_n322), .B2(new_n306), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n291), .B1(new_n323), .B2(new_n298), .ZN(new_n324));
  INV_X1    g0124(.A(new_n315), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(G257), .B2(new_n317), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n326), .A3(G190), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n280), .A2(new_n290), .A3(new_n321), .A4(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(G169), .B1(new_n309), .B2(new_n320), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n324), .A2(new_n326), .A3(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n289), .B1(new_n277), .B2(new_n279), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n328), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT24), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT83), .ZN(new_n336));
  INV_X1    g0136(.A(G87), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(G20), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(new_n270), .A3(new_n272), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT22), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT82), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT82), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT22), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n346), .A2(new_n267), .A3(KEYINPUT83), .A4(new_n338), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n302), .A2(new_n303), .A3(new_n216), .A4(new_n272), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT22), .B1(new_n349), .B2(new_n337), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT23), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n216), .B2(G107), .ZN(new_n353));
  INV_X1    g0153(.A(G107), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(KEYINPUT23), .A3(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G116), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(G20), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n335), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  AOI211_X1 g0160(.A(KEYINPUT24), .B(new_n358), .C1(new_n348), .C2(new_n350), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n279), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n288), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT25), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n282), .B2(G107), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n285), .A2(KEYINPUT25), .A3(new_n354), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n363), .A2(G107), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n319), .A2(G1698), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(G250), .B2(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(G294), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n304), .A2(new_n369), .B1(new_n269), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n291), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n317), .A2(G264), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n315), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n371), .A2(new_n291), .B1(new_n317), .B2(G264), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n315), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n362), .A2(new_n367), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT84), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n362), .A2(KEYINPUT84), .A3(new_n367), .A4(new_n380), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n334), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n267), .A2(G223), .A3(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n267), .A2(new_n294), .ZN(new_n387));
  INV_X1    g0187(.A(G222), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n386), .B1(new_n259), .B2(new_n267), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n291), .ZN(new_n390));
  INV_X1    g0190(.A(G45), .ZN(new_n391));
  AOI21_X1  g0191(.A(G1), .B1(new_n311), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n312), .A2(G274), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n281), .B1(G41), .B2(G45), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n312), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT67), .B(G226), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n378), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(G200), .B2(new_n400), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n281), .A2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n286), .A2(G50), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT8), .B(G58), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n216), .A2(G33), .ZN(new_n406));
  INV_X1    g0206(.A(G150), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n405), .A2(new_n406), .B1(new_n407), .B2(new_n258), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(G20), .B2(new_n203), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n212), .A2(new_n213), .A3(new_n278), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n404), .B1(G50), .B2(new_n282), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT9), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n402), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT70), .ZN(new_n414));
  INV_X1    g0214(.A(new_n400), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n375), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(KEYINPUT10), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(KEYINPUT10), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n402), .A3(new_n412), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n411), .B1(new_n415), .B2(G169), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n400), .A2(G179), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G58), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n244), .ZN(new_n427));
  OAI21_X1  g0227(.A(G20), .B1(new_n427), .B2(new_n201), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n257), .A2(G159), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n303), .A2(new_n272), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT74), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n266), .B(new_n216), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G68), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n266), .B1(new_n304), .B2(new_n216), .ZN(new_n436));
  OAI211_X1 g0236(.A(KEYINPUT16), .B(new_n431), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT16), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n244), .B1(new_n268), .B2(new_n274), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(new_n430), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n279), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n426), .A2(KEYINPUT8), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT8), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G58), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n445), .A2(new_n403), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n286), .A2(new_n446), .B1(new_n285), .B2(new_n405), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G232), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n393), .B1(new_n396), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(G223), .A2(G1698), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G226), .B2(new_n294), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n304), .A2(new_n452), .B1(new_n269), .B2(new_n337), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(new_n291), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G179), .ZN(new_n455));
  INV_X1    g0255(.A(G169), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n454), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n448), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT18), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT18), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n448), .A2(new_n460), .A3(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n453), .A2(new_n291), .ZN(new_n462));
  INV_X1    g0262(.A(new_n450), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(new_n378), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(G200), .B2(new_n454), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(new_n441), .A3(new_n447), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT17), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n465), .A2(new_n441), .A3(KEYINPUT17), .A4(new_n447), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n459), .A2(new_n461), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT73), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G97), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n449), .A2(G1698), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(G226), .B2(G1698), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n474), .B2(new_n273), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n291), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n393), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT71), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n316), .A2(new_n392), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT71), .B1(new_n312), .B2(new_n395), .ZN(new_n480));
  INV_X1    g0280(.A(G238), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT13), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n394), .B1(new_n291), .B2(new_n475), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT13), .ZN(new_n485));
  INV_X1    g0285(.A(new_n480), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n312), .A2(KEYINPUT71), .A3(new_n395), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(G238), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n484), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n483), .A2(G190), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT72), .B1(new_n282), .B2(G68), .ZN(new_n491));
  XOR2_X1   g0291(.A(new_n491), .B(KEYINPUT12), .Z(new_n492));
  NAND2_X1  g0292(.A1(new_n244), .A2(G20), .ZN(new_n493));
  OAI221_X1 g0293(.A(new_n493), .B1(new_n406), .B2(new_n259), .C1(new_n258), .C2(new_n202), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n279), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT11), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(KEYINPUT11), .A3(new_n279), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n286), .A2(G68), .A3(new_n403), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n492), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n490), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n375), .B1(new_n483), .B2(new_n489), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n471), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n483), .A2(new_n489), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(KEYINPUT73), .A3(new_n490), .A4(new_n501), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT14), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n477), .A2(new_n482), .A3(KEYINPUT13), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n485), .B1(new_n484), .B2(new_n488), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(G169), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n483), .A2(G179), .A3(new_n489), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n509), .B1(new_n505), .B2(G169), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n500), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n273), .A2(G107), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n387), .B2(new_n449), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n273), .A2(new_n481), .A3(new_n294), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n291), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n394), .B1(new_n223), .B2(new_n397), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G200), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n405), .A2(new_n258), .B1(new_n216), .B2(new_n259), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT68), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT15), .B(G87), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n525), .A2(new_n526), .B1(new_n406), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n445), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(KEYINPUT68), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n279), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n403), .A2(G77), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n286), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n285), .A2(new_n259), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n521), .A2(G190), .A3(new_n522), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n524), .A2(new_n531), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n523), .A2(new_n456), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n531), .A2(new_n536), .ZN(new_n540));
  INV_X1    g0340(.A(G179), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n521), .A2(new_n541), .A3(new_n522), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n544), .B(KEYINPUT69), .ZN(new_n545));
  NOR4_X1   g0345(.A1(new_n425), .A2(new_n470), .A3(new_n517), .A4(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n374), .A2(G179), .ZN(new_n547));
  AOI21_X1  g0347(.A(G169), .B1(new_n377), .B2(new_n315), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n322), .A2(new_n216), .A3(G87), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(KEYINPUT22), .B1(new_n341), .B2(new_n347), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT24), .B1(new_n551), .B2(new_n358), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n351), .A2(new_n335), .A3(new_n359), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n410), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n367), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n303), .A2(new_n272), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n557), .A2(new_n216), .A3(G68), .A4(new_n302), .ZN(new_n558));
  NOR2_X1   g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n337), .B1(new_n472), .B2(new_n216), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G97), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n560), .A2(new_n561), .B1(new_n406), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n410), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n527), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n282), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT77), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n349), .A2(new_n244), .ZN(new_n568));
  AND4_X1   g0368(.A1(new_n561), .A2(new_n216), .A3(G33), .A4(G97), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n337), .A2(new_n253), .A3(new_n354), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n472), .A2(new_n216), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n572), .B2(KEYINPUT19), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n279), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT77), .ZN(new_n575));
  INV_X1    g0375(.A(new_n566), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n567), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n363), .A2(new_n565), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n305), .A2(G1698), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G238), .B2(G1698), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n357), .B1(new_n304), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n291), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n312), .A2(G250), .A3(new_n313), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n312), .A2(G274), .A3(new_n314), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n541), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n588), .B1(new_n291), .B2(new_n584), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(new_n456), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n581), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(G169), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(G179), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT76), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n580), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n585), .A2(new_n589), .A3(G190), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT78), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n599), .A2(new_n600), .B1(G200), .B2(new_n590), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n288), .A2(new_n337), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT78), .B1(new_n590), .B2(new_n378), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n601), .A2(new_n578), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n556), .A2(new_n598), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n310), .A2(new_n314), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(G270), .A3(new_n312), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n315), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n319), .A2(new_n294), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(G264), .B2(new_n294), .ZN(new_n611));
  INV_X1    g0411(.A(G303), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n304), .A2(new_n611), .B1(new_n612), .B2(new_n267), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n291), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT79), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT79), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n291), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n609), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n410), .A2(G116), .A3(new_n282), .A4(new_n287), .ZN(new_n619));
  INV_X1    g0419(.A(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n285), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(G20), .B1(G33), .B2(G283), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n269), .A2(G97), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n622), .A2(new_n623), .B1(G20), .B2(new_n620), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n624), .A2(new_n279), .A3(KEYINPUT20), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT20), .B1(new_n624), .B2(new_n279), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n619), .B(new_n621), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G169), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT80), .B1(new_n618), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n609), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n613), .A2(new_n616), .A3(new_n291), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n616), .B1(new_n613), .B2(new_n291), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT80), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(G169), .A4(new_n627), .ZN(new_n635));
  XNOR2_X1  g0435(.A(KEYINPUT81), .B(KEYINPUT21), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n629), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n608), .A2(G179), .A3(new_n315), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n627), .B(new_n638), .C1(new_n631), .C2(new_n632), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n618), .A2(new_n628), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(KEYINPUT21), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n627), .B1(new_n633), .B2(G200), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n378), .B2(new_n633), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n637), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n385), .A2(new_n546), .A3(new_n606), .A4(new_n645), .ZN(G372));
  INV_X1    g0446(.A(new_n508), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n516), .B1(new_n647), .B2(new_n543), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n468), .A3(new_n469), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n459), .A2(new_n461), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n423), .B1(new_n652), .B2(new_n420), .ZN(new_n653));
  INV_X1    g0453(.A(new_n546), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n578), .A2(new_n579), .B1(new_n595), .B2(new_n596), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n564), .A2(KEYINPUT77), .A3(new_n566), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n575), .B1(new_n574), .B2(new_n576), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n603), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT85), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT85), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n578), .A2(new_n660), .A3(new_n603), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n599), .B1(G200), .B2(new_n590), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n655), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT88), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT88), .B1(new_n329), .B2(new_n330), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n666), .A2(new_n667), .A3(new_n333), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n664), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n280), .A2(new_n290), .B1(new_n329), .B2(new_n330), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n598), .A2(new_n670), .A3(new_n605), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n655), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT86), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n385), .B2(new_n664), .ZN(new_n675));
  INV_X1    g0475(.A(new_n556), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n637), .A2(new_n642), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT87), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n637), .A2(new_n642), .A3(KEYINPUT87), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n385), .A2(new_n674), .A3(new_n664), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n673), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n653), .B1(new_n654), .B2(new_n684), .ZN(G369));
  NOR2_X1   g0485(.A1(new_n645), .A2(KEYINPUT89), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n281), .A2(new_n216), .A3(G13), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n627), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n645), .A2(KEYINPUT89), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n680), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT87), .B1(new_n637), .B2(new_n642), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n693), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(G330), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n692), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n676), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n552), .A2(new_n553), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n555), .B1(new_n703), .B2(new_n279), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n701), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n383), .B2(new_n384), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n702), .B1(new_n706), .B2(new_n676), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n706), .A2(new_n556), .A3(new_n677), .A4(new_n701), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n702), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n207), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n570), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n220), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(new_n334), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT84), .B1(new_n704), .B2(new_n380), .ZN(new_n722));
  INV_X1    g0522(.A(new_n384), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n660), .B1(new_n578), .B2(new_n603), .ZN(new_n725));
  AOI211_X1 g0525(.A(KEYINPUT85), .B(new_n602), .C1(new_n567), .C2(new_n577), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n663), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n655), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT86), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n556), .B1(new_n697), .B2(new_n698), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n683), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n673), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n692), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n383), .A2(new_n384), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n556), .A2(new_n637), .A3(new_n642), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n664), .A2(new_n737), .A3(new_n721), .A4(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n668), .A2(new_n727), .A3(new_n728), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT26), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n598), .A2(new_n605), .A3(new_n665), .A4(new_n670), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n728), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT91), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n746), .B1(new_n745), .B2(new_n747), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n734), .A2(new_n736), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G330), .ZN(new_n752));
  AND4_X1   g0552(.A1(new_n637), .A2(new_n642), .A3(new_n644), .A4(new_n701), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n385), .A2(new_n753), .A3(new_n606), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n592), .A2(new_n638), .A3(new_n377), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n309), .A2(new_n320), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n615), .A2(new_n617), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n755), .A2(KEYINPUT30), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT30), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n324), .B(new_n326), .C1(new_n631), .C2(new_n632), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n592), .A2(new_n638), .A3(new_n377), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n592), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n324), .A2(new_n326), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n633), .A2(new_n763), .A3(new_n374), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n758), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n766), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n767));
  AOI21_X1  g0567(.A(KEYINPUT31), .B1(new_n766), .B2(new_n692), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n752), .B1(new_n754), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n751), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n720), .B1(new_n771), .B2(G1), .ZN(G364));
  NAND2_X1  g0572(.A1(new_n696), .A2(new_n699), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n215), .B1(G20), .B2(new_n456), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n216), .A2(G179), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(new_n378), .A3(G200), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT96), .Z(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n354), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n378), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n216), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT95), .B(G159), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT32), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G97), .A2(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n793), .B(new_n267), .C1(new_n792), .C2(new_n791), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n780), .A2(G190), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n216), .A2(new_n541), .A3(new_n375), .A4(G190), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n796), .A2(G87), .B1(new_n797), .B2(G68), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n216), .A2(new_n541), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(G190), .A3(G200), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n202), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n784), .A2(new_n794), .A3(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n799), .B(KEYINPUT92), .Z(new_n803));
  INV_X1    g0603(.A(KEYINPUT94), .ZN(new_n804));
  AND3_X1   g0604(.A1(new_n803), .A2(new_n804), .A3(new_n788), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(new_n803), .B2(new_n788), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n803), .A2(G190), .A3(new_n375), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT93), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n802), .B1(new_n259), .B2(new_n807), .C1(new_n426), .C2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n800), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G294), .A2(new_n787), .B1(new_n814), .B2(G326), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT97), .ZN(new_n818));
  INV_X1    g0618(.A(new_n789), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n267), .B1(new_n819), .B2(G329), .ZN(new_n820));
  INV_X1    g0620(.A(G317), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(KEYINPUT33), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(KEYINPUT33), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n797), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G303), .B2(new_n796), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  INV_X1    g0627(.A(G322), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n826), .B1(new_n827), .B2(new_n783), .C1(new_n812), .C2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n813), .B1(new_n818), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n779), .B1(new_n830), .B2(KEYINPUT98), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(KEYINPUT98), .B2(new_n830), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n216), .A2(G13), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n281), .B1(new_n833), .B2(G45), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n715), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n714), .A2(new_n273), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(G355), .B1(new_n620), .B2(new_n714), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n248), .A2(new_n391), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n322), .A2(new_n714), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(G45), .B2(new_n220), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n839), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n778), .A2(new_n776), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n837), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n777), .A2(new_n832), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n773), .A2(new_n752), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n700), .A3(new_n837), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT99), .Z(G396));
  INV_X1    g0650(.A(KEYINPUT102), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n540), .A2(new_n692), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n538), .A2(new_n543), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT101), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n538), .A2(new_n543), .A3(KEYINPUT101), .A4(new_n852), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n543), .A2(new_n701), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n851), .B1(new_n734), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(KEYINPUT102), .B(new_n858), .C1(new_n684), .C2(new_n692), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n732), .A2(new_n733), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n692), .B1(new_n855), .B2(new_n856), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n860), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n770), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n836), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n858), .A2(new_n774), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n778), .A2(new_n774), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n812), .A2(new_n370), .B1(new_n620), .B2(new_n807), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n783), .A2(new_n337), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n273), .B1(new_n789), .B2(new_n816), .C1(new_n786), .C2(new_n253), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n796), .A2(G107), .B1(new_n797), .B2(G283), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n612), .B2(new_n800), .ZN(new_n876));
  NOR4_X1   g0676(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n783), .A2(new_n244), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n304), .B1(new_n819), .B2(G132), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n879), .B1(new_n202), .B2(new_n795), .C1(new_n426), .C2(new_n786), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n814), .A2(G137), .B1(new_n797), .B2(G150), .ZN(new_n881));
  INV_X1    g0681(.A(G143), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n881), .B1(new_n807), .B2(new_n790), .C1(new_n812), .C2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT34), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n878), .B(new_n880), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n877), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n836), .B1(G77), .B2(new_n871), .C1(new_n887), .C2(new_n779), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT100), .Z(new_n889));
  AOI22_X1  g0689(.A1(new_n867), .A2(new_n868), .B1(new_n869), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(G384));
  INV_X1    g0691(.A(new_n264), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n892), .A2(KEYINPUT35), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(KEYINPUT35), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n893), .A2(G116), .A3(new_n217), .A4(new_n894), .ZN(new_n895));
  XOR2_X1   g0695(.A(KEYINPUT103), .B(KEYINPUT36), .Z(new_n896));
  XNOR2_X1  g0696(.A(new_n895), .B(new_n896), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n220), .A2(new_n259), .A3(new_n427), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n281), .B(G13), .C1(new_n898), .C2(new_n243), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n501), .A2(new_n701), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n517), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n508), .B(new_n516), .C1(new_n501), .C2(new_n701), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n858), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n754), .A2(new_n769), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n690), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n448), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n470), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n458), .A2(new_n908), .A3(new_n466), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n458), .A2(new_n908), .A3(new_n913), .A4(new_n466), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT106), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n470), .A2(new_n909), .B1(new_n912), .B2(new_n914), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT106), .B1(new_n919), .B2(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n441), .A2(new_n447), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n437), .A2(new_n279), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n304), .A2(new_n216), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT7), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(G68), .A3(new_n434), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT16), .B1(new_n926), .B2(new_n431), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n447), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n922), .A2(new_n465), .B1(new_n928), .B2(new_n907), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n457), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n913), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n914), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT104), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n928), .A2(new_n907), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n930), .A2(new_n934), .A3(new_n466), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT37), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT104), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n937), .A3(new_n914), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT38), .ZN(new_n939));
  INV_X1    g0739(.A(new_n934), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n939), .B1(new_n470), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n933), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n906), .B1(new_n921), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n904), .A2(new_n905), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n944), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n942), .A2(KEYINPUT105), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT105), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n933), .A2(new_n938), .A3(new_n941), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n470), .A2(new_n940), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n933), .A2(new_n950), .A3(new_n938), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n947), .A2(new_n949), .B1(new_n939), .B2(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n943), .A2(new_n944), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n953), .A2(new_n546), .A3(new_n905), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n546), .B2(new_n905), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n954), .A2(new_n955), .A3(new_n752), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n651), .A2(new_n907), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n902), .A2(new_n903), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n543), .A2(new_n692), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n959), .B1(new_n864), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n952), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT39), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n916), .A2(new_n917), .ZN(new_n966));
  AOI211_X1 g0766(.A(KEYINPUT106), .B(KEYINPUT38), .C1(new_n910), .C2(new_n915), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n965), .B(new_n942), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n952), .B2(new_n965), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n516), .A2(new_n692), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n653), .B1(new_n750), .B2(new_n654), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n956), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n281), .B2(new_n833), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n956), .A2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n900), .B1(new_n977), .B2(new_n978), .ZN(G367));
  NAND2_X1  g0779(.A1(new_n796), .A2(G116), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT46), .Z(new_n981));
  OAI21_X1  g0781(.A(new_n304), .B1(new_n821), .B2(new_n789), .ZN(new_n982));
  INV_X1    g0782(.A(new_n797), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n983), .A2(new_n370), .B1(new_n781), .B2(new_n253), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n786), .A2(new_n354), .B1(new_n800), .B2(new_n816), .ZN(new_n985));
  NOR4_X1   g0785(.A1(new_n981), .A2(new_n982), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n827), .B2(new_n807), .C1(new_n612), .C2(new_n812), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n273), .B1(new_n819), .B2(G137), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n882), .B2(new_n800), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n426), .A2(new_n795), .B1(new_n781), .B2(new_n259), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n983), .A2(new_n790), .B1(new_n244), .B2(new_n786), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n202), .B2(new_n807), .C1(new_n812), .C2(new_n407), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT47), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n778), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n776), .B(new_n778), .C1(new_n714), .C2(new_n565), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n238), .A2(new_n841), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n837), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n659), .A2(new_n661), .A3(new_n692), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n664), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n728), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n776), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n996), .B(new_n999), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n710), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT108), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n692), .B1(new_n637), .B2(new_n642), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1008), .B1(new_n707), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n700), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n700), .A2(new_n1011), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1007), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1014), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1016), .A2(new_n1012), .A3(new_n710), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n721), .B1(new_n333), .B2(new_n701), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n668), .A2(new_n692), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n710), .A2(new_n702), .A3(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1021), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT44), .B1(new_n711), .B2(new_n1025), .ZN(new_n1026));
  AND3_X1   g0826(.A1(new_n711), .A2(KEYINPUT44), .A3(new_n1025), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n709), .B(new_n1024), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1024), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1026), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n708), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n771), .B1(new_n1018), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT109), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n715), .B(KEYINPUT41), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1034), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n834), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1025), .B(new_n712), .C1(KEYINPUT42), .C2(new_n702), .ZN(new_n1039));
  OAI21_X1  g0839(.A(KEYINPUT42), .B1(new_n1025), .B2(new_n710), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n670), .A2(new_n701), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT43), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1003), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1039), .A2(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1043), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n708), .A2(new_n1021), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1006), .B1(new_n1038), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(G387));
  INV_X1    g0851(.A(new_n717), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n838), .A2(new_n1052), .B1(new_n354), .B2(new_n714), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n235), .A2(new_n391), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n445), .A2(new_n202), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n717), .B(new_n391), .C1(new_n244), .C2(new_n259), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n841), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1053), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n837), .B1(new_n1059), .B2(new_n844), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n786), .A2(new_n527), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G159), .B2(new_n814), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n304), .B1(new_n819), .B2(G150), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n796), .A2(G77), .B1(new_n797), .B2(new_n445), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n812), .A2(new_n202), .B1(new_n244), .B2(new_n807), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G97), .C2(new_n782), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n787), .A2(G283), .B1(new_n796), .B2(G294), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n814), .A2(G322), .B1(new_n797), .B2(G311), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n807), .B2(new_n612), .C1(new_n812), .C2(new_n821), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT110), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT49), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n322), .B1(G326), .B2(new_n819), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n620), .B2(new_n781), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1074), .B2(KEYINPUT49), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1067), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1060), .B1(new_n1079), .B2(new_n779), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n707), .B2(new_n776), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1018), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1081), .B1(new_n835), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n771), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n715), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1082), .A2(new_n771), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(G393));
  INV_X1    g0887(.A(new_n1032), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n835), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n844), .B1(new_n253), .B2(new_n207), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n242), .A2(new_n714), .A3(new_n322), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n836), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n812), .A2(new_n816), .B1(new_n821), .B2(new_n800), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT52), .Z(new_n1094));
  NOR2_X1   g0894(.A1(new_n795), .A2(new_n827), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n273), .B1(new_n789), .B2(new_n828), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n983), .A2(new_n612), .B1(new_n620), .B2(new_n786), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n784), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n370), .B2(new_n807), .ZN(new_n1099));
  INV_X1    g0899(.A(G159), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n812), .A2(new_n1100), .B1(new_n407), .B2(new_n800), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT51), .Z(new_n1102));
  OAI21_X1  g0902(.A(new_n322), .B1(new_n882), .B2(new_n789), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n983), .A2(new_n202), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n787), .A2(G77), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n244), .B2(new_n795), .ZN(new_n1106));
  NOR4_X1   g0906(.A1(new_n873), .A2(new_n1103), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n405), .B2(new_n807), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1094), .A2(new_n1099), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1092), .B1(new_n1109), .B2(new_n778), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1004), .B2(new_n1021), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1089), .A2(new_n1111), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1018), .A2(new_n770), .A3(new_n751), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n716), .B1(new_n1113), .B2(new_n1088), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1084), .A2(new_n1032), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(G390));
  OAI21_X1  g0917(.A(new_n942), .B1(new_n966), .B2(new_n967), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n863), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n743), .B1(KEYINPUT26), .B2(new_n740), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n739), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n958), .B1(new_n1121), .B2(new_n960), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n970), .B(KEYINPUT111), .Z(new_n1123));
  NAND3_X1  g0923(.A1(new_n1118), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n961), .B1(new_n684), .B2(new_n1119), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n971), .B1(new_n1125), .B2(new_n958), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1124), .B1(new_n1126), .B2(new_n969), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n770), .A2(new_n904), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n770), .A2(new_n904), .A3(KEYINPUT112), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT112), .B1(new_n770), .B2(new_n904), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1124), .B(new_n1133), .C1(new_n1126), .C2(new_n969), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n835), .A3(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1105), .B1(new_n800), .B2(new_n827), .C1(new_n354), .C2(new_n983), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n273), .B1(new_n789), .B2(new_n370), .C1(new_n337), .C2(new_n795), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n878), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n253), .B2(new_n807), .C1(new_n620), .C2(new_n812), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1140));
  NAND3_X1  g0940(.A1(new_n796), .A2(G150), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n273), .B1(new_n819), .B2(G125), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n1100), .C2(new_n786), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n797), .A2(G137), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n800), .A2(new_n1145), .B1(new_n781), .B2(new_n202), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1140), .B1(new_n796), .B2(G150), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  INV_X1    g0949(.A(G132), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1148), .B1(new_n807), .B2(new_n1149), .C1(new_n812), .C2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n779), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n837), .B(new_n1152), .C1(new_n405), .C2(new_n870), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n969), .B2(new_n775), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1135), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n958), .B1(new_n770), .B2(new_n859), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1129), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n960), .B1(new_n862), .B2(new_n863), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT112), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1128), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n770), .A2(new_n904), .A3(KEYINPUT112), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n960), .B1(new_n745), .B2(new_n863), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n752), .B(new_n858), .C1(new_n754), .C2(new_n769), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n958), .ZN(new_n1166));
  OAI21_X1  g0966(.A(KEYINPUT113), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1164), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(new_n1156), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT113), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1133), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1159), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n546), .A2(new_n770), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n653), .B(new_n1173), .C1(new_n750), .C2(new_n654), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT115), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1124), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n947), .A2(new_n949), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n951), .A2(new_n939), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n965), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n968), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n970), .B1(new_n1158), .B2(new_n959), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1177), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1134), .B1(new_n1184), .B2(new_n1128), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n716), .B1(new_n1176), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT114), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1125), .B1(new_n1129), .B2(new_n1156), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1170), .B1(new_n1133), .B2(new_n1169), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1166), .A2(new_n1131), .A3(new_n1132), .A4(KEYINPUT113), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1174), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1187), .B1(new_n1185), .B2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1175), .A2(KEYINPUT114), .A3(new_n1130), .A4(new_n1134), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1155), .B1(new_n1186), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(G378));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1174), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n411), .A2(new_n907), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT55), .Z(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n425), .B(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1205));
  XNOR2_X1  g1005(.A(new_n1204), .B(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n953), .A2(G330), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1206), .B1(new_n953), .B2(G330), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1208), .A2(new_n973), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n946), .A2(new_n952), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n944), .B1(new_n1118), .B2(new_n945), .ZN(new_n1212));
  OAI21_X1  g1012(.A(G330), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1206), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1215), .A2(new_n1207), .B1(new_n972), .B2(new_n964), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1210), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1199), .B1(new_n1200), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT121), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT121), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n1199), .C1(new_n1200), .C2(new_n1217), .ZN(new_n1221));
  OAI21_X1  g1021(.A(KEYINPUT120), .B1(new_n1210), .B2(new_n1216), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT120), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1215), .A2(new_n1207), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n1224), .B2(new_n973), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1199), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1196), .A2(new_n1192), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n716), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1219), .A2(new_n1221), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n836), .B1(new_n871), .B2(G50), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n819), .C2(G124), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n781), .B2(new_n790), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n983), .A2(new_n1150), .B1(new_n795), .B2(new_n1149), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n812), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(G128), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G150), .A2(new_n787), .B1(new_n814), .B2(G125), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT117), .Z(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n807), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1233), .B(new_n1238), .C1(G137), .C2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1232), .B1(new_n1241), .B2(KEYINPUT59), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(KEYINPUT59), .B2(new_n1241), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n786), .A2(new_n244), .B1(new_n795), .B2(new_n259), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n311), .B1(new_n789), .B2(new_n827), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1244), .A2(new_n322), .A3(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n814), .A2(G116), .B1(new_n797), .B2(G97), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1246), .B(new_n1247), .C1(new_n426), .C2(new_n781), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n807), .A2(new_n527), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n1234), .C2(G107), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n311), .B1(new_n304), .B2(new_n269), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1250), .A2(KEYINPUT58), .B1(new_n202), .B2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1243), .B(new_n1252), .C1(KEYINPUT58), .C2(new_n1250), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1230), .B1(new_n1253), .B2(new_n778), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1206), .B2(new_n775), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT119), .Z(new_n1256));
  INV_X1    g1056(.A(new_n1217), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1257), .B2(new_n835), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1229), .A2(new_n1258), .ZN(G375));
  NAND2_X1  g1059(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1176), .A2(new_n1035), .A3(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n958), .A2(new_n775), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1234), .A2(G283), .B1(G107), .B2(new_n1239), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n796), .A2(G97), .B1(new_n797), .B2(G116), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n370), .B2(new_n800), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n273), .B1(new_n789), .B2(new_n612), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1265), .A2(new_n1061), .A3(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1263), .B(new_n1267), .C1(new_n259), .C2(new_n783), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1234), .A2(G137), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1239), .A2(G150), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n800), .A2(new_n1150), .B1(new_n795), .B2(new_n1100), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G50), .B2(new_n787), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n983), .A2(new_n1149), .B1(new_n426), .B2(new_n781), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n304), .B(new_n1273), .C1(G128), .C2(new_n819), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1269), .A2(new_n1270), .A3(new_n1272), .A4(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n779), .B1(new_n1268), .B2(new_n1275), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n837), .B(new_n1276), .C1(new_n244), .C2(new_n870), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT122), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1172), .A2(new_n834), .B1(new_n1262), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1261), .A2(new_n1280), .ZN(G381));
  NOR4_X1   g1081(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1282));
  AND4_X1   g1082(.A1(new_n1050), .A2(new_n1282), .A3(new_n1280), .A4(new_n1261), .ZN(new_n1283));
  INV_X1    g1083(.A(G375), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n1284), .A3(new_n1197), .ZN(G407));
  NAND2_X1  g1085(.A1(new_n691), .A2(G213), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(new_n1197), .A3(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(G407), .A2(new_n1288), .A3(G213), .ZN(G409));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1229), .A2(G378), .A3(new_n1258), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1227), .A2(KEYINPUT123), .A3(new_n1035), .A4(new_n1257), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n835), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(new_n1255), .A3(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1200), .A2(new_n1217), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT123), .B1(new_n1296), .B2(new_n1035), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1197), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1291), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1286), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1172), .A2(KEYINPUT60), .A3(new_n1174), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n715), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1193), .A2(KEYINPUT60), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1260), .B2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n890), .B1(new_n1304), .B2(new_n1279), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1302), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1260), .B1(new_n1175), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(G384), .A3(new_n1280), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1290), .B1(new_n1300), .B2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G384), .B1(new_n1309), .B2(new_n1280), .ZN(new_n1313));
  AOI211_X1 g1113(.A(new_n890), .B(new_n1279), .C1(new_n1306), .C2(new_n1308), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT125), .B1(new_n1315), .B2(KEYINPUT124), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  OAI211_X1 g1117(.A(G2897), .B(new_n1287), .C1(new_n1311), .C2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT125), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1311), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1316), .A2(new_n1318), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1287), .A2(G2897), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1315), .B2(KEYINPUT124), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1319), .B1(new_n1311), .B2(new_n1317), .ZN(new_n1324));
  AOI211_X1 g1124(.A(KEYINPUT124), .B(KEYINPUT125), .C1(new_n1305), .C2(new_n1310), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1323), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1321), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT61), .B1(new_n1300), .B2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(G393), .B(G396), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(new_n1050), .B2(G390), .ZN(new_n1332));
  AOI211_X1 g1132(.A(new_n1006), .B(new_n1116), .C1(new_n1038), .C2(new_n1049), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1050), .A2(G390), .ZN(new_n1334));
  OAI22_X1  g1134(.A1(new_n1330), .A2(new_n1332), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(G387), .A2(new_n1116), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1050), .A2(G390), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1336), .A2(new_n1331), .A3(new_n1337), .A4(new_n1329), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1335), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1287), .B1(new_n1291), .B2(new_n1298), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(KEYINPUT63), .A3(new_n1315), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1312), .A2(new_n1328), .A3(new_n1339), .A4(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1340), .A2(new_n1343), .A3(new_n1315), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1321), .A2(new_n1326), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1345), .B1(new_n1340), .B2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1343), .B1(new_n1340), .B2(new_n1315), .ZN(new_n1348));
  NOR3_X1   g1148(.A1(new_n1344), .A2(new_n1347), .A3(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1342), .B1(new_n1349), .B2(new_n1339), .ZN(G405));
  NAND3_X1  g1150(.A1(G375), .A2(new_n1197), .A3(new_n1315), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1315), .B1(G375), .B2(new_n1197), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1338), .B(new_n1335), .C1(new_n1352), .C2(new_n1353), .ZN(new_n1354));
  AND2_X1   g1154(.A1(new_n1291), .A2(KEYINPUT127), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1353), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1356), .A2(new_n1339), .A3(new_n1351), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1354), .A2(new_n1355), .A3(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1355), .B1(new_n1354), .B2(new_n1357), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1358), .A2(new_n1359), .ZN(G402));
endmodule


