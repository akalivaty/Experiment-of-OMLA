//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT86), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT87), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G122), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G107), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT77), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n195), .B(new_n200), .C1(new_n197), .C2(new_n196), .ZN(new_n201));
  INV_X1    g015(.A(new_n195), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G104), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n199), .A2(new_n201), .A3(new_n203), .A4(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT4), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G101), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n210));
  INV_X1    g024(.A(G113), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT65), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(KEYINPUT2), .B2(G113), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT2), .A2(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G116), .ZN(new_n219));
  INV_X1    g033(.A(G116), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G119), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n222), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n215), .A3(new_n216), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n209), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT78), .B(G101), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(new_n205), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n199), .A2(new_n201), .A3(new_n229), .A4(new_n203), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT79), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n198), .A2(KEYINPUT77), .B1(KEYINPUT3), .B2(new_n202), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(KEYINPUT79), .A3(new_n201), .A4(new_n229), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n208), .B1(new_n207), .B2(G101), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n227), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(G101), .B1(new_n195), .B2(new_n205), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n219), .B(new_n221), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(G116), .A3(new_n218), .A4(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n244), .A3(G113), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT82), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT82), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n244), .A3(new_n247), .A4(G113), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n246), .A2(new_n225), .A3(new_n248), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n235), .A2(new_n238), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n193), .B1(new_n237), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n238), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n232), .B2(new_n234), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n249), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n235), .A2(new_n236), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n254), .B(new_n192), .C1(new_n255), .C2(new_n227), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(KEYINPUT6), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G143), .B(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n261), .A2(new_n259), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n260), .B1(new_n262), .B2(new_n258), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G125), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n266));
  INV_X1    g080(.A(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G143), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G146), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(KEYINPUT1), .A3(G146), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n271), .B(new_n272), .C1(G128), .C2(new_n258), .ZN(new_n273));
  INV_X1    g087(.A(G125), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  OR2_X1    g090(.A1(new_n276), .A2(KEYINPUT83), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(KEYINPUT83), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G224), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G953), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n283), .B(new_n193), .C1(new_n237), .C2(new_n250), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n257), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT84), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n244), .B(G113), .C1(new_n287), .C2(new_n222), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n225), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n253), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n192), .B(KEYINPUT8), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n246), .A2(new_n225), .A3(new_n248), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(new_n253), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n286), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n281), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n276), .B1(KEYINPUT85), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n296), .A2(KEYINPUT7), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n235), .A2(new_n238), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n249), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n301), .A2(KEYINPUT84), .A3(new_n290), .A4(new_n292), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n295), .A2(new_n299), .A3(new_n302), .A4(new_n256), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n191), .B1(new_n285), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n257), .A2(new_n282), .A3(new_n284), .ZN(new_n307));
  INV_X1    g121(.A(new_n190), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n307), .A2(new_n304), .A3(new_n303), .A4(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n188), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(G469), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n235), .A2(new_n236), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n209), .A2(new_n263), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G137), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(G134), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G131), .ZN(new_n319));
  INV_X1    g133(.A(G134), .ZN(new_n320));
  OAI211_X1 g134(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n320), .C2(G137), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(G134), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT11), .B1(new_n323), .B2(KEYINPUT64), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n319), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT64), .B1(new_n320), .B2(G137), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT11), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n318), .B1(new_n328), .B2(new_n321), .ZN(new_n329));
  INV_X1    g143(.A(G131), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n325), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT80), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n273), .A2(new_n238), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n232), .B2(new_n234), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI211_X1 g150(.A(KEYINPUT10), .B(new_n333), .C1(new_n232), .C2(new_n234), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n316), .B(new_n332), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G110), .B(G140), .ZN(new_n339));
  INV_X1    g153(.A(G953), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n340), .A2(G227), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n339), .B(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n273), .B1(new_n235), .B2(new_n238), .ZN(new_n345));
  OAI211_X1 g159(.A(KEYINPUT12), .B(new_n331), .C1(new_n345), .C2(new_n334), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n331), .B1(new_n345), .B2(new_n334), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT12), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n344), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n316), .B1(new_n336), .B2(new_n337), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n331), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n343), .B1(new_n352), .B2(new_n338), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n313), .B(new_n304), .C1(new_n350), .C2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n338), .A3(new_n343), .ZN(new_n355));
  INV_X1    g169(.A(new_n333), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n235), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT10), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n334), .A2(new_n335), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n358), .A2(new_n359), .B1(new_n314), .B2(new_n315), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n349), .A2(new_n346), .B1(new_n360), .B2(new_n332), .ZN(new_n361));
  OAI211_X1 g175(.A(G469), .B(new_n355), .C1(new_n361), .C2(new_n343), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n313), .A2(new_n304), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n354), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n310), .A2(new_n312), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT92), .B(G122), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G116), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n369));
  INV_X1    g183(.A(G122), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G116), .ZN(new_n371));
  OR2_X1    g185(.A1(KEYINPUT92), .A2(G122), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT92), .A2(G122), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n220), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n369), .B(G107), .C1(new_n371), .C2(new_n374), .ZN(new_n375));
  OAI221_X1 g189(.A(new_n368), .B1(KEYINPUT14), .B2(new_n204), .C1(G116), .C2(new_n370), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT93), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n269), .B2(G128), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n265), .A2(KEYINPUT93), .A3(G143), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n269), .A2(G128), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT94), .B(G134), .Z(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n382), .A2(new_n383), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n375), .A2(new_n376), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT13), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n388), .A2(G134), .B1(new_n381), .B2(new_n380), .ZN(new_n389));
  AND4_X1   g203(.A1(KEYINPUT13), .A2(new_n380), .A3(G134), .A4(new_n381), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n374), .A2(new_n371), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(new_n204), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n374), .A2(G107), .A3(new_n371), .ZN(new_n393));
  OAI22_X1  g207(.A1(new_n389), .A2(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G217), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n311), .A2(new_n395), .A3(G953), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n396), .B(KEYINPUT95), .Z(new_n397));
  NAND3_X1  g211(.A1(new_n386), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n386), .B2(new_n394), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT96), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI211_X1 g215(.A(KEYINPUT96), .B(new_n397), .C1(new_n394), .C2(new_n386), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n304), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT15), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G478), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n340), .A2(G952), .ZN(new_n407));
  NAND2_X1  g221(.A1(G234), .A2(G237), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(G902), .A3(G953), .ZN(new_n411));
  XOR2_X1   g225(.A(new_n411), .B(KEYINPUT97), .Z(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT21), .B(G898), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  NOR2_X1   g232(.A1(G475), .A2(G902), .ZN(new_n419));
  XNOR2_X1  g233(.A(G113), .B(G122), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n370), .A2(G113), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n211), .A2(G122), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n423), .A2(new_n424), .A3(new_n421), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(G104), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n420), .A2(new_n421), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n428), .A2(new_n425), .A3(new_n194), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(G237), .A2(G953), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G214), .ZN(new_n432));
  NOR2_X1   g246(.A1(KEYINPUT88), .A2(G143), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(KEYINPUT88), .A2(G143), .ZN(new_n435));
  NAND2_X1  g249(.A1(KEYINPUT88), .A2(G143), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n435), .A2(new_n436), .B1(new_n431), .B2(G214), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT18), .B(G131), .C1(new_n434), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n432), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(G214), .A3(new_n431), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT18), .A2(G131), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G125), .B(G140), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT72), .B1(new_n444), .B2(new_n267), .ZN(new_n445));
  INV_X1    g259(.A(G140), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G125), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n274), .A2(G140), .ZN(new_n448));
  AND4_X1   g262(.A1(KEYINPUT72), .A2(new_n447), .A3(new_n448), .A4(new_n267), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G140), .B1(new_n274), .B2(KEYINPUT71), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT71), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n446), .A3(G125), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n267), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n438), .B(new_n443), .C1(new_n450), .C2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n453), .A3(KEYINPUT16), .ZN(new_n456));
  OR3_X1    g270(.A1(new_n274), .A2(KEYINPUT16), .A3(G140), .ZN(new_n457));
  AOI21_X1  g271(.A(G146), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(G146), .A3(new_n457), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT17), .ZN(new_n461));
  OAI21_X1  g275(.A(G131), .B1(new_n434), .B2(new_n437), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n440), .A2(new_n330), .A3(new_n441), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n462), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n430), .B(new_n455), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n464), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n451), .A2(new_n453), .A3(KEYINPUT19), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n444), .A2(KEYINPUT19), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n267), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n460), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n430), .B1(new_n471), .B2(new_n455), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n466), .B1(new_n472), .B2(KEYINPUT90), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT90), .ZN(new_n474));
  AOI211_X1 g288(.A(new_n474), .B(new_n430), .C1(new_n455), .C2(new_n471), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n418), .B(new_n419), .C1(new_n473), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT91), .B1(new_n473), .B2(new_n475), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n455), .ZN(new_n479));
  INV_X1    g293(.A(new_n430), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n472), .A2(KEYINPUT90), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n466), .A4(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n478), .A2(new_n485), .A3(new_n419), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n477), .B1(new_n486), .B2(KEYINPUT20), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n455), .B1(new_n463), .B2(new_n465), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n480), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n466), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n304), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n491), .A2(G475), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n417), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n395), .B1(G234), .B2(new_n304), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT23), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n218), .B2(G128), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n218), .A2(G128), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n265), .A2(KEYINPUT23), .A3(G119), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT24), .B(G110), .Z(new_n501));
  XNOR2_X1  g315(.A(G119), .B(G128), .ZN(new_n502));
  OAI22_X1  g316(.A1(new_n500), .A2(G110), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n460), .C1(new_n445), .C2(new_n449), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n502), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n456), .A2(G146), .A3(new_n457), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(new_n458), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n500), .A2(KEYINPUT70), .A3(G110), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT70), .B1(new_n500), .B2(G110), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n504), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n504), .B(KEYINPUT73), .C1(new_n507), .C2(new_n510), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n340), .A2(G221), .A3(G234), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT22), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n317), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n511), .A2(new_n517), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n304), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT74), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n495), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n518), .A2(new_n519), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n518), .A2(KEYINPUT75), .A3(new_n519), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n495), .A2(G902), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(G472), .A2(G902), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT32), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G101), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT27), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n431), .A2(new_n540), .A3(G210), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n540), .B1(new_n431), .B2(G210), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT26), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT26), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n431), .A2(G210), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT27), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n547), .B2(new_n541), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n539), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT26), .B1(new_n542), .B2(new_n543), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n545), .A3(new_n541), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(G101), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n320), .A2(G137), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n330), .B1(new_n323), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n328), .A2(new_n321), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(new_n319), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n331), .A2(new_n263), .B1(new_n273), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n223), .A2(new_n225), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT31), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n558), .A2(KEYINPUT30), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n258), .B1(new_n261), .B2(new_n259), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n258), .A2(new_n259), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n554), .B1(new_n322), .B2(new_n324), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G131), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n565), .B1(new_n567), .B2(new_n325), .ZN(new_n568));
  INV_X1    g382(.A(new_n555), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n325), .A2(new_n273), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT30), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n226), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n560), .B(new_n561), .C1(new_n562), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT66), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n331), .A2(new_n263), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n570), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT30), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(KEYINPUT30), .A3(new_n570), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n226), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT66), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n561), .A4(new_n560), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n576), .A2(new_n226), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n566), .A2(G131), .B1(new_n556), .B2(new_n319), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n559), .B(new_n570), .C1(new_n587), .C2(new_n565), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n585), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT28), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n553), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n560), .B1(new_n562), .B2(new_n572), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT31), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n538), .B1(new_n583), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT69), .ZN(new_n598));
  INV_X1    g412(.A(new_n588), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n559), .B1(new_n575), .B2(new_n570), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n584), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n591), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n602), .A2(new_n553), .B1(KEYINPUT31), .B2(new_n594), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n574), .A2(new_n582), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT69), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n538), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n580), .A2(new_n588), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n553), .ZN(new_n610));
  INV_X1    g424(.A(new_n553), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n602), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT29), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n590), .B1(new_n586), .B2(new_n588), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n592), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(KEYINPUT29), .A3(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n304), .ZN(new_n617));
  OAI21_X1  g431(.A(G472), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n536), .B1(new_n603), .B2(new_n604), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT68), .A3(new_n537), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT68), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n619), .B2(KEYINPUT32), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n608), .A2(new_n618), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n366), .A2(new_n494), .A3(new_n534), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(new_n228), .ZN(G3));
  NAND2_X1  g440(.A1(new_n386), .A2(new_n394), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n627), .A2(KEYINPUT98), .A3(new_n397), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n397), .B1(new_n627), .B2(KEYINPUT98), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT33), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(G478), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(G902), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n401), .A2(new_n402), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n630), .B(new_n632), .C1(new_n633), .C2(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n403), .A2(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n636), .B(new_n416), .C1(new_n487), .C2(new_n492), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n190), .B1(new_n285), .B2(new_n305), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n188), .B1(new_n639), .B2(new_n309), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n638), .A2(new_n640), .A3(KEYINPUT99), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT99), .B1(new_n638), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n312), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n338), .B1(new_n360), .B2(new_n587), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n342), .ZN(new_n646));
  INV_X1    g460(.A(new_n346), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n357), .B1(new_n273), .B2(new_n253), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT12), .B1(new_n648), .B2(new_n331), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n338), .B(new_n343), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n363), .B1(new_n651), .B2(new_n313), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n644), .B1(new_n652), .B2(new_n362), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n605), .A2(new_n304), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n619), .B1(new_n654), .B2(G472), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n534), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n643), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT100), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n657), .B(new_n659), .ZN(G6));
  NAND2_X1  g474(.A1(new_n639), .A2(new_n309), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n187), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT101), .B1(new_n486), .B2(KEYINPUT20), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(KEYINPUT20), .B2(new_n486), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n406), .A2(new_n492), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n478), .A2(new_n485), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n666), .A2(KEYINPUT101), .A3(new_n418), .A4(new_n419), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n664), .A2(new_n665), .A3(new_n416), .A4(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n662), .B1(KEYINPUT102), .B2(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n656), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT103), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n672), .B(new_n674), .ZN(G9));
  NAND2_X1  g489(.A1(new_n513), .A2(new_n514), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n517), .A2(KEYINPUT36), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n676), .B(new_n677), .Z(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n531), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n525), .A2(new_n679), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n417), .A2(new_n493), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n366), .A2(new_n655), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  OR2_X1    g498(.A1(new_n412), .A2(G900), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n409), .B(KEYINPUT104), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n664), .A2(new_n665), .A3(new_n667), .A4(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AOI221_X4 g503(.A(new_n188), .B1(new_n525), .B2(new_n679), .C1(new_n639), .C2(new_n309), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n624), .A2(new_n689), .A3(new_n690), .A4(new_n653), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  XNOR2_X1  g506(.A(new_n687), .B(KEYINPUT39), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n653), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT40), .Z(new_n695));
  AOI21_X1  g509(.A(new_n553), .B1(new_n580), .B2(new_n588), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n586), .A2(new_n588), .A3(new_n553), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n304), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT105), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n608), .A2(new_n621), .A3(new_n623), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n306), .A2(new_n309), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT38), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n486), .A2(KEYINPUT20), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n476), .ZN(new_n706));
  INV_X1    g520(.A(new_n492), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n406), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n704), .A2(new_n188), .A3(new_n680), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n695), .A2(new_n701), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  OAI211_X1 g526(.A(new_n636), .B(new_n687), .C1(new_n487), .C2(new_n492), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n624), .A2(new_n690), .A3(new_n653), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  INV_X1    g530(.A(new_n344), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n349), .A2(new_n346), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n717), .A2(new_n718), .B1(new_n645), .B2(new_n342), .ZN(new_n719));
  OAI21_X1  g533(.A(G469), .B1(new_n719), .B2(G902), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n312), .A3(new_n354), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n720), .A2(KEYINPUT106), .A3(new_n312), .A4(new_n354), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n624), .A3(new_n534), .A4(new_n724), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n643), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  AND2_X1   g542(.A1(new_n721), .A2(new_n722), .ZN(new_n729));
  INV_X1    g543(.A(new_n724), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n624), .A2(new_n534), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n732), .A3(new_n670), .A4(new_n669), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  NOR2_X1   g548(.A1(new_n662), .A2(new_n721), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n624), .A3(new_n681), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  NAND3_X1  g551(.A1(new_n640), .A2(new_n416), .A3(new_n708), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n729), .A2(new_n730), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n654), .A2(KEYINPUT108), .A3(G472), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  AOI21_X1  g555(.A(G902), .B1(new_n603), .B2(new_n604), .ZN(new_n742));
  INV_X1    g556(.A(G472), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n604), .A2(new_n595), .ZN(new_n746));
  OR3_X1    g560(.A1(new_n614), .A2(new_n592), .A3(KEYINPUT107), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT107), .B1(new_n614), .B2(new_n592), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n553), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n536), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n745), .A2(new_n534), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n750), .B1(new_n740), .B2(new_n744), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(KEYINPUT109), .A3(new_n534), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n739), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  AND3_X1   g573(.A1(new_n745), .A2(new_n680), .A3(new_n751), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n735), .A3(new_n714), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  OAI211_X1 g576(.A(new_n618), .B(new_n597), .C1(KEYINPUT32), .C2(new_n619), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(new_n534), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n644), .A2(new_n188), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n306), .A2(new_n309), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n362), .A2(KEYINPUT110), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n338), .B1(new_n647), .B2(new_n649), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n342), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n770), .A3(G469), .A4(new_n355), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n767), .A2(new_n354), .A3(new_n771), .A4(new_n364), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n764), .A2(new_n773), .A3(KEYINPUT42), .A4(new_n714), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n534), .A3(new_n624), .A4(new_n714), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT42), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT112), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n330), .ZN(G33));
  NAND3_X1  g596(.A1(new_n732), .A2(new_n689), .A3(new_n773), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n493), .A2(new_n636), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT43), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(KEYINPUT43), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n620), .B1(new_n743), .B2(new_n742), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(new_n680), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(KEYINPUT44), .A3(new_n791), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n702), .A2(new_n188), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT45), .B1(new_n769), .B2(new_n355), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n313), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n769), .A2(KEYINPUT45), .A3(new_n355), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n363), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n354), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n312), .ZN(new_n806));
  INV_X1    g620(.A(new_n693), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n798), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n805), .A2(KEYINPUT113), .A3(new_n312), .A4(new_n693), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n797), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(new_n317), .ZN(G39));
  NAND2_X1  g625(.A1(new_n806), .A2(KEYINPUT47), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n805), .A2(new_n813), .A3(new_n312), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n796), .A2(new_n533), .A3(new_n714), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n624), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  NAND2_X1  g632(.A1(new_n720), .A2(new_n354), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n820), .A2(new_n821), .A3(new_n785), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n534), .A2(new_n765), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT114), .ZN(new_n824));
  INV_X1    g638(.A(new_n701), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n704), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n310), .A2(new_n365), .A3(new_n312), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n406), .B(KEYINPUT117), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n493), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n534), .A2(new_n655), .A3(new_n416), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n755), .A2(KEYINPUT109), .A3(new_n534), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT109), .B1(new_n755), .B2(new_n534), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n708), .A2(new_n661), .A3(new_n187), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n723), .A3(new_n416), .A4(new_n724), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n832), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n682), .B(new_n736), .C1(new_n643), .C2(new_n725), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n671), .A2(new_n725), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n790), .A2(new_n533), .A3(new_n415), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n636), .B1(new_n487), .B2(new_n492), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT115), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n366), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n625), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n842), .B1(new_n625), .B2(new_n846), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n624), .A2(new_n653), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n664), .A2(new_n667), .ZN(new_n852));
  INV_X1    g666(.A(new_n687), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n828), .A2(new_n852), .A3(new_n492), .A4(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n851), .A2(new_n680), .A3(new_n854), .A4(new_n796), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n760), .A2(new_n773), .A3(new_n714), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n783), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n841), .A2(new_n780), .A3(new_n850), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n680), .A2(new_n644), .A3(new_n853), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n836), .A2(new_n701), .A3(new_n772), .A4(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n761), .A2(new_n691), .A3(new_n862), .A4(new_n715), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n640), .A2(new_n680), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n688), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n714), .A2(new_n640), .A3(new_n680), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n653), .B(new_n624), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT52), .A3(new_n761), .A4(new_n862), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT53), .B1(new_n860), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n865), .A2(KEYINPUT119), .A3(new_n870), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n880), .A2(new_n859), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT54), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n880), .B2(new_n859), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n831), .B1(new_n739), .B2(new_n757), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n682), .A2(new_n736), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n726), .A3(new_n733), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n625), .A2(new_n846), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT116), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n847), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n774), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n775), .A2(new_n777), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT111), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n857), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n891), .A4(new_n897), .ZN(new_n898));
  XOR2_X1   g712(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n899));
  NAND3_X1  g713(.A1(new_n884), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n883), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n721), .A2(new_n702), .A3(new_n188), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n410), .A2(new_n902), .A3(new_n534), .A4(new_n825), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n493), .A3(new_n635), .A4(new_n634), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n788), .A2(new_n686), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n902), .A3(new_n760), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n905), .A2(new_n757), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n721), .A2(new_n187), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n704), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(KEYINPUT50), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT50), .B1(new_n908), .B2(new_n910), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n907), .B(KEYINPUT51), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n819), .A2(new_n312), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n812), .B2(new_n814), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n908), .A2(new_n796), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT122), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n904), .A2(KEYINPUT51), .A3(new_n906), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n908), .A2(new_n910), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT50), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n923), .B2(new_n911), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n924), .B(new_n925), .C1(new_n916), .C2(new_n917), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT51), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT121), .B1(new_n912), .B2(new_n913), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n923), .A2(new_n911), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n931), .A3(new_n907), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n932), .B2(new_n918), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n908), .A2(new_n735), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n903), .B(new_n636), .C1(new_n492), .C2(new_n487), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n905), .A2(new_n764), .A3(new_n902), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT123), .B(KEYINPUT48), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n935), .B(new_n407), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n934), .B(new_n938), .C1(new_n936), .C2(new_n937), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n927), .A2(new_n933), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n901), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(G952), .A2(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n826), .B1(new_n941), .B2(new_n942), .ZN(G75));
  NAND2_X1  g757(.A1(new_n257), .A2(new_n284), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n282), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT124), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT55), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n304), .B1(new_n884), .B2(new_n898), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n190), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT56), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n340), .A2(G952), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n947), .A2(new_n950), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n948), .B2(new_n191), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(G51));
  XNOR2_X1  g769(.A(new_n363), .B(KEYINPUT57), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n884), .A2(new_n898), .A3(new_n899), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n899), .B1(new_n884), .B2(new_n898), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n719), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n948), .A2(new_n801), .A3(new_n800), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n952), .B1(new_n961), .B2(new_n962), .ZN(G54));
  NAND3_X1  g777(.A1(new_n948), .A2(KEYINPUT58), .A3(G475), .ZN(new_n964));
  INV_X1    g778(.A(new_n666), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n952), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n948), .A2(KEYINPUT58), .A3(G475), .A4(new_n666), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(G60));
  OR2_X1    g783(.A1(new_n633), .A2(KEYINPUT33), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n970), .A2(new_n630), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n972));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n971), .B1(new_n901), .B2(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n971), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n957), .B2(new_n958), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n967), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n975), .A2(new_n978), .ZN(G63));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT60), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n879), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT119), .B1(new_n865), .B2(new_n870), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT53), .B1(new_n860), .B2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n865), .A2(new_n873), .A3(new_n870), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n873), .B1(new_n865), .B2(new_n870), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n989), .A2(new_n859), .A3(new_n881), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n982), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n530), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(KEYINPUT126), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n981), .B1(new_n884), .B2(new_n898), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(new_n530), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n952), .B1(new_n995), .B2(new_n678), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n993), .A2(new_n996), .A3(new_n997), .A4(KEYINPUT61), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n678), .B(new_n982), .C1(new_n986), .C2(new_n990), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n967), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n995), .A2(new_n530), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n998), .A2(new_n1003), .ZN(G66));
  NOR3_X1   g818(.A1(new_n414), .A2(new_n280), .A3(new_n340), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n891), .B2(new_n340), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n944), .B1(G898), .B2(new_n340), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(G69));
  NAND2_X1  g822(.A1(new_n578), .A2(new_n579), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n468), .A2(new_n469), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G900), .A2(G953), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n869), .A2(new_n761), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT127), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1014), .A2(new_n783), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n808), .A2(new_n809), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n764), .A2(new_n836), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n797), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1015), .A2(new_n1019), .A3(new_n780), .A4(new_n817), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1011), .B(new_n1012), .C1(new_n1020), .C2(G953), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1014), .A2(new_n711), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(KEYINPUT62), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT62), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1014), .A2(new_n1024), .A3(new_n711), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n845), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n694), .B1(new_n1027), .B2(new_n829), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1028), .A2(new_n732), .A3(new_n796), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n817), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1030), .A2(new_n810), .ZN(new_n1031));
  AOI21_X1  g845(.A(G953), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1021), .B1(new_n1032), .B2(new_n1011), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n340), .B1(G227), .B2(G900), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1034), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1021), .B(new_n1036), .C1(new_n1032), .C2(new_n1011), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1035), .A2(new_n1037), .ZN(G72));
  NAND4_X1  g852(.A1(new_n1031), .A2(new_n1023), .A3(new_n891), .A4(new_n1025), .ZN(new_n1039));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  NAND2_X1  g855(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n952), .B1(new_n1042), .B2(new_n696), .ZN(new_n1043));
  INV_X1    g857(.A(new_n891), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1041), .B1(new_n1020), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1045), .A2(new_n609), .A3(new_n553), .ZN(new_n1046));
  AND2_X1   g860(.A1(new_n610), .A2(new_n1041), .ZN(new_n1047));
  OAI221_X1 g861(.A(new_n1047), .B1(new_n609), .B2(new_n553), .C1(new_n876), .C2(new_n882), .ZN(new_n1048));
  AND3_X1   g862(.A1(new_n1043), .A2(new_n1046), .A3(new_n1048), .ZN(G57));
endmodule


