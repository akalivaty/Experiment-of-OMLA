//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT67), .B(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g0023(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n214), .B1(KEYINPUT1), .B2(new_n223), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT68), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G13), .ZN(new_n245));
  NOR3_X1   g0045(.A1(new_n245), .A2(new_n209), .A3(G1), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G1), .A2(G13), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n201), .B1(new_n208), .B2(G20), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(new_n251), .B1(new_n201), .B2(new_n246), .ZN(new_n252));
  OR2_X1    g0052(.A1(new_n252), .A2(KEYINPUT70), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(KEYINPUT70), .ZN(new_n254));
  OAI21_X1  g0054(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n255));
  INV_X1    g0055(.A(G150), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n209), .A2(G33), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n255), .B1(new_n256), .B2(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n253), .A2(new_n254), .B1(new_n249), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT9), .ZN(new_n263));
  INV_X1    g0063(.A(new_n215), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n264), .A2(new_n267), .B1(new_n273), .B2(G223), .ZN(new_n274));
  INV_X1    g0074(.A(G222), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n276), .B(new_n278), .C1(new_n265), .C2(new_n266), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n274), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n248), .B1(G33), .B2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(G1), .B(G13), .C1(new_n270), .C2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n286), .A3(G274), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n283), .ZN(new_n288));
  INV_X1    g0088(.A(G226), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(G190), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n282), .A2(new_n291), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G200), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n263), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n253), .A2(new_n254), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n261), .A2(new_n249), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT74), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT74), .B1(new_n262), .B2(KEYINPUT9), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n295), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n295), .B2(new_n303), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n260), .ZN(new_n308));
  INV_X1    g0108(.A(G68), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n308), .A2(G77), .B1(G20), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n201), .B2(new_n258), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n246), .A2(new_n309), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT12), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n208), .A2(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n250), .A2(G68), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n312), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT11), .B1(new_n311), .B2(new_n249), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n271), .A2(new_n272), .ZN(new_n320));
  INV_X1    g0120(.A(G232), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(new_n268), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n320), .A2(new_n322), .B1(G33), .B2(G97), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT69), .B(G1698), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n324), .A3(G226), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n286), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G238), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n287), .B1(new_n288), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n327), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n332), .A2(G190), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT13), .B1(new_n326), .B2(new_n329), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n319), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n336), .A3(new_n334), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n327), .A2(new_n330), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(KEYINPUT75), .A3(KEYINPUT13), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(G200), .A3(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n337), .A2(G169), .A3(new_n339), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n332), .A2(G179), .A3(new_n334), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n337), .A2(new_n339), .A3(new_n345), .A4(G169), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n341), .B1(new_n319), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n287), .B1(new_n288), .B2(new_n216), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n320), .A2(G238), .A3(G1698), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT71), .B(G107), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n350), .B1(new_n320), .B2(new_n351), .C1(new_n321), .C2(new_n279), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(new_n352), .B2(new_n281), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n249), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT15), .B(G87), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT72), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n308), .ZN(new_n360));
  INV_X1    g0160(.A(new_n259), .ZN(new_n361));
  AOI22_X1  g0161(.A1(G20), .A2(new_n264), .B1(new_n361), .B2(new_n257), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n356), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n250), .A2(G77), .A3(new_n315), .ZN(new_n364));
  INV_X1    g0164(.A(new_n246), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n264), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n353), .A2(G190), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n355), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n363), .A2(new_n366), .B1(new_n353), .B2(G169), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n370), .A2(KEYINPUT73), .B1(new_n371), .B2(new_n353), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT73), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n373), .B1(new_n353), .B2(G169), .C1(new_n363), .C2(new_n366), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n369), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G169), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n262), .B1(new_n293), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G179), .B2(new_n293), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n307), .A2(new_n348), .A3(new_n375), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n202), .A2(new_n309), .ZN(new_n380));
  NOR2_X1   g0180(.A1(G58), .A2(G68), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n257), .A2(G159), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT16), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NOR4_X1   g0187(.A1(new_n265), .A2(new_n266), .A3(new_n387), .A4(G20), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT76), .B1(new_n265), .B2(new_n266), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT76), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n271), .A2(new_n390), .A3(new_n272), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n391), .A3(new_n209), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(new_n387), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n386), .B1(new_n393), .B2(new_n309), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT77), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT77), .B(new_n386), .C1(new_n393), .C2(new_n309), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n387), .B1(new_n320), .B2(G20), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n309), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n385), .B1(new_n401), .B2(new_n384), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n249), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT78), .ZN(new_n406));
  INV_X1    g0206(.A(new_n250), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n361), .A2(new_n315), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n407), .A2(new_n408), .B1(new_n365), .B2(new_n361), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n403), .B1(new_n396), .B2(new_n397), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT78), .B1(new_n412), .B2(new_n409), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT79), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n276), .A2(new_n278), .A3(G223), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G226), .A2(G1698), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n267), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G87), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n270), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n281), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n281), .A2(new_n284), .ZN(new_n421));
  INV_X1    g0221(.A(G274), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n281), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g0223(.A1(G232), .A2(new_n421), .B1(new_n423), .B2(new_n284), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n414), .B1(new_n425), .B2(new_n371), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n420), .A2(new_n424), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n376), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n427), .A2(KEYINPUT79), .A3(G179), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n411), .A2(new_n413), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT18), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n411), .A2(new_n413), .A3(new_n435), .A4(new_n432), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n409), .B1(new_n398), .B2(new_n404), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n420), .A2(new_n424), .A3(G190), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n425), .B2(new_n354), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT17), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT17), .ZN(new_n442));
  NOR4_X1   g0242(.A1(new_n412), .A2(new_n442), .A3(new_n439), .A4(new_n409), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n434), .A2(new_n436), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n379), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT84), .ZN(new_n447));
  OAI211_X1 g0247(.A(G264), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT82), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n320), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G257), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n271), .B2(new_n272), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n454), .A2(new_n324), .B1(new_n267), .B2(G303), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n286), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n281), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G270), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n459), .A2(new_n286), .A3(G274), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(G200), .B1(new_n456), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n246), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n208), .A2(G33), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n250), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n468), .B2(new_n465), .ZN(new_n469));
  AOI21_X1  g0269(.A(G20), .B1(new_n270), .B2(G97), .ZN(new_n470));
  INV_X1    g0270(.A(G283), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n270), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(G20), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n249), .A2(KEYINPUT83), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT83), .B1(new_n249), .B2(new_n473), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT20), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT20), .B(new_n472), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n447), .B1(new_n464), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n459), .A2(new_n458), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n460), .A2(G270), .B1(new_n483), .B2(new_n423), .ZN(new_n484));
  OAI21_X1  g0284(.A(G257), .B1(new_n265), .B2(new_n266), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n276), .A2(new_n278), .ZN(new_n486));
  INV_X1    g0286(.A(G303), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n485), .A2(new_n486), .B1(new_n320), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n450), .B2(new_n451), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n484), .B1(new_n489), .B2(new_n286), .ZN(new_n490));
  INV_X1    g0290(.A(G190), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n481), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n464), .A2(new_n447), .A3(new_n480), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n478), .A2(new_n479), .ZN(new_n497));
  INV_X1    g0297(.A(new_n469), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n499), .A2(KEYINPUT21), .A3(G169), .A4(new_n490), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  OAI21_X1  g0301(.A(G169), .B1(new_n456), .B2(new_n463), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n480), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n456), .A2(new_n463), .A3(new_n371), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n500), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT85), .B1(new_n496), .B2(new_n506), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n494), .A2(new_n481), .A3(new_n492), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n500), .A2(new_n503), .A3(new_n505), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT85), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n351), .ZN(new_n513));
  INV_X1    g0313(.A(new_n399), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n388), .ZN(new_n515));
  INV_X1    g0315(.A(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(KEYINPUT6), .A3(G97), .ZN(new_n517));
  XOR2_X1   g0317(.A(G97), .B(G107), .Z(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n356), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n246), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n468), .B2(new_n522), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n482), .A2(G257), .A3(new_n286), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n462), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n273), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n279), .B2(new_n216), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n320), .A2(new_n324), .A3(KEYINPUT4), .A4(G244), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n527), .B1(new_n532), .B2(new_n281), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n371), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n533), .A2(G169), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n525), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n521), .A2(new_n524), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n533), .A2(KEYINPUT80), .ZN(new_n538));
  OAI21_X1  g0338(.A(G200), .B1(new_n533), .B2(KEYINPUT80), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT81), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n533), .A2(new_n541), .A3(G190), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n533), .B2(G190), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n536), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n458), .A2(G250), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n457), .A2(G1), .A3(G274), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n546), .A2(new_n281), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n320), .A2(new_n324), .A3(G238), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G116), .ZN(new_n550));
  OAI211_X1 g0350(.A(G244), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n548), .B1(new_n552), .B2(new_n281), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n371), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n320), .A2(new_n209), .A3(G68), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n260), .B2(new_n522), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(G87), .A2(G97), .ZN(new_n559));
  NAND3_X1  g0359(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n351), .A2(new_n559), .B1(new_n209), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n249), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n357), .A2(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n357), .A2(KEYINPUT72), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n246), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n563), .A2(new_n250), .A3(new_n564), .A4(new_n467), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n554), .B(new_n568), .C1(G169), .C2(new_n553), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n551), .A2(new_n550), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n286), .B1(new_n570), .B2(new_n549), .ZN(new_n571));
  OAI21_X1  g0371(.A(G200), .B1(new_n571), .B2(new_n548), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n553), .A2(G190), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n351), .A2(new_n559), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n560), .A2(new_n209), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n557), .A3(new_n555), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n249), .B1(new_n565), .B2(new_n246), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n250), .A2(G87), .A3(new_n467), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n572), .A2(new_n573), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n569), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT87), .B1(new_n582), .B2(KEYINPUT86), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(KEYINPUT87), .B2(new_n582), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n209), .B(G87), .C1(new_n265), .C2(new_n266), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT23), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n516), .A3(G20), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n465), .B2(new_n260), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n351), .A2(G20), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(KEYINPUT23), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n585), .B1(KEYINPUT86), .B2(new_n582), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT24), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n586), .A2(new_n591), .A3(new_n595), .A4(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n249), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT25), .B1(new_n246), .B2(new_n516), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n516), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n516), .B2(new_n468), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n320), .A2(G257), .A3(G1698), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G294), .ZN(new_n606));
  INV_X1    g0406(.A(G250), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n279), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n281), .B1(G264), .B2(new_n460), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(G190), .A3(new_n462), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n281), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n460), .A2(G264), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n462), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G200), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n598), .A2(new_n604), .A3(new_n610), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n376), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n609), .A2(new_n371), .A3(new_n462), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n356), .B1(new_n594), .B2(new_n596), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n603), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n581), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n545), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n446), .A2(new_n512), .A3(new_n621), .ZN(G372));
  INV_X1    g0422(.A(new_n569), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n536), .B(new_n615), .C1(new_n540), .C2(new_n544), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n506), .B2(new_n619), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT88), .B1(new_n578), .B2(new_n579), .ZN(new_n626));
  AND4_X1   g0426(.A1(KEYINPUT88), .A2(new_n562), .A3(new_n566), .A4(new_n579), .ZN(new_n627));
  OAI211_X1 g0427(.A(KEYINPUT89), .B(new_n572), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n573), .ZN(new_n629));
  INV_X1    g0429(.A(new_n572), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n562), .A2(new_n566), .A3(new_n579), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT88), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n578), .A2(KEYINPUT88), .A3(new_n579), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(KEYINPUT89), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n569), .B1(new_n629), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n623), .B1(new_n625), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n536), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n640), .B(new_n569), .C1(new_n629), .C2(new_n636), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(KEYINPUT90), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n640), .A2(new_n581), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT90), .B1(new_n641), .B2(new_n642), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n639), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n446), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n378), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n430), .B1(new_n426), .B2(new_n428), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT18), .B1(new_n437), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n437), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(new_n435), .A3(new_n432), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n372), .A2(new_n374), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n335), .A2(new_n340), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n656), .A2(new_n657), .B1(new_n347), .B2(new_n319), .ZN(new_n658));
  INV_X1    g0458(.A(new_n444), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n652), .B(new_n654), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n650), .B1(new_n660), .B2(new_n307), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n649), .A2(new_n661), .ZN(G369));
  NAND3_X1  g0462(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT91), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  INV_X1    g0466(.A(G213), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(KEYINPUT92), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(KEYINPUT92), .ZN(new_n671));
  OAI211_X1 g0471(.A(G343), .B(new_n668), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n512), .B1(new_n480), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n672), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n509), .A2(new_n499), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n619), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n674), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n674), .B1(new_n618), .B2(new_n603), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n615), .A2(new_n679), .A3(new_n619), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n676), .A2(G330), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n509), .A2(new_n672), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT93), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n681), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n672), .A2(KEYINPUT94), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n672), .A2(KEYINPUT94), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n677), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n682), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n212), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n574), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n225), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT95), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  MUX2_X1   g0499(.A(new_n644), .B(new_n641), .S(KEYINPUT26), .Z(new_n700));
  NAND2_X1  g0500(.A1(new_n506), .A2(new_n619), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n540), .A2(new_n544), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n702), .A3(new_n536), .A4(new_n615), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n569), .B1(new_n703), .B2(new_n637), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT29), .B(new_n672), .C1(new_n700), .C2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n648), .A2(new_n688), .ZN(new_n706));
  XOR2_X1   g0506(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G330), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n621), .B(new_n688), .C1(new_n507), .C2(new_n511), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n533), .A2(new_n609), .A3(new_n553), .ZN(new_n711));
  OAI211_X1 g0511(.A(G179), .B(new_n484), .C1(new_n489), .C2(new_n286), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT30), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n609), .A2(new_n553), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(new_n504), .A4(new_n533), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n553), .A2(G179), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n718), .A2(new_n490), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n533), .B1(new_n462), .B2(new_n609), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT31), .B1(new_n722), .B2(new_n674), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n713), .A2(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n724), .A2(new_n688), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n709), .B1(new_n710), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n708), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n699), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n676), .A2(G330), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT97), .Z(new_n733));
  NAND2_X1  g0533(.A1(new_n676), .A2(G330), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n245), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n208), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n733), .B(new_n734), .C1(new_n693), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n693), .A2(new_n737), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT98), .Z(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n692), .A2(new_n267), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n742), .A2(G355), .B1(new_n465), .B2(new_n692), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n389), .A2(new_n391), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n692), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G45), .B2(new_n226), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n240), .A2(new_n457), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n248), .B1(G20), .B2(new_n376), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n741), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n752), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n209), .A2(new_n371), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n757), .A2(new_n491), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G322), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n209), .A2(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n759), .A2(new_n760), .B1(new_n487), .B2(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n320), .B(new_n763), .C1(G311), .C2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n761), .A2(new_n491), .A3(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n756), .A2(G200), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT99), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(KEYINPUT33), .B(G317), .Z(new_n771));
  OAI221_X1 g0571(.A(new_n765), .B1(new_n471), .B2(new_n766), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n761), .A2(new_n491), .A3(new_n354), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT100), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n772), .B1(G329), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n768), .A2(new_n491), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n491), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n209), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n780), .A2(G326), .B1(G294), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT102), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n320), .B1(new_n762), .B2(new_n418), .C1(new_n516), .C2(new_n766), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT101), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n770), .B2(new_n309), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G50), .B2(new_n780), .ZN(new_n789));
  INV_X1    g0589(.A(new_n764), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n202), .A2(new_n759), .B1(new_n790), .B2(new_n215), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n782), .A2(new_n522), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n778), .A2(G159), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(KEYINPUT101), .B2(new_n786), .C1(KEYINPUT32), .C2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(KEYINPUT32), .B2(new_n794), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n779), .A2(new_n785), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n751), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n754), .B1(new_n755), .B2(new_n797), .C1(new_n676), .C2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n738), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n370), .A2(KEYINPUT73), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n353), .A2(new_n371), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n367), .A2(new_n672), .ZN(new_n804));
  AND4_X1   g0604(.A1(new_n374), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n804), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(new_n375), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n688), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n648), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n706), .B2(new_n808), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n739), .B1(new_n812), .B2(new_n729), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n729), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n752), .A2(new_n749), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n740), .B1(G77), .B2(new_n816), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n790), .A2(new_n465), .B1(new_n516), .B2(new_n762), .ZN(new_n818));
  INV_X1    g0618(.A(G294), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n267), .B1(new_n759), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n766), .A2(new_n418), .ZN(new_n821));
  NOR4_X1   g0621(.A1(new_n818), .A2(new_n820), .A3(new_n792), .A4(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n769), .A2(G283), .B1(new_n778), .B2(G311), .ZN(new_n823));
  INV_X1    g0623(.A(new_n780), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n823), .C1(new_n487), .C2(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G143), .A2(new_n758), .B1(new_n764), .B2(G159), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n824), .B2(new_n827), .C1(new_n256), .C2(new_n770), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  INV_X1    g0629(.A(new_n744), .ZN(new_n830));
  INV_X1    g0630(.A(new_n762), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(G50), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n766), .A2(new_n309), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G58), .B2(new_n783), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n832), .B(new_n834), .C1(new_n835), .C2(new_n777), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n825), .B1(new_n829), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n817), .B1(new_n837), .B2(new_n752), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n808), .B2(new_n750), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n814), .A2(new_n839), .ZN(G384));
  NOR2_X1   g0640(.A1(new_n735), .A2(new_n208), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n382), .B(new_n383), .C1(new_n393), .C2(new_n309), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n356), .B1(new_n842), .B2(new_n385), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n409), .B1(new_n398), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n670), .A2(new_n671), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n668), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n445), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n405), .A2(new_n410), .A3(new_n440), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n651), .B2(new_n844), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n850), .B2(new_n847), .ZN(new_n851));
  INV_X1    g0651(.A(new_n846), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n411), .A2(new_n413), .A3(new_n852), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n412), .A2(new_n409), .A3(new_n439), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n433), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT104), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n848), .A2(KEYINPUT104), .A3(KEYINPUT38), .A4(new_n857), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n854), .A2(KEYINPUT17), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n849), .A2(new_n442), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n654), .A2(new_n862), .A3(new_n863), .A4(new_n652), .ZN(new_n864));
  INV_X1    g0664(.A(new_n853), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n856), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n854), .B1(new_n653), .B2(new_n432), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n853), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n860), .A2(new_n861), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n724), .A2(new_n725), .A3(new_n672), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n723), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n710), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n347), .A2(new_n319), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n674), .A2(new_n319), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n657), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n319), .B(new_n674), .C1(new_n341), .C2(new_n347), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n807), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n877), .A2(new_n882), .ZN(new_n887));
  AOI221_X4 g0687(.A(new_n872), .B1(new_n851), .B2(new_n856), .C1(new_n445), .C2(new_n847), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n848), .B2(new_n857), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n886), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n446), .A2(new_n877), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n709), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n654), .A2(new_n652), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n846), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n880), .A2(new_n881), .ZN(new_n897));
  INV_X1    g0697(.A(new_n647), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n645), .A3(new_n643), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n809), .B1(new_n899), .B2(new_n639), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n655), .A2(new_n674), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n848), .A2(new_n857), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n872), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n858), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n896), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n878), .A2(new_n674), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT39), .B1(new_n871), .B2(new_n872), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n860), .A2(new_n910), .A3(new_n861), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT39), .B1(new_n888), .B2(new_n889), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n907), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n446), .B(new_n705), .C1(new_n706), .C2(new_n707), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(new_n661), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n914), .B(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n841), .B1(new_n894), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n917), .B2(new_n894), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n215), .A2(new_n225), .A3(new_n380), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n201), .B2(G68), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n921), .A2(new_n208), .A3(G13), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT103), .Z(new_n923));
  INV_X1    g0723(.A(KEYINPUT36), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n465), .B(new_n224), .C1(new_n519), .C2(KEYINPUT35), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(KEYINPUT35), .B2(new_n519), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n924), .B2(new_n926), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n919), .A2(new_n928), .ZN(G367));
  INV_X1    g0729(.A(new_n745), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n753), .B1(new_n212), .B2(new_n565), .C1(new_n930), .C2(new_n236), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n740), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n778), .A2(G317), .ZN(new_n933));
  INV_X1    g0733(.A(G311), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n933), .B1(new_n824), .B2(new_n934), .C1(new_n819), .C2(new_n770), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n759), .A2(new_n487), .B1(new_n790), .B2(new_n471), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n744), .ZN(new_n937));
  INV_X1    g0737(.A(new_n766), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(G97), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n831), .A2(KEYINPUT46), .A3(G116), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT46), .B1(new_n831), .B2(G116), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n513), .B2(new_n783), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n780), .A2(G143), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n267), .B1(new_n764), .B2(G50), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n758), .A2(G150), .B1(G58), .B2(new_n831), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n783), .A2(G68), .B1(new_n938), .B2(new_n264), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n944), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(G159), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n770), .A2(new_n949), .B1(new_n827), .B2(new_n777), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n935), .A2(new_n943), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT47), .Z(new_n952));
  NAND3_X1  g0752(.A1(new_n674), .A2(new_n633), .A3(new_n634), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n638), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n569), .B2(new_n953), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n932), .B1(new_n755), .B2(new_n952), .C1(new_n955), .C2(new_n798), .ZN(new_n956));
  INV_X1    g0756(.A(new_n681), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n734), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n958), .A2(new_n682), .A3(new_n684), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n684), .B1(new_n958), .B2(new_n682), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n702), .B(new_n536), .C1(new_n537), .C2(new_n688), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n640), .B1(new_n686), .B2(new_n687), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n685), .A2(new_n689), .A3(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT45), .Z(new_n966));
  NOR2_X1   g0766(.A1(new_n690), .A2(new_n964), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(KEYINPUT44), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT44), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n690), .A2(new_n969), .A3(new_n964), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n966), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n682), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n966), .B(new_n682), .C1(new_n968), .C2(new_n970), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n961), .A2(new_n973), .A3(new_n730), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n730), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n693), .B(KEYINPUT41), .Z(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n737), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT42), .ZN(new_n980));
  INV_X1    g0780(.A(new_n964), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(new_n685), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n964), .A2(KEYINPUT42), .A3(new_n681), .A4(new_n684), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n536), .B1(new_n962), .B2(new_n619), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n982), .A2(new_n983), .B1(new_n688), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n955), .B(KEYINPUT43), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT105), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT105), .B1(new_n985), .B2(new_n986), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n985), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n972), .A2(new_n964), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n995), .B1(KEYINPUT106), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(KEYINPUT106), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n956), .B1(new_n979), .B2(new_n999), .ZN(G387));
  AND2_X1   g0800(.A1(new_n961), .A2(new_n730), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1001), .A2(new_n694), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n730), .B2(new_n961), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n233), .A2(G45), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT107), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n361), .A2(new_n201), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT50), .ZN(new_n1007));
  AOI21_X1  g0807(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n695), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1005), .B(new_n745), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n742), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(G107), .B2(new_n212), .C1(new_n695), .C2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n741), .B1(new_n1012), .B2(new_n753), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n681), .B2(new_n798), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n762), .A2(new_n215), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n758), .B2(G50), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n309), .B2(new_n790), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n830), .B(new_n1017), .C1(G97), .C2(new_n938), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n359), .A2(new_n783), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n778), .A2(G150), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G159), .A2(new_n780), .B1(new_n769), .B2(new_n361), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n778), .A2(G326), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n744), .B1(G116), .B2(new_n938), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n782), .A2(new_n471), .B1(new_n762), .B2(new_n819), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G303), .A2(new_n764), .B1(new_n758), .B2(G317), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n824), .B2(new_n760), .C1(new_n934), .C2(new_n770), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT49), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1023), .B(new_n1024), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1022), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1014), .B1(new_n752), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n961), .B2(new_n737), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1003), .A2(new_n1036), .ZN(G393));
  NAND3_X1  g0837(.A1(new_n973), .A2(KEYINPUT108), .A3(new_n974), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT108), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n971), .A2(new_n1039), .A3(new_n972), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(KEYINPUT109), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT109), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1038), .A2(new_n1043), .A3(new_n1040), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n737), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n693), .B(new_n975), .C1(new_n1041), .C2(new_n1001), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n753), .B1(new_n522), .B2(new_n212), .C1(new_n930), .C2(new_n243), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n740), .A2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n780), .A2(G317), .B1(G311), .B2(new_n758), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT52), .Z(new_n1050));
  OAI22_X1  g0850(.A1(new_n782), .A2(new_n465), .B1(new_n766), .B2(new_n516), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n267), .B1(new_n471), .B2(new_n762), .C1(new_n790), .C2(new_n819), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G303), .C2(new_n769), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1050), .B(new_n1053), .C1(new_n760), .C2(new_n777), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT110), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n780), .A2(G150), .B1(G159), .B2(new_n758), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT51), .Z(new_n1058));
  NAND2_X1  g0858(.A1(new_n778), .A2(G143), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n769), .A2(G50), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n744), .B1(new_n309), .B2(new_n762), .C1(new_n790), .C2(new_n259), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n821), .B(new_n1061), .C1(G77), .C2(new_n783), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1056), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1048), .B1(new_n1065), .B2(new_n752), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n981), .A2(new_n751), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1045), .A2(new_n1046), .A3(new_n1068), .ZN(G390));
  INV_X1    g0869(.A(new_n897), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n901), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1070), .B1(new_n811), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n912), .B(new_n911), .C1(new_n1072), .C2(new_n908), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n672), .B(new_n808), .C1(new_n700), .C2(new_n704), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n1071), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n897), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n909), .A3(new_n874), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n709), .B1(new_n710), .B2(new_n876), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n882), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n729), .A2(new_n807), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n897), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1073), .A2(new_n1077), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n736), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n741), .B1(new_n259), .B2(new_n815), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n320), .B1(new_n759), .B2(new_n835), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G159), .B2(new_n783), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT54), .B(G143), .Z(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT111), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n831), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT53), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n762), .B2(new_n256), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1092), .A2(new_n764), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1090), .B(new_n1096), .C1(new_n201), .C2(new_n766), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n780), .A2(G128), .B1(new_n778), .B2(G125), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n827), .B2(new_n770), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(KEYINPUT112), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n320), .B1(new_n831), .B2(G87), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n759), .B2(new_n465), .C1(new_n522), .C2(new_n790), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n833), .B(new_n1103), .C1(G77), .C2(new_n783), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n769), .A2(new_n513), .B1(new_n778), .B2(G294), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(new_n471), .C2(new_n824), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(KEYINPUT112), .B2(new_n1100), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n911), .A2(new_n912), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1088), .B1(new_n755), .B2(new_n1108), .C1(new_n1109), .C2(new_n750), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT113), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1087), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1075), .B1(new_n897), .B2(new_n1083), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1079), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1070), .B1(new_n1114), .B2(new_n807), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1080), .B1(new_n1083), .B2(new_n897), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n811), .A2(new_n1071), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1113), .A2(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n446), .A2(new_n1079), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n915), .A2(new_n661), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1086), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n693), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1112), .A2(new_n1125), .ZN(G378));
  INV_X1    g0926(.A(new_n1120), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n709), .B1(new_n890), .B2(new_n884), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n874), .A2(new_n885), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT117), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n852), .A2(new_n298), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT116), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n378), .B1(new_n305), .B2(new_n306), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1133), .B(new_n378), .C1(new_n306), .C2(new_n305), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1131), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1141), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(KEYINPUT117), .A3(new_n1139), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1129), .A2(new_n1130), .A3(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n914), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1147), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n883), .B1(new_n904), .B2(new_n858), .ZN(new_n1151));
  OAI21_X1  g0951(.A(G330), .B1(new_n1151), .B2(KEYINPUT40), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1150), .B1(new_n886), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1109), .A2(new_n908), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1072), .A2(new_n905), .B1(new_n895), .B2(new_n846), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1129), .A2(new_n1145), .A3(new_n1130), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1153), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1149), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT57), .B1(new_n1128), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT118), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1124), .A2(new_n1127), .B1(new_n1149), .B2(new_n1158), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT118), .B1(new_n1163), .B2(KEYINPUT57), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1128), .A2(KEYINPUT57), .A3(new_n1159), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1162), .A2(new_n1164), .A3(new_n693), .A4(new_n1165), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n522), .A2(new_n770), .B1(new_n824), .B2(new_n465), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n777), .A2(new_n471), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n830), .B1(new_n202), .B2(new_n766), .C1(new_n309), .C2(new_n782), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G41), .B(new_n1015), .C1(G107), .C2(new_n758), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n565), .B2(new_n790), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G41), .B1(new_n744), .B2(G33), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1173), .A2(KEYINPUT58), .B1(G50), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(KEYINPUT58), .B2(new_n1173), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n780), .A2(G125), .B1(G150), .B2(new_n783), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT115), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1092), .A2(new_n831), .B1(G128), .B2(new_n758), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT114), .Z(new_n1180));
  AOI22_X1  g0980(.A1(new_n769), .A2(G132), .B1(G137), .B2(new_n764), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n778), .A2(G124), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n938), .C2(G159), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n755), .B1(new_n1176), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n739), .B1(G50), .B2(new_n816), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n1145), .C2(new_n749), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1159), .B2(new_n737), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1166), .A2(KEYINPUT119), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT119), .B1(new_n1166), .B2(new_n1191), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(G375));
  INV_X1    g0995(.A(new_n1118), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1070), .A2(new_n749), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n740), .B1(G68), .B2(new_n816), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n267), .B1(new_n759), .B2(new_n471), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n790), .A2(new_n351), .B1(new_n522), .B2(new_n762), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G77), .C2(new_n938), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n778), .A2(G303), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G116), .A2(new_n769), .B1(new_n780), .B2(G294), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1019), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n769), .A2(new_n1092), .B1(G137), .B2(new_n758), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n835), .B2(new_n824), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT120), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n778), .A2(G128), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n764), .A2(G150), .B1(G159), .B2(new_n831), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n783), .A2(G50), .B1(new_n938), .B2(G58), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1208), .A2(new_n744), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1204), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1198), .B1(new_n1212), .B2(new_n752), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1196), .A2(new_n737), .B1(new_n1197), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1122), .A2(new_n978), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1196), .A2(new_n1127), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(G381));
  AOI21_X1  g1017(.A(new_n736), .B1(new_n1041), .B2(KEYINPUT109), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1218), .A2(new_n1044), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n977), .B1(new_n975), .B2(new_n730), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n998), .B(new_n997), .C1(new_n1220), .C2(new_n737), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(new_n956), .A3(new_n1221), .A4(new_n1046), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1003), .A2(new_n800), .A3(new_n1036), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1223), .A2(G381), .A3(G384), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G378), .A2(G375), .A3(new_n1222), .A4(new_n1224), .ZN(G407));
  INV_X1    g1025(.A(G378), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(G343), .C2(new_n1227), .ZN(G409));
  NAND2_X1  g1028(.A1(G387), .A2(G390), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1222), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1231), .A2(new_n1223), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT61), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1223), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n1229), .A3(new_n1222), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT125), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1233), .A2(KEYINPUT125), .A3(new_n1234), .A4(new_n1236), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n667), .A2(G343), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1163), .A2(new_n978), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT121), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n736), .B1(new_n1159), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1149), .A2(new_n1158), .A3(KEYINPUT121), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1190), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT122), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1243), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI211_X1 g1049(.A(KEYINPUT122), .B(new_n1190), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1226), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n693), .B(new_n1165), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1163), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G378), .B(new_n1191), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1242), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1118), .A2(new_n1120), .A3(KEYINPUT60), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT123), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1256), .B(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT60), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1259), .A2(new_n1121), .A3(new_n694), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n814), .A2(KEYINPUT124), .A3(new_n839), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1261), .A2(new_n1214), .A3(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(G384), .B(KEYINPUT124), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1261), .B2(new_n1214), .ZN(new_n1265));
  INV_X1    g1065(.A(G2897), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1242), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n1263), .A2(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1261), .A2(new_n1214), .A3(new_n1262), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1267), .A2(new_n1266), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1261), .A2(new_n1214), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1269), .B(new_n1270), .C1(new_n1271), .C2(new_n1264), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1268), .A2(new_n1272), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1255), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1255), .A2(KEYINPUT63), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1255), .A2(new_n1275), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1241), .A2(new_n1274), .A3(new_n1276), .A4(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1234), .B1(new_n1255), .B2(new_n1273), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT126), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(new_n1234), .C1(new_n1255), .C2(new_n1273), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT62), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1277), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1255), .A2(KEYINPUT62), .A3(new_n1275), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1282), .A2(new_n1284), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1289));
  XOR2_X1   g1089(.A(new_n1289), .B(KEYINPUT127), .Z(new_n1290));
  OAI21_X1  g1090(.A(new_n1280), .B1(new_n1288), .B2(new_n1290), .ZN(G405));
  INV_X1    g1091(.A(new_n1289), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1166), .A2(new_n1191), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT119), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G378), .B1(new_n1295), .B2(new_n1192), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(G378), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1292), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1227), .A2(new_n1289), .A3(new_n1297), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1299), .A2(new_n1275), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1275), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(G402));
endmodule


