//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT88), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(new_n206), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n204), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n202), .B1(new_n210), .B2(KEYINPUT89), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n205), .B(new_n206), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(G1gat), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OAI221_X1 g013(.A(new_n210), .B1(KEYINPUT89), .B2(new_n202), .C1(G1gat), .C2(new_n212), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G29gat), .A2(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT15), .A4(new_n223), .ZN(new_n227));
  XNOR2_X1  g026(.A(G43gat), .B(G50gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n227), .A2(new_n228), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT87), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT87), .A2(KEYINPUT17), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n234), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n231), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT90), .B1(new_n216), .B2(new_n231), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n243));
  AOI211_X1 g042(.A(new_n243), .B(new_n232), .C1(new_n214), .C2(new_n215), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n240), .B(new_n241), .C1(new_n242), .C2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT92), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n249), .A3(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n217), .A2(new_n232), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(new_n242), .B2(new_n244), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n241), .B(KEYINPUT13), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G113gat), .B(G141gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G197gat), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT11), .B(G169gat), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT12), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n255), .B(new_n260), .C1(new_n246), .C2(new_n245), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n251), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n255), .B1(new_n246), .B2(new_n245), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT91), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n255), .B(new_n265), .C1(new_n246), .C2(new_n245), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n247), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n260), .B(KEYINPUT86), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G64gat), .B(G92gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  AND2_X1   g071(.A1(G226gat), .A2(G233gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(KEYINPUT23), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n278), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(G183gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(G190gat), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT24), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n283), .A2(new_n281), .A3(KEYINPUT24), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT64), .B(G169gat), .Z(new_n290));
  INV_X1    g089(.A(G176gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n274), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G183gat), .B(G190gat), .Z(new_n295));
  AOI21_X1  g094(.A(new_n286), .B1(new_n295), .B2(KEYINPUT24), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n278), .A2(G169gat), .A3(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(KEYINPUT25), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n296), .A2(KEYINPUT66), .A3(new_n280), .A4(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n280), .A2(new_n285), .A3(new_n299), .A4(new_n287), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n294), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT27), .B(G183gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(KEYINPUT28), .A3(new_n281), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT27), .B1(new_n308), .B2(new_n283), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT27), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n309), .A2(new_n310), .A3(new_n281), .A4(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n283), .A2(KEYINPUT27), .ZN(new_n316));
  AOI21_X1  g115(.A(G190gat), .B1(new_n316), .B2(KEYINPUT67), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n310), .B1(new_n317), .B2(new_n309), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n307), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n276), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(KEYINPUT26), .ZN(new_n321));
  INV_X1    g120(.A(new_n289), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(new_n320), .B2(KEYINPUT26), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n321), .A2(new_n323), .B1(G183gat), .B2(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n304), .A2(new_n305), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n305), .B1(new_n304), .B2(new_n325), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n273), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G211gat), .B(G218gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n332));
  OR2_X1    g131(.A1(G197gat), .A2(G204gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G197gat), .A2(G204gat), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n331), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n304), .A2(new_n325), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n273), .A2(KEYINPUT29), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n328), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(KEYINPUT73), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n304), .A2(new_n305), .A3(new_n325), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n304), .A2(new_n273), .A3(new_n325), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n337), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n272), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n345), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n336), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n328), .A2(new_n337), .A3(new_n340), .ZN(new_n350));
  INV_X1    g149(.A(new_n272), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(KEYINPUT74), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n347), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n349), .A2(new_n350), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT74), .B(KEYINPUT30), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n272), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT83), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361));
  INV_X1    g160(.A(G120gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G113gat), .ZN(new_n363));
  INV_X1    g162(.A(G113gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G120gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G127gat), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n369), .A2(KEYINPUT69), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(KEYINPUT69), .ZN(new_n371));
  OAI21_X1  g170(.A(G134gat), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G134gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n368), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT1), .B1(new_n363), .B2(new_n365), .ZN(new_n376));
  XNOR2_X1  g175(.A(G127gat), .B(G134gat), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(KEYINPUT70), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT70), .B1(new_n376), .B2(new_n377), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G141gat), .B(G148gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT2), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(G155gat), .B2(G162gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G141gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G148gat), .ZN(new_n389));
  INV_X1    g188(.A(G148gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G141gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G155gat), .B(G162gat), .ZN(new_n393));
  INV_X1    g192(.A(G155gat), .ZN(new_n394));
  INV_X1    g193(.A(G162gat), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT2), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n361), .B1(new_n380), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n387), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(KEYINPUT3), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n380), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n366), .A2(new_n377), .A3(new_n367), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT70), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n376), .A2(KEYINPUT70), .A3(new_n377), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n387), .A2(new_n397), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n409), .A2(new_n410), .A3(new_n375), .A4(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n399), .A2(new_n403), .A3(new_n404), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT5), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n404), .A2(KEYINPUT5), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n387), .A2(new_n397), .A3(new_n400), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n400), .B1(new_n387), .B2(new_n397), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n420), .B2(new_n380), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n366), .A2(new_n367), .B1(new_n369), .B2(new_n373), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n407), .A2(new_n408), .B1(new_n372), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n361), .A4(new_n410), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n409), .A2(new_n361), .A3(new_n410), .A4(new_n375), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT76), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n411), .B1(new_n423), .B2(new_n410), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n421), .B(new_n425), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT0), .ZN(new_n431));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n380), .A2(new_n398), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT77), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n409), .A2(new_n410), .A3(new_n375), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n404), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n380), .A2(KEYINPUT77), .A3(new_n398), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n416), .A2(new_n429), .A3(new_n433), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n360), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n441), .A2(new_n442), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n441), .A2(new_n442), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n416), .A2(new_n429), .A3(new_n440), .ZN(new_n446));
  INV_X1    g245(.A(new_n433), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n443), .B1(new_n449), .B2(new_n360), .ZN(new_n450));
  XNOR2_X1  g249(.A(G78gat), .B(G106gat), .ZN(new_n451));
  INV_X1    g250(.A(G50gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G22gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(KEYINPUT80), .A2(G22gat), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n400), .B1(new_n336), .B2(KEYINPUT29), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n398), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT79), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G228gat), .A2(G233gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n336), .B1(KEYINPUT29), .B2(new_n418), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n462), .A2(new_n463), .B1(G228gat), .B2(G233gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n468), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n460), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n466), .A2(new_n469), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n468), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n459), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT35), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n359), .A2(new_n450), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n338), .A2(new_n423), .ZN(new_n479));
  INV_X1    g278(.A(G227gat), .ZN(new_n480));
  INV_X1    g279(.A(G233gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n304), .A2(new_n380), .A3(new_n325), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT32), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(G71gat), .B(G99gat), .Z(new_n488));
  XNOR2_X1  g287(.A(G15gat), .B(G43gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n485), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(KEYINPUT33), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n484), .A2(KEYINPUT32), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n304), .A2(new_n380), .A3(new_n325), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n380), .B1(new_n304), .B2(new_n325), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n495), .A2(new_n496), .B1(new_n480), .B2(new_n481), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT34), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n499));
  OAI221_X1 g298(.A(new_n499), .B1(new_n480), .B2(new_n481), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n485), .A2(new_n487), .A3(new_n490), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n493), .A2(new_n498), .A3(new_n500), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT71), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n493), .A2(new_n498), .A3(new_n500), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT71), .B1(new_n507), .B2(new_n491), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n502), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT84), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n511), .B(new_n502), .C1(new_n506), .C2(new_n508), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n478), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n478), .A2(new_n510), .A3(KEYINPUT85), .A4(new_n512), .ZN(new_n516));
  INV_X1    g315(.A(new_n449), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n359), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n494), .A2(new_n501), .B1(new_n507), .B2(new_n491), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n473), .A2(new_n476), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT35), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n526));
  INV_X1    g325(.A(new_n509), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(KEYINPUT36), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n450), .B1(new_n356), .B2(new_n272), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n328), .A2(new_n336), .A3(new_n340), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT37), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT38), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n272), .B1(new_n356), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n356), .B2(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT38), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n529), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n399), .A2(new_n413), .A3(new_n403), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n438), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n437), .A2(new_n439), .ZN(new_n545));
  OAI211_X1 g344(.A(KEYINPUT39), .B(new_n544), .C1(new_n545), .C2(new_n438), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n544), .A2(KEYINPUT39), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT81), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n547), .A2(new_n548), .A3(new_n447), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n547), .B2(new_n447), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT40), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(KEYINPUT40), .B(new_n546), .C1(new_n549), .C2(new_n550), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n441), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n520), .B1(new_n555), .B2(new_n359), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n525), .B(new_n528), .C1(new_n542), .C2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n269), .B1(new_n523), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT98), .ZN(new_n559));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(G176gat), .B(G204gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(G57gat), .A2(G64gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G57gat), .A2(G64gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT93), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n577), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n571), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n582), .A2(KEYINPUT96), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n572), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n570), .B(new_n582), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n577), .A2(new_n580), .ZN(new_n587));
  INV_X1    g386(.A(new_n580), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n573), .B(new_n574), .C1(new_n578), .C2(KEYINPUT9), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n589), .B2(KEYINPUT93), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n584), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G230gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(new_n481), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT97), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n593), .A2(new_n598), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT10), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n592), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n595), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n563), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n600), .A2(new_n563), .A3(new_n604), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n559), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n607), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(KEYINPUT98), .A3(new_n605), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n572), .B1(new_n235), .B2(new_n238), .ZN(new_n612));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613));
  AND2_X1   g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(new_n232), .B2(new_n586), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n612), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n613), .B1(new_n612), .B2(new_n616), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT94), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AND4_X1   g421(.A1(KEYINPUT95), .A2(new_n617), .A3(new_n618), .A4(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n625), .A2(new_n622), .B1(new_n617), .B2(new_n618), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n587), .A2(new_n590), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n369), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n217), .B1(new_n630), .B2(new_n629), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G155gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n558), .A2(new_n611), .A3(new_n628), .A4(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n517), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(new_n203), .ZN(G1324gat));
  NOR2_X1   g445(.A1(new_n644), .A2(new_n359), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n202), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT16), .B(G8gat), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n644), .A2(new_n359), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT42), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(KEYINPUT42), .B2(new_n650), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n510), .A2(new_n512), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n644), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT99), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n644), .A2(new_n653), .A3(new_n528), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n644), .A2(new_n520), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  INV_X1    g460(.A(new_n643), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(new_n611), .A3(new_n627), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n558), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n218), .A3(new_n449), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT100), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n662), .A2(new_n611), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n269), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n628), .B1(new_n523), .B2(new_n557), .ZN(new_n674));
  AND2_X1   g473(.A1(KEYINPUT101), .A2(KEYINPUT44), .ZN(new_n675));
  NOR2_X1   g474(.A1(KEYINPUT101), .A2(KEYINPUT44), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AOI211_X1 g478(.A(new_n628), .B(new_n675), .C1(new_n523), .C2(new_n557), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n673), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G29gat), .B1(new_n683), .B2(new_n517), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n670), .A3(new_n684), .ZN(G1328gat));
  INV_X1    g484(.A(new_n359), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n665), .A2(new_n219), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT46), .Z(new_n688));
  OAI21_X1  g487(.A(G36gat), .B1(new_n683), .B2(new_n359), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1329gat));
  NOR2_X1   g489(.A1(new_n654), .A2(G43gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n558), .A2(new_n664), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT103), .Z(new_n693));
  INV_X1    g492(.A(new_n528), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n694), .B(new_n672), .C1(new_n678), .C2(new_n680), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G43gat), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT102), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1330gat));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n524), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G50gat), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n520), .A2(G50gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n665), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT104), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n665), .A2(new_n706), .A3(new_n703), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n705), .A2(KEYINPUT48), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n700), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n452), .B1(new_n682), .B2(new_n524), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n705), .A2(KEYINPUT48), .A3(new_n707), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT105), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n701), .A2(G50gat), .B1(new_n665), .B2(new_n703), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n709), .A2(new_n712), .B1(KEYINPUT48), .B2(new_n713), .ZN(G1331gat));
  NAND2_X1  g513(.A1(new_n267), .A2(new_n268), .ZN(new_n715));
  INV_X1    g514(.A(new_n262), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(new_n662), .A3(new_n627), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n608), .A2(new_n610), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT106), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n557), .B2(new_n523), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n449), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G57gat), .ZN(G1332gat));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n359), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT49), .B(G64gat), .Z(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(G1333gat));
  NAND2_X1  g529(.A1(new_n722), .A2(new_n694), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n654), .A2(G71gat), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n731), .A2(G71gat), .B1(new_n722), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1334gat));
  NAND2_X1  g534(.A1(new_n722), .A2(new_n524), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g536(.A1(new_n717), .A2(new_n611), .A3(new_n643), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n678), .B2(new_n680), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n517), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n523), .A2(new_n557), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n717), .A2(new_n643), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(new_n627), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n674), .A2(KEYINPUT51), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n719), .A2(new_n567), .A3(new_n449), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n740), .B1(new_n748), .B2(new_n749), .ZN(G1336gat));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751));
  INV_X1    g550(.A(new_n726), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(G92gat), .A3(new_n611), .ZN(new_n753));
  INV_X1    g552(.A(new_n746), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT51), .B1(new_n674), .B2(new_n742), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n747), .A2(KEYINPUT111), .A3(new_n753), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n726), .B(new_n738), .C1(new_n678), .C2(new_n680), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(G92gat), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n751), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT111), .B1(new_n747), .B2(new_n753), .ZN(new_n765));
  INV_X1    g564(.A(new_n753), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n757), .B(new_n766), .C1(new_n745), .C2(new_n746), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n763), .B(new_n751), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n745), .A2(new_n770), .A3(new_n746), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n755), .A2(KEYINPUT109), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n753), .A3(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n686), .B(new_n738), .C1(new_n678), .C2(new_n680), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT110), .B1(new_n776), .B2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n778), .B(new_n779), .C1(new_n773), .C2(new_n775), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n764), .A2(new_n769), .B1(new_n777), .B2(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n739), .B2(new_n528), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n654), .A2(G99gat), .A3(new_n611), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n748), .B2(new_n783), .ZN(G1338gat));
  NOR3_X1   g583(.A1(new_n611), .A2(new_n520), .A3(G106gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n771), .A2(new_n772), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G106gat), .B1(new_n739), .B2(new_n520), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n747), .A2(new_n785), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1339gat));
  NAND2_X1  g592(.A1(new_n718), .A2(new_n611), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n602), .A2(new_n595), .A3(new_n603), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n796), .A2(new_n604), .A3(new_n797), .ZN(new_n798));
  AOI211_X1 g597(.A(KEYINPUT54), .B(new_n595), .C1(new_n602), .C2(new_n603), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n800), .A3(new_n562), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n602), .A2(new_n603), .ZN(new_n802));
  INV_X1    g601(.A(new_n595), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT115), .B1(new_n804), .B2(new_n563), .ZN(new_n805));
  OAI211_X1 g604(.A(KEYINPUT55), .B(new_n798), .C1(new_n801), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n609), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n796), .A2(new_n604), .A3(new_n797), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n800), .B1(new_n799), .B2(new_n562), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n804), .A2(KEYINPUT115), .A3(new_n563), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(KEYINPUT55), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n795), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n607), .B1(new_n811), .B2(KEYINPUT55), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n798), .B1(new_n801), .B2(new_n805), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(KEYINPUT116), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n242), .A2(new_n244), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n241), .B1(new_n820), .B2(new_n240), .ZN(new_n821));
  INV_X1    g620(.A(new_n254), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n252), .B(new_n822), .C1(new_n242), .C2(new_n244), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n259), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n627), .B(new_n825), .C1(new_n251), .C2(new_n261), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n251), .B2(new_n261), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(new_n611), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n819), .B2(new_n269), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n827), .B1(new_n830), .B2(new_n628), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n794), .B1(new_n831), .B2(new_n643), .ZN(new_n832));
  AND4_X1   g631(.A1(new_n520), .A2(new_n832), .A3(new_n510), .A4(new_n512), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n726), .A2(new_n517), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(new_n364), .A3(new_n269), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n832), .A2(new_n449), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n837), .A2(new_n520), .A3(new_n519), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n752), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n717), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n836), .B1(new_n840), .B2(new_n364), .ZN(G1340gat));
  NOR3_X1   g640(.A1(new_n835), .A2(new_n362), .A3(new_n611), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n719), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n362), .ZN(G1341gat));
  NOR2_X1   g643(.A1(new_n370), .A2(new_n371), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n845), .A3(new_n643), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n835), .A2(new_n662), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n845), .B2(new_n847), .ZN(G1342gat));
  NAND2_X1  g647(.A1(new_n359), .A2(new_n627), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT117), .Z(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n838), .A2(new_n373), .A3(new_n851), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n835), .B2(new_n628), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G1343gat));
  NAND2_X1  g655(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n694), .A2(new_n520), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n837), .A2(new_n752), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n717), .A2(new_n388), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n811), .B2(KEYINPUT55), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n815), .A2(KEYINPUT119), .A3(new_n816), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n807), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n268), .ZN(new_n865));
  INV_X1    g664(.A(new_n247), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n263), .B2(KEYINPUT91), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n867), .B2(new_n266), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n864), .B1(new_n868), .B2(new_n262), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n627), .B1(new_n869), .B2(new_n829), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n662), .B1(new_n870), .B2(new_n827), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(KEYINPUT120), .B(new_n662), .C1(new_n870), .C2(new_n827), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n794), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n520), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n832), .A2(new_n524), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n875), .A2(new_n877), .B1(new_n878), .B2(new_n876), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n834), .A2(new_n528), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT118), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n879), .A2(new_n269), .A3(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G141gat), .ZN(new_n885));
  OAI221_X1 g684(.A(new_n857), .B1(new_n859), .B2(new_n860), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n859), .A2(new_n887), .A3(new_n860), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n879), .B2(new_n882), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n878), .A2(new_n876), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n794), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n819), .A2(new_n826), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n828), .A2(new_n611), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n717), .B2(new_n864), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n895), .B2(new_n627), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT120), .B1(new_n896), .B2(new_n662), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n877), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(KEYINPUT121), .A3(new_n881), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n890), .A2(new_n717), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n888), .B1(new_n901), .B2(G141gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n886), .B1(new_n902), .B2(new_n884), .ZN(G1344gat));
  INV_X1    g702(.A(new_n859), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n390), .A3(new_n719), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G148gat), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT121), .B1(new_n899), .B2(new_n881), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n889), .B(new_n882), .C1(new_n891), .C2(new_n898), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(new_n910), .B2(new_n719), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n832), .A2(new_n877), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n814), .A2(new_n627), .A3(new_n817), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(KEYINPUT124), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(KEYINPUT124), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n915), .A2(new_n916), .A3(new_n828), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n662), .B1(new_n870), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n520), .B1(new_n918), .B2(new_n794), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n912), .A2(new_n913), .B1(new_n919), .B2(KEYINPUT57), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n912), .A2(new_n913), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n719), .B(new_n881), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n906), .B1(new_n922), .B2(G148gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n905), .B1(new_n911), .B2(new_n923), .ZN(G1345gat));
  AOI21_X1  g723(.A(G155gat), .B1(new_n904), .B2(new_n643), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n643), .A2(G155gat), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT125), .Z(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n910), .B2(new_n927), .ZN(G1346gat));
  NOR3_X1   g727(.A1(new_n908), .A2(new_n909), .A3(new_n628), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n837), .A2(new_n858), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n851), .A2(new_n395), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n929), .A2(new_n395), .B1(new_n930), .B2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n359), .A2(new_n449), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n833), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n269), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n832), .A2(new_n517), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n752), .A2(new_n521), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n269), .A2(new_n290), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  OAI21_X1  g739(.A(G176gat), .B1(new_n934), .B2(new_n611), .ZN(new_n941));
  INV_X1    g740(.A(new_n938), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n291), .A3(new_n719), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1349gat));
  OAI21_X1  g743(.A(G183gat), .B1(new_n934), .B2(new_n662), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n942), .A2(new_n306), .A3(new_n643), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n947), .B(new_n948), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n942), .A2(new_n281), .A3(new_n627), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n281), .B1(new_n951), .B2(KEYINPUT61), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n952), .B1(new_n934), .B2(new_n628), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n951), .A2(KEYINPUT61), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(G1351gat));
  NOR3_X1   g756(.A1(new_n694), .A2(new_n752), .A3(new_n520), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n936), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n717), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n920), .A2(new_n921), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n528), .A2(new_n933), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n717), .A2(G197gat), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(G1352gat));
  OAI21_X1  g766(.A(G204gat), .B1(new_n964), .B2(new_n611), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n959), .A2(G204gat), .A3(new_n611), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(G1353gat));
  OR3_X1    g770(.A1(new_n959), .A2(G211gat), .A3(new_n662), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n643), .B(new_n963), .C1(new_n920), .C2(new_n921), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  OAI21_X1  g775(.A(G218gat), .B1(new_n964), .B2(new_n628), .ZN(new_n977));
  OR3_X1    g776(.A1(new_n959), .A2(G218gat), .A3(new_n628), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1355gat));
endmodule


