//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G116), .A2(G270), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G107), .A2(G264), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G68), .A2(G238), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR3_X1   g0016(.A1(new_n210), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G58), .A2(G232), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n205), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT1), .Z(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  INV_X1    g0021(.A(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n205), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n221), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G68), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n231), .A2(new_n204), .A3(new_n232), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n220), .A2(new_n227), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n232), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT67), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n229), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n255), .B1(new_n258), .B2(new_n214), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT11), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n203), .A2(G20), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n222), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n229), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT12), .ZN(new_n265));
  INV_X1    g0065(.A(new_n251), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G68), .A3(new_n262), .ZN(new_n267));
  XOR2_X1   g0067(.A(new_n267), .B(KEYINPUT74), .Z(new_n268));
  AND3_X1   g0068(.A1(new_n261), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n232), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n212), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n275), .B(new_n277), .C1(G232), .C2(new_n276), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G97), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n272), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT64), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n271), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(KEYINPUT64), .A2(G33), .A3(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n270), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n281), .ZN(new_n289));
  INV_X1    g0089(.A(G238), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n284), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n280), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT13), .B1(new_n280), .B2(new_n291), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G169), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT14), .ZN(new_n298));
  INV_X1    g0098(.A(new_n296), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G179), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT14), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n296), .A2(new_n301), .A3(G169), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT75), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT75), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n298), .A2(new_n300), .A3(new_n305), .A4(new_n302), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n269), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n296), .A2(G200), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n299), .A2(G190), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n269), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g0111(.A(KEYINPUT8), .B(G58), .Z(new_n312));
  INV_X1    g0112(.A(KEYINPUT68), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT68), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(new_n257), .B1(G150), .B2(new_n254), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT69), .ZN(new_n319));
  OAI21_X1  g0119(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n253), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n263), .A2(new_n211), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n252), .A2(new_n262), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G50), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n275), .A2(new_n214), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n276), .A2(G222), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT65), .B(G223), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n276), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n327), .B1(new_n330), .B2(new_n275), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT66), .ZN(new_n332));
  INV_X1    g0132(.A(new_n272), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n289), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n283), .B1(new_n335), .B2(G226), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(new_n340), .A3(new_n336), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n326), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n254), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n344), .A2(KEYINPUT70), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(KEYINPUT70), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n312), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT15), .B(G87), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n349), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n347), .B1(new_n204), .B2(new_n214), .C1(new_n352), .C2(new_n258), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n251), .B1(new_n214), .B2(new_n263), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n266), .A2(G77), .A3(new_n262), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n276), .A2(G232), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n275), .B(new_n357), .C1(new_n290), .C2(new_n276), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n333), .C1(G107), .C2(new_n275), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n284), .C1(new_n215), .C2(new_n289), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n338), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(G179), .B2(new_n360), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(G200), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n356), .B(new_n364), .C1(new_n365), .C2(new_n360), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n337), .A2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n334), .A2(G190), .A3(new_n336), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n368), .B(new_n372), .C1(new_n373), .C2(KEYINPUT9), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT9), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n326), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n371), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n371), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(KEYINPUT9), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n326), .A2(new_n375), .B1(G200), .B2(new_n337), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n372), .ZN(new_n381));
  AOI211_X1 g0181(.A(new_n343), .B(new_n367), .C1(new_n377), .C2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT73), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n311), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n377), .A2(new_n381), .ZN(new_n385));
  INV_X1    g0185(.A(new_n367), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n385), .A2(new_n383), .A3(new_n342), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n212), .A2(G1698), .ZN(new_n388));
  AND2_X1   g0188(.A1(KEYINPUT3), .A2(G33), .ZN(new_n389));
  NOR2_X1   g0189(.A1(KEYINPUT3), .A2(G33), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n388), .B1(G223), .B2(G1698), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n333), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n288), .A2(G232), .A3(new_n281), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n394), .A2(G179), .A3(new_n284), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n284), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n272), .B1(new_n391), .B2(new_n392), .ZN(new_n398));
  OAI21_X1  g0198(.A(G169), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n389), .A2(new_n390), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n402), .B2(new_n204), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  NOR4_X1   g0204(.A1(new_n389), .A2(new_n390), .A3(new_n404), .A4(G20), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n254), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G58), .A2(G68), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n230), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n406), .A2(KEYINPUT16), .A3(new_n407), .A4(new_n410), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n251), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n263), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n317), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n324), .B2(new_n317), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(KEYINPUT76), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT76), .B1(new_n415), .B2(new_n418), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n401), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT18), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n394), .A2(new_n284), .A3(new_n395), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT77), .B(G190), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(G200), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n415), .A2(new_n426), .A3(new_n427), .A4(new_n418), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT17), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n401), .C1(new_n420), .C2(new_n421), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n423), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n387), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n384), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n263), .B1(new_n203), .B2(G33), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n252), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n437), .A2(G107), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT23), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n204), .B2(G107), .ZN(new_n442));
  INV_X1    g0242(.A(G107), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(KEYINPUT23), .A3(G20), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G116), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G20), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n204), .B(G87), .C1(new_n389), .C2(new_n390), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT22), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT22), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n275), .A2(new_n450), .A3(new_n204), .A4(G87), .ZN(new_n451));
  AOI211_X1 g0251(.A(new_n445), .B(new_n447), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n440), .B1(new_n452), .B2(KEYINPUT86), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n447), .B1(new_n449), .B2(new_n451), .ZN(new_n454));
  INV_X1    g0254(.A(new_n445), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT86), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(new_n439), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n452), .A2(KEYINPUT86), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n453), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n438), .B1(new_n460), .B2(new_n251), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n443), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT87), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT25), .B1(new_n263), .B2(new_n443), .ZN(new_n464));
  XOR2_X1   g0264(.A(new_n463), .B(new_n464), .Z(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n288), .A2(new_n471), .A3(G264), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT88), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT88), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n288), .A2(new_n471), .A3(new_n474), .A4(G264), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n224), .A2(G1698), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n275), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G250), .A2(G1698), .ZN(new_n479));
  INV_X1    g0279(.A(G294), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n478), .A2(new_n479), .B1(new_n256), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n333), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n468), .B(G274), .C1(new_n470), .C2(new_n469), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n476), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT89), .B1(new_n484), .B2(G169), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n484), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G179), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n484), .A2(KEYINPUT89), .A3(G169), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n466), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(G33), .B2(G283), .ZN(new_n492));
  INV_X1    g0292(.A(G97), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(G33), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n495), .A2(KEYINPUT20), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G20), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n494), .A2(new_n496), .A3(new_n251), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(KEYINPUT20), .ZN(new_n500));
  XNOR2_X1  g0300(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n251), .A2(new_n497), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n436), .A2(new_n502), .B1(new_n497), .B2(new_n263), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n276), .A2(G257), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n275), .B(new_n505), .C1(new_n225), .C2(new_n276), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n506), .B(new_n333), .C1(G303), .C2(new_n275), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n288), .A2(new_n471), .A3(G270), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n483), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(G169), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT21), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n501), .A2(new_n503), .ZN(new_n514));
  OR3_X1    g0314(.A1(new_n514), .A2(new_n340), .A3(new_n509), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n473), .A2(new_n475), .B1(new_n481), .B2(new_n333), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n365), .A3(new_n483), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(KEYINPUT90), .C1(new_n487), .C2(G200), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n518), .A2(KEYINPUT90), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n461), .A2(new_n519), .A3(new_n465), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n509), .A2(G200), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n514), .B(new_n522), .C1(new_n425), .C2(new_n509), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n491), .A2(new_n516), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n215), .A2(G1698), .ZN(new_n525));
  OAI221_X1 g0325(.A(new_n525), .B1(G238), .B2(G1698), .C1(new_n389), .C2(new_n390), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n272), .B1(new_n526), .B2(new_n446), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n221), .B1(new_n467), .B2(G1), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n468), .A2(new_n282), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n288), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT83), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT83), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n288), .A2(new_n532), .A3(new_n528), .A4(new_n529), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n527), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G179), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n338), .B2(new_n534), .ZN(new_n536));
  INV_X1    g0336(.A(new_n352), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n437), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n352), .A2(new_n263), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n275), .A2(new_n204), .A3(G68), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  INV_X1    g0341(.A(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n279), .A2(new_n204), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(KEYINPUT19), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n279), .A2(G20), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n540), .B(new_n545), .C1(KEYINPUT19), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n251), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n538), .A2(new_n539), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n536), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n534), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n252), .A2(G87), .A3(new_n436), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n539), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n534), .A2(G190), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n416), .A2(G97), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n252), .A2(G97), .A3(new_n436), .ZN(new_n560));
  OAI21_X1  g0360(.A(G107), .B1(new_n403), .B2(new_n405), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT6), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n493), .A2(new_n443), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(new_n541), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n443), .A2(KEYINPUT6), .A3(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G20), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n561), .B(new_n567), .C1(new_n214), .C2(new_n344), .ZN(new_n568));
  AOI211_X1 g0368(.A(new_n559), .B(new_n560), .C1(new_n568), .C2(new_n251), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(new_n276), .C1(new_n389), .C2(new_n390), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT78), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n571), .A2(KEYINPUT4), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n275), .A2(G244), .A3(new_n276), .A4(new_n572), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n275), .A2(G250), .A3(G1698), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n571), .A2(KEYINPUT4), .B1(G33), .B2(G283), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n333), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n288), .A2(new_n471), .A3(G257), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT79), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n483), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n583), .B1(new_n582), .B2(new_n483), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT80), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(new_n483), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT79), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT80), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n590), .A3(new_n584), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n581), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G200), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n569), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n580), .A2(new_n589), .A3(G190), .A4(new_n584), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT81), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n585), .A2(new_n586), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(KEYINPUT81), .A3(G190), .A4(new_n580), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT82), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n597), .A2(new_n599), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT80), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n590), .B1(new_n589), .B2(new_n584), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n580), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G200), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT82), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n602), .A2(new_n606), .A3(new_n607), .A4(new_n569), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n560), .B1(new_n568), .B2(new_n251), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G97), .B2(new_n416), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n598), .A2(new_n580), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n338), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n612), .C1(G179), .C2(new_n605), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n601), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n524), .A2(new_n558), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n435), .A2(new_n615), .ZN(G372));
  NAND2_X1  g0416(.A1(new_n415), .A2(new_n418), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT95), .B1(new_n617), .B2(new_n401), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(KEYINPUT95), .A3(new_n401), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n430), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT95), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n622), .B(new_n400), .C1(new_n415), .C2(new_n418), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT18), .B1(new_n623), .B2(new_n618), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n363), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n310), .A2(new_n308), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n307), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n429), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n343), .B1(new_n630), .B2(new_n385), .ZN(new_n631));
  INV_X1    g0431(.A(new_n435), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n601), .A2(new_n608), .A3(new_n613), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT92), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT91), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n534), .A2(new_n338), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n340), .B(new_n527), .C1(new_n531), .C2(new_n533), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n535), .B(KEYINPUT91), .C1(new_n338), .C2(new_n534), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n635), .B1(new_n641), .B2(new_n549), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n521), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n633), .A2(new_n634), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n491), .A2(new_n516), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n521), .A2(new_n642), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT92), .B1(new_n614), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n569), .B1(new_n340), .B2(new_n592), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n554), .B1(new_n551), .B2(G200), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n650), .A2(new_n556), .B1(new_n536), .B2(new_n549), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n649), .A2(new_n651), .A3(KEYINPUT26), .A4(new_n612), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n641), .A2(KEYINPUT93), .A3(new_n549), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT93), .B1(new_n641), .B2(new_n549), .ZN(new_n654));
  OAI22_X1  g0454(.A1(new_n652), .A2(KEYINPUT94), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n613), .A2(new_n558), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n613), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n642), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n655), .B1(new_n660), .B2(KEYINPUT94), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n648), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n631), .B1(new_n632), .B2(new_n663), .ZN(G369));
  NAND2_X1  g0464(.A1(new_n491), .A2(new_n521), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n222), .A2(G20), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n203), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n665), .B1(new_n466), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n489), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n485), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n488), .A2(new_n675), .B1(new_n461), .B2(new_n465), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n673), .B1(new_n676), .B2(new_n672), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n516), .B2(new_n672), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n516), .A2(new_n523), .ZN(new_n679));
  INV_X1    g0479(.A(new_n672), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n514), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g0481(.A(new_n679), .B(new_n516), .S(new_n681), .Z(new_n682));
  INV_X1    g0482(.A(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n665), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n516), .A2(new_n672), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n676), .A2(new_n680), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(G399));
  OR2_X1    g0493(.A1(new_n223), .A2(G41), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G1), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n541), .A2(new_n542), .A3(new_n497), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n695), .A2(new_n696), .B1(new_n231), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n611), .A2(new_n509), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n517), .A3(new_n638), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT96), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n700), .B(new_n702), .Z(new_n703));
  NOR3_X1   g0503(.A1(new_n592), .A2(new_n487), .A3(new_n534), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n704), .A2(new_n340), .A3(new_n509), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n672), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(KEYINPUT31), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n615), .B2(new_n680), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n707), .B1(new_n709), .B2(new_n706), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n683), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n672), .B1(new_n648), .B2(new_n661), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT97), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(KEYINPUT97), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT98), .B1(new_n676), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT98), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n491), .A2(new_n720), .A3(new_n516), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n719), .A2(new_n633), .A3(new_n721), .A4(new_n643), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n656), .B1(new_n658), .B2(new_n642), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n653), .A2(new_n654), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n613), .A2(new_n558), .A3(KEYINPUT26), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n672), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT29), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n712), .B1(new_n717), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n698), .B1(new_n729), .B2(G1), .ZN(G364));
  INV_X1    g0530(.A(new_n684), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n695), .B1(G45), .B2(new_n666), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n682), .A2(new_n683), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(G20), .B1(KEYINPUT100), .B2(G169), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(KEYINPUT100), .A2(G169), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n232), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n204), .A2(new_n340), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n593), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n275), .B1(new_n744), .B2(new_n214), .C1(new_n229), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n204), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G159), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  OR3_X1    g0554(.A1(new_n593), .A2(KEYINPUT101), .A3(G179), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT101), .B1(new_n593), .B2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n757), .A2(new_n204), .A3(new_n365), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n754), .B1(G87), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n757), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n749), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n759), .B1(new_n443), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n745), .A2(new_n425), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n748), .B(new_n762), .C1(G50), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n742), .A2(new_n425), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n750), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n764), .B1(new_n228), .B2(new_n766), .C1(new_n493), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n758), .ZN(new_n771));
  INV_X1    g0571(.A(G303), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n771), .A2(new_n772), .B1(new_n761), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n275), .B1(new_n765), .B2(G322), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n752), .A2(G329), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n775), .B(new_n776), .C1(new_n480), .C2(new_n769), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n774), .B(new_n777), .C1(new_n746), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  INV_X1    g0580(.A(G326), .ZN(new_n781));
  INV_X1    g0581(.A(new_n763), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n779), .B1(new_n780), .B2(new_n744), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n740), .B1(new_n770), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n682), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n223), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n275), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT99), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G355), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n223), .A2(new_n275), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n231), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(new_n467), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n245), .B2(new_n467), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n792), .B(new_n797), .C1(G116), .C2(new_n789), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n739), .A2(new_n787), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n788), .A2(new_n800), .A3(new_n732), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n735), .B1(new_n784), .B2(new_n801), .ZN(G396));
  OR2_X1    g0602(.A1(new_n356), .A2(new_n680), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n386), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(KEYINPUT102), .B1(new_n803), .B2(new_n362), .ZN(new_n805));
  OR3_X1    g0605(.A1(new_n803), .A2(KEYINPUT102), .A3(new_n362), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n662), .A2(new_n680), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n714), .A2(new_n716), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(new_n807), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n712), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n808), .B1(new_n683), .B2(new_n711), .C1(new_n809), .C2(new_n807), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n811), .A2(new_n812), .A3(new_n733), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT103), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n402), .B1(new_n751), .B2(new_n780), .C1(new_n769), .C2(new_n493), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n743), .A2(G116), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n816), .B1(new_n761), .B2(new_n542), .C1(new_n771), .C2(new_n443), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(G294), .C2(new_n765), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n818), .B1(new_n773), .B2(new_n747), .C1(new_n772), .C2(new_n782), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G143), .A2(new_n765), .B1(new_n743), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n782), .C1(new_n822), .C2(new_n747), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n761), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n823), .A2(new_n824), .B1(G68), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n768), .A2(G58), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n402), .B1(new_n752), .B2(G132), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n825), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n771), .A2(new_n211), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n819), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n739), .A2(new_n785), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n832), .A2(new_n739), .B1(new_n214), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n807), .B2(new_n786), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n732), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n813), .A2(new_n814), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n814), .B1(new_n813), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(G384));
  OAI211_X1 g0639(.A(G20), .B(new_n270), .C1(new_n566), .C2(KEYINPUT35), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n497), .B(new_n840), .C1(KEYINPUT35), .C2(new_n566), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT36), .Z(new_n842));
  NAND3_X1  g0642(.A1(new_n795), .A2(G77), .A3(new_n408), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT104), .Z(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(G50), .B2(new_n229), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(G1), .A3(new_n222), .ZN(new_n846));
  XNOR2_X1  g0646(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n847));
  INV_X1    g0647(.A(new_n670), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n413), .A2(new_n253), .A3(new_n414), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n418), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n432), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n421), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n419), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n400), .A2(new_n670), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n428), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n850), .A2(new_n854), .ZN(new_n857));
  INV_X1    g0657(.A(new_n428), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT37), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n851), .A2(KEYINPUT38), .A3(new_n860), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n524), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n867), .A2(new_n651), .A3(new_n633), .A4(new_n680), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n706), .A2(KEYINPUT31), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n304), .A2(new_n306), .ZN(new_n871));
  INV_X1    g0671(.A(new_n269), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n672), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n627), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n307), .A2(new_n672), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n869), .A2(new_n870), .A3(new_n877), .A4(new_n807), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n847), .B1(new_n866), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n848), .B1(new_n420), .B2(new_n421), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n625), .B2(new_n429), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(new_n619), .A3(new_n428), .A4(new_n620), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .B1(new_n855), .B2(new_n428), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n862), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n864), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT106), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT40), .B(new_n885), .C1(new_n878), .C2(new_n886), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n878), .A2(new_n886), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n879), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n435), .A2(new_n710), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n889), .B(new_n890), .Z(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(G330), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT107), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n435), .A2(new_n717), .A3(new_n728), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n631), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n875), .A2(new_n876), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n363), .A2(new_n672), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n808), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n865), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n621), .A2(new_n624), .A3(new_n670), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n885), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n863), .A2(KEYINPUT39), .A3(new_n864), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n307), .A2(new_n680), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n901), .A2(new_n902), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n896), .B(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n666), .A2(new_n203), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n842), .B(new_n846), .C1(new_n911), .C2(new_n912), .ZN(G367));
  NAND2_X1  g0713(.A1(new_n554), .A2(new_n672), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n653), .A2(new_n654), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n642), .B2(new_n914), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT43), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n633), .B1(new_n569), .B2(new_n680), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n613), .A2(new_n680), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT108), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT109), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n613), .B1(new_n924), .B2(new_n491), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n680), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n922), .A2(new_n690), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT42), .Z(new_n928));
  AOI21_X1  g0728(.A(new_n918), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n916), .A2(new_n917), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n926), .A2(new_n917), .A3(new_n916), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n685), .B2(new_n924), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n685), .A2(new_n924), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n203), .B1(new_n666), .B2(G45), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n694), .B(KEYINPUT41), .Z(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n678), .A2(new_n684), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n691), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n689), .A2(new_n692), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(new_n922), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT44), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n922), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT45), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n942), .A2(new_n948), .A3(new_n729), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n940), .B1(new_n949), .B2(new_n729), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n934), .B(new_n936), .C1(new_n938), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n241), .A2(new_n793), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n952), .B(new_n799), .C1(new_n789), .C2(new_n352), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT110), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n826), .A2(G97), .ZN(new_n955));
  INV_X1    g0755(.A(G317), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n955), .B(new_n402), .C1(new_n956), .C2(new_n751), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT112), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(G283), .B2(new_n743), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT111), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n771), .B2(new_n497), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT46), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n765), .A2(G303), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n746), .A2(G294), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n780), .B2(new_n782), .C1(new_n961), .C2(KEYINPUT46), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G107), .B2(new_n768), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n959), .A2(new_n962), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n275), .B1(new_n821), .B2(new_n751), .C1(new_n766), .C2(new_n822), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n826), .A2(G77), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n763), .A2(G143), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(new_n228), .C2(new_n771), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n968), .B(new_n971), .C1(G50), .C2(new_n743), .ZN(new_n972));
  INV_X1    g0772(.A(G159), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n972), .B1(new_n229), .B2(new_n769), .C1(new_n973), .C2(new_n747), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n967), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n733), .B(new_n954), .C1(new_n976), .C2(new_n739), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT113), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n916), .A2(new_n787), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n951), .A2(new_n980), .ZN(G387));
  NAND2_X1  g0781(.A1(new_n942), .A2(new_n938), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n402), .B1(new_n317), .B2(new_n746), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n955), .B(new_n983), .C1(new_n211), .C2(new_n766), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n537), .A2(new_n768), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n752), .A2(G150), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n763), .A2(KEYINPUT114), .A3(G159), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT114), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n782), .B2(new_n973), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n771), .A2(new_n214), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n744), .A2(new_n229), .ZN(new_n992));
  NOR4_X1   g0792(.A1(new_n984), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT115), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G311), .A2(new_n746), .B1(new_n763), .B2(G322), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n772), .B2(new_n744), .C1(new_n956), .C2(new_n766), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT116), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT48), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n773), .B2(new_n769), .C1(new_n480), .C2(new_n771), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT49), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n402), .B1(new_n781), .B2(new_n751), .C1(new_n761), .C2(new_n497), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n994), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n739), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n238), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n793), .B1(new_n1004), .B2(new_n467), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n791), .A2(new_n696), .ZN(new_n1006));
  AOI211_X1 g0806(.A(G45), .B(new_n696), .C1(G68), .C2(G77), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n315), .A2(G50), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1005), .A2(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n789), .A2(G107), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n799), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n677), .A2(new_n787), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1003), .A2(new_n732), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n942), .A2(new_n729), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n694), .B(KEYINPUT117), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n942), .A2(new_n729), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n982), .B(new_n1014), .C1(new_n1017), .C2(new_n1018), .ZN(G393));
  NAND2_X1  g0819(.A1(new_n948), .A2(new_n686), .ZN(new_n1020));
  OR3_X1    g0820(.A1(new_n945), .A2(new_n686), .A3(new_n947), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n938), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n733), .B1(new_n924), .B2(new_n787), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n799), .B1(new_n493), .B2(new_n789), .C1(new_n248), .C2(new_n794), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G311), .A2(new_n765), .B1(new_n763), .B2(G317), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT52), .Z(new_n1026));
  AOI21_X1  g0826(.A(new_n275), .B1(new_n752), .B2(G322), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n443), .C2(new_n761), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n747), .A2(new_n772), .B1(new_n744), .B2(new_n480), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G116), .B2(new_n768), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT118), .Z(new_n1031));
  AOI211_X1 g0831(.A(new_n1028), .B(new_n1031), .C1(G283), .C2(new_n758), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G150), .A2(new_n763), .B1(new_n765), .B2(G159), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT51), .Z(new_n1034));
  AOI22_X1  g0834(.A1(new_n743), .A2(new_n312), .B1(G143), .B2(new_n752), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n211), .C2(new_n747), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n771), .A2(new_n229), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n769), .A2(new_n214), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n275), .B1(new_n761), .B2(new_n542), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n739), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1023), .A2(new_n1024), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1022), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT119), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1022), .A2(KEYINPUT119), .A3(new_n1042), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n1015), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n949), .A3(new_n1016), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1050), .ZN(G390));
  INV_X1    g0851(.A(KEYINPUT120), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n904), .A2(new_n905), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n900), .B2(new_n907), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n722), .A2(new_n726), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n680), .A3(new_n807), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n897), .B1(new_n1056), .B2(new_n899), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n885), .A2(new_n906), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n710), .A2(G330), .A3(new_n807), .A4(new_n877), .ZN(new_n1061));
  AND4_X1   g0861(.A1(new_n1052), .A2(new_n1054), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n898), .B1(new_n713), .B2(new_n807), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n906), .B1(new_n1063), .B2(new_n897), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1059), .B1(new_n1064), .B2(new_n1053), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n1052), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1061), .B1(new_n1065), .B2(new_n1052), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1062), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n869), .A2(G330), .A3(new_n870), .A4(new_n807), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n897), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n898), .B1(new_n727), .B2(new_n807), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1061), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT121), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT121), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1061), .A2(new_n1070), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1063), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1073), .B1(new_n1077), .B2(new_n1072), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n435), .A2(G330), .A3(new_n710), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n894), .A2(new_n1079), .A3(new_n631), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1068), .B1(new_n1082), .B2(KEYINPUT122), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1065), .A2(new_n1052), .A3(new_n1061), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1061), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(KEYINPUT120), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(KEYINPUT120), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT122), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n1090), .A3(new_n1081), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1083), .A2(new_n1016), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n786), .B1(new_n904), .B2(new_n905), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n833), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(new_n317), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n771), .A2(new_n822), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT53), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1096), .A2(new_n1097), .B1(new_n744), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1097), .B2(new_n1096), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G132), .A2(new_n765), .B1(new_n746), .B2(G137), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1101), .B(new_n275), .C1(new_n973), .C2(new_n769), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G50), .B2(new_n826), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G125), .B2(new_n752), .ZN(new_n1105));
  INV_X1    g0905(.A(G128), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n782), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n771), .A2(new_n542), .B1(new_n761), .B2(new_n229), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n493), .A2(new_n744), .B1(new_n782), .B2(new_n773), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n402), .B1(new_n751), .B2(new_n480), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n1108), .A2(new_n1038), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n443), .B2(new_n747), .C1(new_n497), .C2(new_n766), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n740), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  NOR4_X1   g0913(.A1(new_n1093), .A2(new_n733), .A3(new_n1095), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1068), .B2(new_n938), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1092), .A2(new_n1115), .ZN(G378));
  INV_X1    g0916(.A(KEYINPUT57), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n894), .A2(new_n1079), .A3(new_n631), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1068), .B2(new_n1078), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n385), .A2(new_n342), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n385), .B2(new_n342), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1123), .A2(new_n1124), .B1(new_n373), .B2(new_n670), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1124), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n373), .A2(new_n670), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n1122), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n889), .B2(new_n683), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n878), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT106), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n878), .A2(new_n886), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1133), .A2(KEYINPUT40), .A3(new_n885), .A4(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1135), .A2(G330), .A3(new_n879), .A4(new_n1129), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n909), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1131), .A2(new_n1136), .A3(new_n910), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1117), .B1(new_n1119), .B2(new_n1140), .ZN(new_n1141));
  AND4_X1   g0941(.A1(KEYINPUT121), .A2(new_n1061), .A3(new_n1071), .A4(new_n1070), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1132), .A2(G330), .B1(new_n1069), .B2(new_n897), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT121), .B1(new_n1143), .B2(new_n1063), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1072), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1080), .B1(new_n1089), .B2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1131), .A2(new_n1136), .A3(new_n910), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n910), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1150), .A3(KEYINPUT57), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1141), .A2(new_n1016), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n211), .B1(new_n389), .B2(G41), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n402), .B1(new_n751), .B2(new_n773), .C1(new_n769), .C2(new_n229), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1154), .B(new_n991), .C1(G97), .C2(new_n746), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n761), .A2(new_n228), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n352), .A2(new_n744), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n766), .A2(new_n443), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(G41), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1155), .B(new_n1159), .C1(new_n497), .C2(new_n782), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT58), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n763), .A2(G125), .B1(G150), .B2(new_n768), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT123), .Z(new_n1163));
  INV_X1    g0963(.A(G132), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n747), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G137), .B2(new_n743), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n1106), .B2(new_n766), .C1(new_n771), .C2(new_n1098), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(new_n1167), .B2(KEYINPUT59), .ZN(new_n1168));
  AOI21_X1  g0968(.A(G33), .B1(new_n752), .B2(G124), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n973), .C2(new_n761), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1167), .A2(KEYINPUT59), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1153), .B(new_n1161), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n733), .B1(new_n1172), .B2(new_n739), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(G50), .B2(new_n1094), .C1(new_n1130), .C2(new_n786), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1150), .B2(new_n938), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1152), .A2(new_n1176), .ZN(G375));
  INV_X1    g0977(.A(KEYINPUT124), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1146), .A2(KEYINPUT124), .A3(new_n1118), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n939), .A3(new_n1081), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n937), .B(KEYINPUT125), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1078), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n897), .A2(new_n785), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n833), .A2(new_n229), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1156), .B1(G50), .B2(new_n768), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n1164), .B2(new_n782), .C1(new_n747), .C2(new_n1098), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n744), .A2(new_n822), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n751), .A2(new_n1106), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n275), .B1(new_n766), .B2(new_n821), .C1(new_n771), .C2(new_n973), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n969), .B(new_n985), .C1(new_n493), .C2(new_n771), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n275), .B1(new_n765), .B2(G283), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n772), .B2(new_n751), .C1(new_n443), .C2(new_n744), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n747), .A2(new_n497), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n782), .A2(new_n480), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n739), .B1(new_n1192), .B2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1185), .A2(new_n732), .A3(new_n1186), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1184), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1182), .A2(new_n1202), .ZN(G381));
  NOR2_X1   g1003(.A1(G375), .A2(G378), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(G381), .A2(G384), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1047), .A2(new_n951), .A3(new_n980), .A4(new_n1050), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1206), .A2(G396), .A3(G393), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(G407));
  INV_X1    g1008(.A(new_n1204), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G407), .B(G213), .C1(G343), .C2(new_n1209), .ZN(G409));
  NAND2_X1  g1010(.A1(G375), .A2(G378), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n671), .A2(G213), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1119), .A2(new_n940), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1150), .B1(new_n1213), .B2(new_n1183), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1214), .A2(new_n1115), .A3(new_n1092), .A4(new_n1174), .ZN(new_n1215));
  INV_X1    g1015(.A(G384), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1016), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1081), .A2(KEYINPUT60), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1181), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1216), .B1(new_n1220), .B2(new_n1201), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1179), .A2(new_n1180), .B1(new_n1081), .B2(KEYINPUT60), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G384), .B(new_n1202), .C1(new_n1222), .C2(new_n1218), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1211), .A2(new_n1212), .A3(new_n1215), .A4(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT62), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1211), .A2(new_n1212), .A3(new_n1215), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n671), .A2(G213), .A3(G2897), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT127), .Z(new_n1229));
  AND3_X1   g1029(.A1(new_n1221), .A2(new_n1223), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1227), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT61), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G375), .A2(G378), .B1(G213), .B2(new_n671), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT62), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1215), .A4(new_n1224), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1226), .A2(new_n1233), .A3(new_n1234), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G390), .A2(G387), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1206), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(G396), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1239), .A2(new_n1206), .A3(new_n1241), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1238), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1227), .A2(KEYINPUT126), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT126), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1235), .A2(new_n1248), .A3(new_n1215), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1232), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1243), .A2(new_n1234), .A3(new_n1244), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1225), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1225), .A2(new_n1252), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1250), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1246), .A2(new_n1255), .ZN(G405));
  NAND3_X1  g1056(.A1(new_n1245), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1211), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1243), .B(new_n1244), .C1(new_n1258), .C2(new_n1204), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1257), .A2(new_n1259), .A3(new_n1224), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1224), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(G402));
endmodule


