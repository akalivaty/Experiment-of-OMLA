//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1294, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(KEYINPUT64), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(KEYINPUT64), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G97), .ZN(new_n231));
  INV_X1    g0031(.A(G257), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n209), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n212), .B(new_n221), .C1(KEYINPUT1), .C2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G97), .B(G107), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n216), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OR2_X1    g0054(.A1(KEYINPUT64), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT64), .A2(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G33), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n255), .A2(KEYINPUT65), .A3(G33), .A4(new_n256), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G77), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n262), .A2(G50), .B1(G20), .B2(new_n223), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n254), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n264), .A2(KEYINPUT11), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(KEYINPUT11), .ZN(new_n266));
  INV_X1    g0066(.A(G13), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n267), .A2(new_n207), .A3(G1), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n253), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n206), .A2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G68), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT12), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n268), .A2(new_n223), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(KEYINPUT70), .B2(KEYINPUT12), .ZN(new_n275));
  AOI211_X1 g0075(.A(new_n272), .B(new_n273), .C1(new_n268), .C2(new_n223), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n265), .A2(new_n266), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT14), .ZN(new_n279));
  INV_X1    g0079(.A(G226), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n230), .A2(G1698), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n282), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G97), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n286), .A2(KEYINPUT69), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT69), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G45), .ZN(new_n294));
  AOI21_X1  g0094(.A(G1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(new_n291), .A3(G274), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n296), .B1(new_n224), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT13), .B1(new_n292), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n286), .A2(new_n287), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT69), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n286), .A2(KEYINPUT69), .A3(new_n287), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  INV_X1    g0107(.A(new_n299), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n279), .B1(new_n310), .B2(G169), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  AOI211_X1 g0112(.A(KEYINPUT14), .B(new_n312), .C1(new_n300), .C2(new_n309), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n300), .A2(G179), .A3(new_n309), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT71), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT71), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n300), .A2(new_n317), .A3(G179), .A4(new_n309), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n278), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n291), .B1(new_n301), .B2(new_n302), .ZN(new_n321));
  AOI211_X1 g0121(.A(KEYINPUT13), .B(new_n299), .C1(new_n321), .C2(new_n304), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G190), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n310), .A2(G200), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(new_n278), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT72), .B1(new_n320), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n278), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n316), .A2(new_n318), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT14), .B1(new_n324), .B2(new_n312), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n310), .A2(new_n279), .A3(G169), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n330), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT72), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n336), .A3(new_n327), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT3), .B(G33), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(G232), .A3(new_n281), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(G238), .A3(G1698), .ZN(new_n340));
  INV_X1    g0140(.A(G107), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n339), .B(new_n340), .C1(new_n341), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n305), .ZN(new_n343));
  INV_X1    g0143(.A(G244), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n296), .B1(new_n344), .B2(new_n298), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G200), .ZN(new_n348));
  XOR2_X1   g0148(.A(KEYINPUT15), .B(G87), .Z(new_n349));
  NAND3_X1  g0149(.A1(new_n259), .A2(new_n260), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT8), .B(G58), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n255), .A2(new_n256), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n352), .A2(new_n262), .B1(new_n353), .B2(G77), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n254), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n269), .A2(G77), .A3(new_n270), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n267), .A2(G1), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G20), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(G77), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n345), .B1(new_n342), .B2(new_n305), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G190), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n348), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n361), .A2(G169), .B1(new_n355), .B2(new_n359), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n364), .A2(KEYINPUT67), .ZN(new_n365));
  INV_X1    g0165(.A(G179), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n364), .A2(KEYINPUT67), .B1(new_n366), .B2(new_n361), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n296), .B1(new_n280), .B2(new_n298), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n338), .A2(G222), .A3(new_n281), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n338), .A2(G223), .A3(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G77), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n338), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n373), .B2(new_n305), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT68), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n374), .A2(G190), .B1(new_n377), .B2(KEYINPUT10), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n377), .A2(KEYINPUT10), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n259), .A2(new_n260), .A3(new_n352), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n262), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n254), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n269), .A2(G50), .A3(new_n270), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(G50), .B2(new_n358), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT9), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT9), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n384), .B2(new_n386), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n379), .A2(new_n381), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n388), .A2(new_n376), .A3(new_n378), .A4(new_n390), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n380), .ZN(new_n393));
  INV_X1    g0193(.A(new_n387), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n374), .A2(KEYINPUT66), .A3(new_n366), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT66), .B1(new_n374), .B2(new_n366), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n394), .B1(G169), .B2(new_n374), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n368), .A2(new_n391), .A3(new_n393), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n351), .B1(new_n206), .B2(G20), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n269), .B1(new_n268), .B2(new_n351), .ZN(new_n400));
  INV_X1    g0200(.A(G223), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n281), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n280), .A2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n284), .C2(new_n285), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n305), .ZN(new_n407));
  INV_X1    g0207(.A(G190), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n293), .A2(new_n294), .ZN(new_n409));
  AND2_X1   g0209(.A1(G1), .A2(G13), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n206), .A2(new_n409), .B1(new_n410), .B2(new_n290), .ZN(new_n411));
  INV_X1    g0211(.A(G274), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n410), .B2(new_n290), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n411), .A2(G232), .B1(new_n413), .B2(new_n295), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n407), .A2(new_n408), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n291), .B1(new_n404), .B2(new_n405), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n291), .A2(G232), .A3(new_n297), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n296), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n375), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g0220(.A1(KEYINPUT3), .A2(G33), .ZN(new_n421));
  NAND2_X1  g0221(.A1(KEYINPUT3), .A2(G33), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n207), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n223), .B1(new_n423), .B2(KEYINPUT7), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n284), .A2(new_n285), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT7), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n215), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n229), .A2(new_n223), .ZN(new_n429));
  OAI21_X1  g0229(.A(G20), .B1(new_n429), .B2(new_n201), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n262), .A2(G159), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT16), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n253), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT7), .B1(new_n353), .B2(new_n338), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n425), .A2(new_n426), .A3(new_n207), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(G68), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT16), .B1(new_n439), .B2(new_n433), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n400), .B(new_n420), .C1(new_n436), .C2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT17), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n400), .B1(new_n436), .B2(new_n440), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n407), .A2(new_n366), .A3(new_n414), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n312), .B1(new_n416), .B2(new_n418), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(KEYINPUT73), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT74), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT73), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n407), .A2(new_n414), .A3(new_n448), .A4(new_n366), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n446), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n443), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT18), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n443), .C1(new_n450), .C2(new_n451), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n442), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n398), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n329), .A2(new_n337), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n215), .A2(new_n338), .A3(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n215), .A2(new_n338), .A3(new_n461), .A4(G87), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT23), .A2(G107), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(G20), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT23), .A2(G107), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n353), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT24), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT24), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n463), .A2(new_n471), .A3(new_n468), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n254), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G33), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n269), .B1(G1), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT25), .B1(new_n268), .B2(new_n341), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n268), .A2(KEYINPUT25), .A3(new_n341), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n476), .A2(G107), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n206), .B(G45), .C1(new_n293), .C2(KEYINPUT5), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT78), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n294), .A2(G1), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G41), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(KEYINPUT78), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n486), .A2(G41), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n484), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(G264), .A3(new_n291), .ZN(new_n492));
  OAI211_X1 g0292(.A(G257), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n493));
  OAI211_X1 g0293(.A(G250), .B(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G294), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n305), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n489), .B1(new_n482), .B2(new_n483), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(new_n413), .A3(new_n488), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n492), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT85), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n501), .A3(G169), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n305), .B1(new_n498), .B2(new_n488), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G264), .B1(new_n305), .B2(new_n496), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(G179), .A3(new_n499), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n501), .B1(new_n500), .B2(G169), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n473), .A2(new_n481), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n476), .A2(new_n349), .ZN(new_n509));
  INV_X1    g0309(.A(new_n349), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n268), .ZN(new_n511));
  NAND3_X1  g0311(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n255), .A2(new_n256), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n225), .A2(KEYINPUT82), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT82), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G87), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n215), .A2(new_n338), .A3(G68), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT19), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n259), .A2(G97), .A3(new_n260), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT83), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n253), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n522), .ZN(new_n527));
  INV_X1    g0327(.A(new_n521), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n527), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n509), .B(new_n511), .C1(new_n526), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT81), .ZN(new_n531));
  OAI21_X1  g0331(.A(G250), .B1(new_n294), .B2(G1), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(new_n305), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n532), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n291), .A3(KEYINPUT81), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n533), .A2(new_n535), .B1(new_n413), .B2(new_n485), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n344), .A2(new_n281), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n285), .B2(new_n284), .ZN(new_n538));
  OAI211_X1 g0338(.A(G238), .B(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G116), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n305), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(G179), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n312), .B2(new_n543), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n530), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n527), .A2(new_n528), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT83), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n524), .A2(new_n525), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n253), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n543), .A2(new_n375), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G190), .B2(new_n543), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n476), .A2(G87), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n550), .A2(new_n552), .A3(new_n511), .A4(new_n553), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n463), .A2(new_n471), .A3(new_n468), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n471), .B1(new_n463), .B2(new_n468), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n253), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n504), .A2(G190), .A3(new_n499), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n500), .A2(G200), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n557), .A2(new_n480), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n508), .A2(new_n546), .A3(new_n554), .A4(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n269), .B(G116), .C1(G1), .C2(new_n474), .ZN(new_n562));
  INV_X1    g0362(.A(G116), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n268), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n474), .A2(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G283), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n255), .A2(new_n565), .A3(new_n256), .A4(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n252), .A2(new_n216), .B1(G20), .B2(new_n563), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT20), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n567), .A2(KEYINPUT20), .A3(new_n568), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n562), .B(new_n564), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G264), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n572));
  OAI211_X1 g0372(.A(G257), .B(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n573));
  INV_X1    g0373(.A(G303), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n572), .B(new_n573), .C1(new_n574), .C2(new_n338), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n305), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n491), .A2(G270), .A3(new_n291), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n577), .A3(new_n499), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n578), .A2(KEYINPUT21), .A3(G169), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n366), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n571), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n571), .B1(G200), .B2(new_n578), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n408), .B2(new_n578), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n578), .A2(new_n571), .A3(G169), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT21), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n584), .A2(KEYINPUT84), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT84), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n581), .B(new_n583), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n561), .A2(new_n588), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n484), .A2(new_n488), .A3(new_n490), .ZN(new_n590));
  AOI22_X1  g0390(.A1(G257), .A2(new_n503), .B1(new_n590), .B2(new_n413), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT79), .ZN(new_n592));
  OAI211_X1 g0392(.A(G244), .B(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n338), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n338), .A2(G250), .A3(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n566), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n305), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n591), .A2(new_n592), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n592), .B1(new_n591), .B2(new_n599), .ZN(new_n601));
  OAI21_X1  g0401(.A(G190), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT76), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT6), .ZN(new_n604));
  AND2_X1   g0404(.A1(G97), .A2(G107), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(new_n517), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n341), .A2(KEYINPUT6), .A3(G97), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n353), .B1(G77), .B2(new_n262), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n437), .A2(G107), .A3(new_n438), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n253), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT75), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n358), .B2(G97), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n268), .A2(KEYINPUT75), .A3(new_n231), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n475), .B2(new_n231), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n603), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n254), .B1(new_n609), .B2(new_n610), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n620), .A2(KEYINPUT76), .A3(new_n617), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n598), .A2(KEYINPUT77), .A3(new_n305), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT77), .B1(new_n598), .B2(new_n305), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n591), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G200), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n602), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT80), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n598), .A2(new_n305), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n491), .A2(new_n291), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n499), .B1(new_n631), .B2(new_n232), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT79), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n591), .A2(new_n592), .A3(new_n599), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n312), .A3(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n366), .B(new_n591), .C1(new_n624), .C2(new_n625), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n612), .A2(new_n618), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n628), .A2(new_n629), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n629), .B1(new_n628), .B2(new_n638), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n589), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n458), .A2(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n397), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n365), .A2(new_n367), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT86), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT86), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n365), .A2(new_n367), .A3(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n645), .A2(new_n327), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n442), .B1(new_n648), .B2(new_n320), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n453), .A3(new_n455), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n391), .A2(new_n393), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n643), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n508), .B(new_n581), .C1(new_n587), .C2(new_n586), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n554), .A2(new_n560), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n638), .A4(new_n628), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n546), .A2(new_n554), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n612), .A2(new_n603), .A3(new_n618), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT76), .B1(new_n620), .B2(new_n617), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n635), .A2(new_n660), .A3(new_n636), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n656), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n657), .A2(new_n656), .A3(new_n638), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n655), .B(new_n546), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n652), .B1(new_n458), .B2(new_n666), .ZN(G369));
  NAND2_X1  g0467(.A1(new_n215), .A2(new_n357), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n571), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT87), .Z(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n588), .B2(KEYINPUT88), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(KEYINPUT88), .B2(new_n588), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n581), .B1(new_n586), .B2(new_n587), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n673), .B1(new_n473), .B2(new_n481), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT89), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n508), .A2(new_n560), .ZN(new_n684));
  INV_X1    g0484(.A(new_n506), .ZN(new_n685));
  INV_X1    g0485(.A(new_n507), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n685), .A2(new_n686), .B1(new_n557), .B2(new_n480), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n683), .A2(new_n684), .B1(new_n687), .B2(new_n673), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n673), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n683), .A2(new_n678), .A3(new_n684), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n690), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n689), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n210), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n206), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n518), .A2(G116), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n220), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  OAI21_X1  g0500(.A(new_n656), .B1(new_n657), .B2(new_n638), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT92), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n635), .A2(new_n660), .A3(new_n636), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(KEYINPUT26), .A3(new_n546), .A4(new_n554), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT91), .ZN(new_n706));
  INV_X1    g0506(.A(new_n657), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT91), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT26), .A4(new_n704), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT92), .B(new_n656), .C1(new_n657), .C2(new_n638), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n703), .A2(new_n706), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n628), .A2(new_n638), .A3(new_n554), .A4(new_n560), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n678), .A2(new_n687), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n546), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(KEYINPUT29), .A3(new_n690), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n665), .A2(new_n690), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  INV_X1    g0524(.A(new_n625), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n632), .B1(new_n725), .B2(new_n623), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n578), .A2(new_n500), .A3(new_n366), .A4(new_n543), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n633), .A2(new_n634), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT90), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n492), .A2(new_n497), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n730), .B1(new_n731), .B2(new_n543), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n504), .A2(KEYINPUT90), .A3(new_n542), .A4(new_n536), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n580), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n728), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n729), .A2(new_n734), .A3(KEYINPUT30), .A4(new_n580), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n724), .B(new_n690), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n580), .B1(new_n600), .B2(new_n601), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n732), .A2(new_n733), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n728), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT31), .B1(new_n744), .B2(new_n673), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n589), .B(new_n690), .C1(new_n640), .C2(new_n639), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n723), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n722), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n700), .B1(new_n749), .B2(G1), .ZN(G364));
  XOR2_X1   g0550(.A(new_n681), .B(KEYINPUT94), .Z(new_n751));
  NOR3_X1   g0551(.A1(new_n353), .A2(new_n267), .A3(new_n294), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT95), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n697), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n751), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n680), .A2(G330), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT93), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n680), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n757), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n210), .A2(new_n338), .ZN(new_n768));
  INV_X1    g0568(.A(G355), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(new_n769), .B1(G116), .B2(new_n210), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n247), .A2(new_n294), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n210), .A2(new_n425), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n294), .B2(new_n220), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n216), .B1(G20), .B2(new_n312), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n765), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n767), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n215), .A2(new_n366), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G190), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n215), .A2(G190), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G179), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G311), .A2(new_n782), .B1(new_n786), .B2(G329), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n215), .B1(G190), .B2(new_n784), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n783), .A2(new_n366), .A3(G200), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT97), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(KEYINPUT97), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n787), .B1(new_n788), .B2(new_n789), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n779), .A2(G190), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G322), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(new_n375), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G326), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n366), .A2(new_n375), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n783), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n207), .A2(new_n408), .A3(new_n375), .A4(G179), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n338), .B1(new_n806), .B2(G303), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n798), .A2(new_n800), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n785), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT32), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n341), .B2(new_n793), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G50), .A2(new_n799), .B1(new_n797), .B2(G58), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n782), .A2(G77), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n514), .A2(new_n516), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n425), .B1(new_n806), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n789), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n803), .A2(G68), .B1(new_n817), .B2(G97), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n795), .A2(new_n808), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n778), .B1(new_n820), .B2(new_n775), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n761), .B1(new_n766), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  NOR2_X1   g0623(.A1(new_n690), .A2(new_n360), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n645), .A2(new_n647), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n368), .B1(new_n360), .B2(new_n690), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n638), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n828), .A2(KEYINPUT26), .A3(new_n546), .A4(new_n554), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n662), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n690), .B(new_n827), .C1(new_n830), .C2(new_n714), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT98), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n665), .A2(KEYINPUT98), .A3(new_n690), .A4(new_n827), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n827), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n718), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n748), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n767), .B1(new_n838), .B2(new_n839), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n836), .A2(new_n763), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n775), .A2(new_n763), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n767), .B1(G77), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n793), .A2(new_n225), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G311), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n563), .A2(new_n781), .B1(new_n785), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G283), .B2(new_n803), .ZN(new_n851));
  INV_X1    g0651(.A(new_n806), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n425), .B1(new_n852), .B2(new_n341), .C1(new_n231), .C2(new_n789), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G294), .B2(new_n797), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n799), .A2(G303), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n848), .A2(new_n851), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n793), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(G68), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n338), .B1(new_n852), .B2(new_n202), .C1(new_n229), .C2(new_n789), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G132), .B2(new_n786), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G150), .A2(new_n803), .B1(new_n782), .B2(G159), .ZN(new_n861));
  INV_X1    g0661(.A(new_n797), .ZN(new_n862));
  INV_X1    g0662(.A(G143), .ZN(new_n863));
  INV_X1    g0663(.A(G137), .ZN(new_n864));
  INV_X1    g0664(.A(new_n799), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n861), .B1(new_n862), .B2(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT34), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n858), .B(new_n860), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n856), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n846), .B1(new_n870), .B2(new_n775), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n841), .A2(new_n842), .B1(new_n843), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  AOI21_X1  g0673(.A(new_n206), .B1(new_n215), .B2(G13), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n319), .A2(new_n332), .A3(new_n333), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n328), .B1(new_n875), .B2(new_n330), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT99), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n278), .A2(new_n690), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n335), .A2(KEYINPUT99), .A3(new_n327), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n314), .A2(new_n319), .A3(new_n327), .A4(new_n879), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(new_n836), .ZN(new_n887));
  INV_X1    g0687(.A(new_n671), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n450), .A2(new_n451), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n432), .B1(new_n427), .B2(new_n424), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n254), .B1(new_n890), .B2(KEYINPUT16), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT100), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n435), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n434), .A2(KEYINPUT100), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n400), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n441), .B1(new_n889), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT101), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT37), .ZN(new_n900));
  INV_X1    g0700(.A(new_n441), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n446), .A2(new_n449), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT74), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(new_n671), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n901), .B1(new_n905), .B2(new_n896), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT101), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n443), .A2(new_n888), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n452), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n441), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n900), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n456), .A2(new_n888), .A3(new_n896), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(KEYINPUT38), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  INV_X1    g0720(.A(new_n745), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n747), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n887), .A2(new_n919), .A3(new_n920), .A4(new_n923), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n878), .A2(new_n880), .B1(new_n882), .B2(new_n884), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n923), .A3(new_n827), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT105), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n918), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n913), .A2(KEYINPUT105), .A3(KEYINPUT38), .A4(new_n914), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT103), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n452), .A2(new_n931), .A3(new_n909), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n452), .A2(new_n441), .A3(new_n909), .ZN(new_n933));
  INV_X1    g0733(.A(new_n911), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n932), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT104), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n910), .B(new_n441), .C1(new_n931), .C2(new_n911), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT104), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n456), .A2(new_n443), .A3(new_n888), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n916), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n926), .B1(new_n930), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n924), .B1(new_n945), .B2(new_n920), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT106), .Z(new_n947));
  AOI21_X1  g0747(.A(new_n458), .B1(new_n747), .B2(new_n746), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n949), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(G330), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n644), .A2(new_n673), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n833), .B2(new_n834), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n919), .A3(new_n925), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n335), .A2(new_n673), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n928), .A2(new_n929), .B1(new_n916), .B2(new_n943), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n957), .B(new_n958), .C1(new_n959), .C2(KEYINPUT39), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n453), .A2(new_n455), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n671), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n956), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n458), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n717), .A2(new_n964), .A3(new_n720), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n652), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n963), .B(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n874), .B1(new_n952), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n952), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n608), .A2(KEYINPUT35), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n608), .A2(KEYINPUT35), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n970), .A2(G116), .A3(new_n217), .A4(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT36), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n219), .A2(new_n372), .A3(new_n429), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n223), .A2(G50), .ZN(new_n975));
  OAI211_X1 g0775(.A(G1), .B(new_n267), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n969), .A2(new_n973), .A3(new_n976), .ZN(G367));
  OAI221_X1 g0777(.A(new_n776), .B1(new_n210), .B2(new_n510), .C1(new_n243), .C2(new_n772), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n767), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n775), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n788), .A2(new_n802), .B1(new_n785), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n852), .A2(new_n563), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n425), .B1(new_n983), .B2(KEYINPUT46), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(G283), .C2(new_n782), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n574), .B2(new_n862), .C1(new_n849), .C2(new_n865), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n857), .A2(G97), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(KEYINPUT46), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT109), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n988), .A2(new_n989), .B1(G107), .B2(new_n817), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(new_n989), .C2(new_n988), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n338), .B1(new_n852), .B2(new_n229), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G137), .B2(new_n786), .ZN(new_n993));
  INV_X1    g0793(.A(G150), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n993), .B1(new_n862), .B2(new_n994), .C1(new_n863), .C2(new_n865), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n857), .A2(G77), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n817), .A2(G68), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G50), .A2(new_n782), .B1(new_n803), .B2(G159), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n986), .A2(new_n991), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT47), .Z(new_n1001));
  NAND3_X1  g0801(.A1(new_n550), .A2(new_n511), .A3(new_n553), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n673), .ZN(new_n1003));
  MUX2_X1   g0803(.A(new_n546), .B(new_n657), .S(new_n1003), .Z(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT107), .Z(new_n1005));
  INV_X1    g0805(.A(new_n765), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n979), .B1(new_n980), .B2(new_n1001), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n628), .B(new_n638), .C1(new_n622), .C2(new_n690), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n635), .A2(new_n660), .A3(new_n636), .A4(new_n673), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n1011), .A2(new_n691), .A3(KEYINPUT108), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT108), .B1(new_n1011), .B2(new_n691), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT42), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n638), .B1(new_n1011), .B2(new_n508), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1014), .A2(KEYINPUT42), .B1(new_n690), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1005), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT43), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1015), .A2(new_n1017), .A3(new_n1020), .A4(new_n1019), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n689), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(new_n1011), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1025), .B(new_n1027), .Z(new_n1028));
  NOR2_X1   g0828(.A1(new_n755), .A2(new_n206), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n693), .A2(new_n1011), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n693), .A2(new_n1011), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT44), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n689), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1032), .A2(new_n1026), .A3(new_n1035), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n678), .A2(new_n690), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n688), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n691), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n751), .A2(new_n1042), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n681), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n749), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n696), .B(KEYINPUT41), .Z(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1030), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1007), .B1(new_n1028), .B2(new_n1049), .ZN(G387));
  INV_X1    g0850(.A(new_n1045), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n688), .A2(new_n765), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n240), .A2(new_n294), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1053), .A2(new_n772), .B1(new_n698), .B2(new_n768), .ZN(new_n1054));
  AOI21_X1  g0854(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n352), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT50), .B1(new_n352), .B2(new_n202), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n698), .B(new_n1055), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1054), .A2(new_n1058), .B1(new_n341), .B2(new_n695), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n767), .B1(new_n1059), .B2(new_n777), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n789), .A2(new_n510), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n802), .B2(new_n351), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G150), .B2(new_n786), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n799), .A2(G159), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n338), .B1(new_n852), .B2(new_n372), .C1(new_n781), .C2(new_n223), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G50), .B2(new_n797), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n987), .A2(new_n1064), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n789), .A2(new_n794), .B1(new_n852), .B2(new_n788), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G303), .A2(new_n782), .B1(new_n803), .B2(G311), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n799), .A2(G322), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n981), .C2(new_n862), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT49), .Z(new_n1076));
  AOI21_X1  g0876(.A(new_n338), .B1(new_n786), .B2(G326), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n793), .B2(new_n563), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1068), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1060), .B1(new_n1079), .B2(new_n775), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1051), .A2(new_n1030), .B1(new_n1052), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1051), .A2(new_n749), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n696), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1051), .A2(new_n749), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(G393));
  INV_X1    g0885(.A(new_n1039), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n1030), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n776), .B1(new_n231), .B2(new_n210), .C1(new_n250), .C2(new_n772), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT110), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1090), .A2(new_n767), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n425), .B1(new_n852), .B2(new_n794), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G294), .A2(new_n782), .B1(new_n786), .B2(G322), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n574), .B2(new_n802), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(G116), .C2(new_n817), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n341), .B2(new_n793), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G311), .A2(new_n797), .B1(new_n799), .B2(G317), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT52), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G143), .A2(new_n786), .B1(new_n782), .B2(new_n352), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n372), .B2(new_n789), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n338), .B1(new_n852), .B2(new_n223), .C1(new_n802), .C2(new_n202), .ZN(new_n1102));
  OR3_X1    g0902(.A1(new_n847), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G150), .A2(new_n799), .B1(new_n797), .B2(G159), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1097), .A2(new_n1099), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT112), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1092), .B1(new_n1006), .B2(new_n1010), .C1(new_n1108), .C2(new_n980), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n696), .B1(new_n1082), .B2(new_n1039), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1086), .B1(new_n749), .B2(new_n1051), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1087), .B(new_n1109), .C1(new_n1110), .C2(new_n1111), .ZN(G390));
  NAND3_X1  g0912(.A1(new_n748), .A2(new_n827), .A3(new_n925), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(KEYINPUT115), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n957), .B1(new_n930), .B2(new_n944), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT113), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n881), .A2(new_n1117), .A3(new_n885), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n879), .B1(new_n876), .B2(new_n877), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n883), .B1(new_n876), .B2(KEYINPUT99), .ZN(new_n1120));
  OAI21_X1  g0920(.A(KEYINPUT113), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n673), .B(new_n836), .C1(new_n711), .C2(new_n715), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n953), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1116), .A2(KEYINPUT114), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT114), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n954), .A2(new_n886), .B1(new_n335), .B2(new_n673), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n958), .B1(new_n959), .B2(KEYINPUT39), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1113), .A2(KEYINPUT115), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1115), .B1(new_n1127), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1131), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1135), .B(new_n1114), .C1(new_n1126), .C2(new_n1125), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1030), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1129), .A2(new_n763), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n767), .B1(new_n352), .B2(new_n845), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT120), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n802), .A2(new_n864), .B1(new_n789), .B2(new_n809), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT54), .B(G143), .Z(new_n1143));
  AND2_X1   g0943(.A1(new_n782), .A2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(G125), .C2(new_n786), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n799), .A2(G128), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n852), .A2(KEYINPUT53), .A3(new_n994), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT53), .B1(new_n852), .B2(new_n994), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n338), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1147), .B(new_n1149), .C1(G132), .C2(new_n797), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n857), .A2(G50), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1145), .A2(new_n1146), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n231), .A2(new_n781), .B1(new_n785), .B2(new_n788), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G107), .B2(new_n803), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n425), .B1(new_n852), .B2(new_n225), .C1(new_n372), .C2(new_n789), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G116), .B2(new_n797), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n799), .A2(G283), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n858), .A2(new_n1154), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1152), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1139), .B(new_n1141), .C1(new_n980), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1138), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n696), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT117), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n923), .A2(G330), .A3(new_n827), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n673), .B1(new_n711), .B2(new_n715), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n953), .B1(new_n1167), .B2(new_n827), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1166), .A2(new_n1113), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1165), .A2(new_n886), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n954), .B1(new_n1113), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT116), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n948), .B2(G330), .ZN(new_n1174));
  AND4_X1   g0974(.A1(new_n1173), .A2(new_n964), .A3(G330), .A4(new_n923), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n652), .B(new_n965), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1164), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(new_n966), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1166), .A2(new_n1113), .A3(new_n1168), .ZN(new_n1180));
  AND4_X1   g0980(.A1(G330), .A2(new_n925), .A3(new_n923), .A4(new_n827), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n925), .B1(new_n748), .B2(new_n827), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1180), .B1(new_n1183), .B2(new_n954), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1179), .A2(new_n1184), .A3(KEYINPUT117), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1177), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1163), .B1(new_n1137), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT119), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT118), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1179), .A2(new_n1184), .A3(KEYINPUT117), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT117), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1177), .A2(KEYINPUT118), .A3(new_n1185), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1187), .A2(new_n1188), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1188), .B1(new_n1187), .B2(new_n1194), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1162), .B1(new_n1195), .B2(new_n1196), .ZN(G378));
  AOI21_X1  g0997(.A(new_n757), .B1(new_n202), .B2(new_n844), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n793), .A2(new_n229), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT121), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n997), .B1(new_n865), .B2(new_n563), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT122), .Z(new_n1202));
  OAI22_X1  g1002(.A1(new_n231), .A2(new_n802), .B1(new_n785), .B2(new_n794), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n338), .A2(G41), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n852), .B2(new_n372), .C1(new_n781), .C2(new_n510), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G107), .C2(new_n797), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1200), .A2(new_n1202), .A3(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT123), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT58), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G50), .B(new_n1204), .C1(new_n474), .C2(new_n293), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G132), .A2(new_n803), .B1(new_n782), .B2(G137), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n817), .A2(G150), .B1(new_n806), .B2(new_n1143), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n797), .A2(G128), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n799), .A2(G125), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n857), .A2(G159), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(G41), .C1(new_n786), .C2(G124), .ZN(new_n1221));
  AND4_X1   g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n651), .A2(new_n397), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n387), .A2(new_n671), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1224), .B(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1226), .B(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1198), .B1(new_n1223), .B2(new_n980), .C1(new_n1229), .C2(new_n764), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n946), .A2(G330), .A3(new_n1229), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1229), .B1(new_n946), .B2(G330), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n963), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n946), .A2(G330), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1228), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n963), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1232), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1231), .B1(new_n1240), .B2(new_n1030), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1136), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1116), .A2(new_n1124), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT114), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1116), .A2(new_n1124), .A3(KEYINPUT114), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1114), .B1(new_n1247), .B2(new_n1135), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1186), .B1(new_n1242), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1179), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1250), .B2(new_n1240), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1176), .B1(new_n1137), .B2(new_n1186), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1233), .A2(new_n1234), .A3(new_n963), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1238), .B1(new_n1237), .B2(new_n1232), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n696), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1241), .B1(new_n1251), .B2(new_n1256), .ZN(G375));
  NAND3_X1  g1057(.A1(new_n1118), .A2(new_n1121), .A3(new_n763), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n767), .B1(G68), .B2(new_n845), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n797), .A2(G283), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n338), .B1(new_n806), .B2(G97), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1062), .A3(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G107), .A2(new_n782), .B1(new_n786), .B2(G303), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n996), .B(new_n1263), .C1(new_n563), .C2(new_n802), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1262), .B(new_n1264), .C1(G294), .C2(new_n799), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(KEYINPUT124), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(KEYINPUT124), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n817), .A2(G50), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G128), .A2(new_n786), .B1(new_n803), .B2(new_n1143), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n338), .B1(new_n852), .B2(new_n809), .C1(new_n781), .C2(new_n994), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n862), .A2(new_n864), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1270), .B(new_n1271), .C1(G132), .C2(new_n799), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1200), .A2(new_n1268), .A3(new_n1269), .A4(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1266), .A2(new_n1267), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1259), .B1(new_n1274), .B2(new_n775), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1184), .A2(new_n1030), .B1(new_n1258), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1048), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1277), .B2(new_n1279), .ZN(G381));
  INV_X1    g1080(.A(new_n1241), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT57), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1163), .B1(new_n1250), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1240), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1282), .B1(new_n1252), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1281), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(KEYINPUT125), .ZN(new_n1288));
  OR4_X1    g1088(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1289));
  OR3_X1    g1089(.A1(new_n1289), .A2(G387), .A3(G381), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1161), .B1(new_n1194), .B2(new_n1187), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OR3_X1    g1092(.A1(new_n1288), .A2(new_n1290), .A3(new_n1292), .ZN(G407));
  NAND2_X1  g1093(.A1(new_n672), .A2(G213), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G407), .B(G213), .C1(new_n1288), .C2(new_n1296), .ZN(G409));
  NAND3_X1  g1097(.A1(new_n1250), .A2(new_n1048), .A3(new_n1240), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1241), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1291), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1277), .A2(new_n1137), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1249), .A2(new_n696), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT119), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1187), .A2(new_n1194), .A3(new_n1188), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1161), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1300), .B1(new_n1305), .B2(G375), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1278), .A2(KEYINPUT126), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT60), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT60), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1278), .A2(KEYINPUT126), .A3(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(new_n696), .A3(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1186), .A2(new_n1278), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1276), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n872), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G384), .B(new_n1276), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1294), .A4(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(G390), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G387), .A2(new_n1319), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(G393), .B(new_n822), .ZN(new_n1321));
  OAI211_X1 g1121(.A(G390), .B(new_n1007), .C1(new_n1049), .C2(new_n1028), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1321), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1323), .A2(new_n1324), .A3(KEYINPUT61), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1318), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1295), .A2(G2897), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1314), .A2(new_n1315), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1327), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(G378), .A2(new_n1287), .B1(new_n1291), .B2(new_n1299), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1330), .B(KEYINPUT127), .C1(new_n1331), .C2(new_n1295), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1306), .A2(new_n1294), .A3(new_n1317), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1330), .B1(new_n1331), .B2(new_n1295), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT127), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1326), .A2(new_n1332), .A3(new_n1335), .A4(new_n1338), .ZN(new_n1339));
  OR2_X1    g1139(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1306), .A2(new_n1341), .A3(new_n1294), .A4(new_n1317), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1336), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(G378), .A2(new_n1287), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1295), .B1(new_n1345), .B2(new_n1300), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1341), .B1(new_n1346), .B2(new_n1317), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1340), .B1(new_n1344), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1339), .A2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(G375), .A2(new_n1291), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1345), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1317), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1345), .A2(new_n1350), .A3(new_n1316), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1354), .B(new_n1340), .ZN(G402));
endmodule


