

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756;

  NOR2_X1 U375 ( .A1(n577), .A2(n694), .ZN(n576) );
  XNOR2_X1 U376 ( .A(n510), .B(n511), .ZN(n735) );
  AND2_X2 U377 ( .A1(n387), .A2(n369), .ZN(n721) );
  INV_X1 U378 ( .A(G953), .ZN(n730) );
  XNOR2_X1 U379 ( .A(n581), .B(n580), .ZN(n678) );
  NOR2_X2 U380 ( .A1(n563), .A2(n605), .ZN(n561) );
  XNOR2_X2 U381 ( .A(n425), .B(KEYINPUT22), .ZN(n563) );
  XNOR2_X2 U382 ( .A(G101), .B(G113), .ZN(n437) );
  XNOR2_X1 U383 ( .A(n527), .B(KEYINPUT19), .ZN(n591) );
  AND2_X1 U384 ( .A1(n374), .A2(n373), .ZN(n372) );
  AND2_X1 U385 ( .A1(n460), .A2(n364), .ZN(n373) );
  NOR2_X1 U386 ( .A1(n380), .A2(n462), .ZN(n461) );
  XNOR2_X1 U387 ( .A(n397), .B(n423), .ZN(n641) );
  AND2_X1 U388 ( .A1(n415), .A2(n427), .ZN(n392) );
  AND2_X1 U389 ( .A1(n408), .A2(n407), .ZN(n452) );
  NOR2_X1 U390 ( .A1(n756), .A2(n753), .ZN(n390) );
  XNOR2_X1 U391 ( .A(n623), .B(KEYINPUT42), .ZN(n756) );
  AND2_X1 U392 ( .A1(n421), .A2(n420), .ZN(n657) );
  XNOR2_X1 U393 ( .A(n424), .B(KEYINPUT41), .ZN(n698) );
  NOR2_X1 U394 ( .A1(n703), .A2(n701), .ZN(n424) );
  XNOR2_X1 U395 ( .A(n382), .B(n381), .ZN(n703) );
  NAND2_X1 U396 ( .A1(n591), .A2(n533), .ZN(n535) );
  NAND2_X1 U397 ( .A1(n595), .A2(n699), .ZN(n527) );
  XNOR2_X1 U398 ( .A(n472), .B(KEYINPUT65), .ZN(n688) );
  OR2_X2 U399 ( .A1(n402), .A2(n401), .ZN(n691) );
  XNOR2_X1 U400 ( .A(n560), .B(n559), .ZN(n684) );
  XOR2_X1 U401 ( .A(G116), .B(G107), .Z(n509) );
  XNOR2_X1 U402 ( .A(n485), .B(n484), .ZN(n590) );
  INV_X1 U403 ( .A(n652), .ZN(n440) );
  AND2_X1 U404 ( .A1(n375), .A2(n602), .ZN(n579) );
  XNOR2_X1 U405 ( .A(n376), .B(KEYINPUT91), .ZN(n375) );
  NOR2_X1 U406 ( .A1(n671), .A2(n657), .ZN(n376) );
  OR2_X1 U407 ( .A1(G237), .A2(G902), .ZN(n523) );
  XNOR2_X1 U408 ( .A(G902), .B(KEYINPUT15), .ZN(n637) );
  XNOR2_X1 U409 ( .A(n675), .B(n453), .ZN(n407) );
  INV_X1 U410 ( .A(KEYINPUT81), .ZN(n453) );
  NAND2_X1 U411 ( .A1(G214), .A2(n523), .ZN(n699) );
  NAND2_X1 U412 ( .A1(n648), .A2(G472), .ZN(n403) );
  OR2_X1 U413 ( .A1(n684), .A2(n683), .ZN(n472) );
  NAND2_X1 U414 ( .A1(n385), .A2(n371), .ZN(n387) );
  XNOR2_X1 U415 ( .A(n384), .B(n386), .ZN(n385) );
  NAND2_X1 U416 ( .A1(n641), .A2(n383), .ZN(n384) );
  NAND2_X1 U417 ( .A1(n454), .A2(n590), .ZN(n622) );
  XNOR2_X1 U418 ( .A(n589), .B(n455), .ZN(n454) );
  XNOR2_X1 U419 ( .A(KEYINPUT28), .B(KEYINPUT103), .ZN(n455) );
  INV_X1 U420 ( .A(KEYINPUT6), .ZN(n409) );
  NAND2_X1 U421 ( .A1(n612), .A2(n664), .ZN(n379) );
  INV_X1 U422 ( .A(KEYINPUT76), .ZN(n378) );
  XNOR2_X1 U423 ( .A(G146), .B(G125), .ZN(n512) );
  AND2_X1 U424 ( .A1(n752), .A2(n457), .ZN(n456) );
  NOR2_X1 U425 ( .A1(n579), .A2(n440), .ZN(n427) );
  XNOR2_X1 U426 ( .A(n524), .B(KEYINPUT75), .ZN(n525) );
  XOR2_X1 U427 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n539) );
  INV_X1 U428 ( .A(KEYINPUT71), .ZN(n540) );
  XNOR2_X1 U429 ( .A(G137), .B(G116), .ZN(n541) );
  XNOR2_X1 U430 ( .A(n480), .B(G143), .ZN(n486) );
  INV_X1 U431 ( .A(G128), .ZN(n480) );
  XNOR2_X1 U432 ( .A(n500), .B(n496), .ZN(n464) );
  XNOR2_X1 U433 ( .A(G113), .B(G143), .ZN(n496) );
  XNOR2_X1 U434 ( .A(G131), .B(KEYINPUT12), .ZN(n497) );
  INV_X1 U435 ( .A(KEYINPUT48), .ZN(n423) );
  XNOR2_X1 U436 ( .A(n519), .B(n451), .ZN(n741) );
  XNOR2_X1 U437 ( .A(n396), .B(G134), .ZN(n451) );
  XNOR2_X1 U438 ( .A(G131), .B(KEYINPUT4), .ZN(n396) );
  XOR2_X1 U439 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n517) );
  AND2_X1 U440 ( .A1(n605), .A2(n699), .ZN(n606) );
  XNOR2_X1 U441 ( .A(n502), .B(n458), .ZN(n572) );
  XNOR2_X1 U442 ( .A(n501), .B(n459), .ZN(n458) );
  INV_X1 U443 ( .A(G475), .ZN(n459) );
  XNOR2_X1 U444 ( .A(n549), .B(n548), .ZN(n553) );
  XNOR2_X1 U445 ( .A(G119), .B(G128), .ZN(n548) );
  XOR2_X1 U446 ( .A(KEYINPUT24), .B(G110), .Z(n549) );
  XOR2_X1 U447 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n552) );
  XNOR2_X1 U448 ( .A(n469), .B(n467), .ZN(n550) );
  XNOR2_X1 U449 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n469) );
  NOR2_X1 U450 ( .A1(n468), .A2(G953), .ZN(n467) );
  INV_X1 U451 ( .A(G234), .ZN(n468) );
  XNOR2_X1 U452 ( .A(n446), .B(n567), .ZN(n709) );
  OR2_X1 U453 ( .A1(n411), .A2(n355), .ZN(n625) );
  NOR2_X1 U454 ( .A1(n709), .A2(n577), .ZN(n568) );
  XNOR2_X1 U455 ( .A(n610), .B(n476), .ZN(n615) );
  INV_X1 U456 ( .A(KEYINPUT72), .ZN(n476) );
  NAND2_X1 U457 ( .A1(n566), .A2(n426), .ZN(n425) );
  AND2_X1 U458 ( .A1(n506), .A2(n505), .ZN(n426) );
  NAND2_X1 U459 ( .A1(n403), .A2(n406), .ZN(n402) );
  NAND2_X1 U460 ( .A1(G472), .A2(G902), .ZN(n406) );
  XOR2_X1 U461 ( .A(n590), .B(KEYINPUT1), .Z(n626) );
  XNOR2_X1 U462 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U463 ( .A1(n372), .A2(n370), .ZN(n369) );
  NAND2_X1 U464 ( .A1(n371), .A2(n461), .ZN(n370) );
  NOR2_X1 U465 ( .A1(G953), .A2(G237), .ZN(n537) );
  AND2_X1 U466 ( .A1(n377), .A2(n359), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n379), .B(n378), .ZN(n377) );
  INV_X1 U468 ( .A(KEYINPUT69), .ZN(n428) );
  NAND2_X1 U469 ( .A1(n640), .A2(n641), .ZN(n380) );
  INV_X1 U470 ( .A(KEYINPUT78), .ZN(n462) );
  AND2_X1 U471 ( .A1(n639), .A2(KEYINPUT2), .ZN(n383) );
  NAND2_X1 U472 ( .A1(G234), .A2(G237), .ZN(n528) );
  INV_X1 U473 ( .A(KEYINPUT105), .ZN(n381) );
  NAND2_X1 U474 ( .A1(n574), .A2(n572), .ZN(n701) );
  INV_X1 U475 ( .A(n699), .ZN(n410) );
  INV_X1 U476 ( .A(n701), .ZN(n506) );
  NAND2_X1 U477 ( .A1(n546), .A2(n405), .ZN(n404) );
  INV_X1 U478 ( .A(G902), .ZN(n405) );
  XNOR2_X1 U479 ( .A(n438), .B(n545), .ZN(n648) );
  XNOR2_X1 U480 ( .A(n439), .B(n544), .ZN(n438) );
  XNOR2_X1 U481 ( .A(G134), .B(G122), .ZN(n489) );
  XNOR2_X1 U482 ( .A(n499), .B(n466), .ZN(n465) );
  XNOR2_X1 U483 ( .A(n741), .B(n450), .ZN(n545) );
  INV_X1 U484 ( .A(G146), .ZN(n450) );
  INV_X1 U485 ( .A(G101), .ZN(n481) );
  XNOR2_X1 U486 ( .A(G107), .B(G104), .ZN(n482) );
  XNOR2_X1 U487 ( .A(n429), .B(n522), .ZN(n644) );
  XNOR2_X1 U488 ( .A(n735), .B(n515), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n399), .B(n617), .ZN(n633) );
  AND2_X1 U490 ( .A1(n616), .A2(n621), .ZN(n400) );
  NOR2_X1 U491 ( .A1(n626), .A2(n445), .ZN(n575) );
  INV_X1 U492 ( .A(n688), .ZN(n445) );
  NOR2_X1 U493 ( .A1(n622), .A2(n592), .ZN(n593) );
  XNOR2_X1 U494 ( .A(n691), .B(n547), .ZN(n605) );
  INV_X1 U495 ( .A(KEYINPUT95), .ZN(n547) );
  XNOR2_X1 U496 ( .A(n471), .B(n740), .ZN(n650) );
  XNOR2_X1 U497 ( .A(n545), .B(n447), .ZN(n724) );
  XNOR2_X1 U498 ( .A(n449), .B(n448), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n554), .B(n357), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n483), .B(n513), .ZN(n449) );
  NOR2_X1 U501 ( .A1(KEYINPUT2), .A2(n371), .ZN(n679) );
  NOR2_X1 U502 ( .A1(n625), .A2(n629), .ZN(n600) );
  INV_X1 U503 ( .A(KEYINPUT35), .ZN(n442) );
  NAND2_X1 U504 ( .A1(n569), .A2(n354), .ZN(n443) );
  XNOR2_X1 U505 ( .A(n389), .B(KEYINPUT32), .ZN(n755) );
  OR2_X1 U506 ( .A1(n353), .A2(n597), .ZN(n388) );
  NAND2_X1 U507 ( .A1(n611), .A2(n354), .ZN(n664) );
  XNOR2_X1 U508 ( .A(n474), .B(n473), .ZN(n611) );
  INV_X1 U509 ( .A(KEYINPUT102), .ZN(n473) );
  INV_X1 U510 ( .A(KEYINPUT89), .ZN(n422) );
  INV_X1 U511 ( .A(KEYINPUT83), .ZN(n413) );
  INV_X1 U512 ( .A(KEYINPUT56), .ZN(n393) );
  OR2_X1 U513 ( .A1(n583), .A2(n626), .ZN(n353) );
  XOR2_X1 U514 ( .A(n565), .B(KEYINPUT97), .Z(n354) );
  XNOR2_X1 U515 ( .A(n691), .B(n409), .ZN(n597) );
  OR2_X1 U516 ( .A1(n618), .A2(n410), .ZN(n355) );
  AND2_X1 U517 ( .A1(n590), .A2(n609), .ZN(n356) );
  AND2_X1 U518 ( .A1(G227), .A2(n730), .ZN(n357) );
  NOR2_X1 U519 ( .A1(KEYINPUT2), .A2(n742), .ZN(n358) );
  NAND2_X1 U520 ( .A1(n594), .A2(n603), .ZN(n359) );
  XOR2_X1 U521 ( .A(n642), .B(n477), .Z(n360) );
  XOR2_X1 U522 ( .A(n648), .B(KEYINPUT62), .Z(n361) );
  XOR2_X1 U523 ( .A(n724), .B(n478), .Z(n362) );
  XOR2_X1 U524 ( .A(n650), .B(KEYINPUT122), .Z(n363) );
  OR2_X1 U525 ( .A1(n636), .A2(n635), .ZN(n364) );
  XOR2_X1 U526 ( .A(n646), .B(n645), .Z(n365) );
  XOR2_X1 U527 ( .A(n624), .B(KEYINPUT46), .Z(n366) );
  NOR2_X1 U528 ( .A1(G952), .A2(n730), .ZN(n729) );
  INV_X1 U529 ( .A(n729), .ZN(n434) );
  XNOR2_X1 U530 ( .A(KEYINPUT60), .B(KEYINPUT121), .ZN(n367) );
  XOR2_X1 U531 ( .A(KEYINPUT63), .B(KEYINPUT107), .Z(n368) );
  INV_X1 U532 ( .A(n678), .ZN(n371) );
  NAND2_X1 U533 ( .A1(n678), .A2(n462), .ZN(n374) );
  NAND2_X1 U534 ( .A1(n688), .A2(n590), .ZN(n608) );
  NAND2_X1 U535 ( .A1(n688), .A2(n356), .ZN(n610) );
  NAND2_X1 U536 ( .A1(n380), .A2(n462), .ZN(n460) );
  NAND2_X1 U537 ( .A1(n621), .A2(n699), .ZN(n382) );
  XNOR2_X2 U538 ( .A(n613), .B(n614), .ZN(n621) );
  AND2_X1 U539 ( .A1(n641), .A2(n639), .ZN(n742) );
  INV_X1 U540 ( .A(n387), .ZN(n681) );
  INV_X1 U541 ( .A(KEYINPUT80), .ZN(n386) );
  OR2_X1 U542 ( .A1(n563), .A2(n597), .ZN(n414) );
  NOR2_X1 U543 ( .A1(n563), .A2(n388), .ZN(n389) );
  XNOR2_X1 U544 ( .A(n390), .B(n366), .ZN(n398) );
  AND2_X1 U545 ( .A1(n391), .A2(n434), .ZN(G54) );
  XNOR2_X1 U546 ( .A(n725), .B(n362), .ZN(n391) );
  NAND2_X1 U547 ( .A1(n417), .A2(n392), .ZN(n581) );
  XNOR2_X1 U548 ( .A(n394), .B(n393), .ZN(G51) );
  NAND2_X1 U549 ( .A1(n433), .A2(n434), .ZN(n394) );
  XNOR2_X1 U550 ( .A(n395), .B(n367), .ZN(G60) );
  NAND2_X1 U551 ( .A1(n435), .A2(n434), .ZN(n395) );
  XNOR2_X1 U552 ( .A(n418), .B(n428), .ZN(n417) );
  NAND2_X1 U553 ( .A1(n398), .A2(n452), .ZN(n397) );
  NOR2_X1 U554 ( .A1(n633), .A2(n618), .ZN(n620) );
  NAND2_X1 U555 ( .A1(n615), .A2(n400), .ZN(n399) );
  NOR2_X1 U556 ( .A1(n648), .A2(n404), .ZN(n401) );
  NAND2_X1 U557 ( .A1(n601), .A2(n687), .ZN(n675) );
  XNOR2_X1 U558 ( .A(n598), .B(n412), .ZN(n411) );
  INV_X1 U559 ( .A(KEYINPUT98), .ZN(n412) );
  XNOR2_X1 U560 ( .A(n414), .B(n413), .ZN(n570) );
  NAND2_X1 U561 ( .A1(n416), .A2(KEYINPUT44), .ZN(n415) );
  NAND2_X1 U562 ( .A1(n419), .A2(n752), .ZN(n416) );
  NAND2_X1 U563 ( .A1(n419), .A2(n456), .ZN(n418) );
  XNOR2_X1 U564 ( .A(n564), .B(KEYINPUT84), .ZN(n419) );
  INV_X1 U565 ( .A(n691), .ZN(n420) );
  XNOR2_X1 U566 ( .A(n578), .B(n422), .ZN(n421) );
  XNOR2_X2 U567 ( .A(n535), .B(n534), .ZN(n566) );
  XNOR2_X1 U568 ( .A(n430), .B(n368), .ZN(G57) );
  NAND2_X1 U569 ( .A1(n441), .A2(n434), .ZN(n430) );
  AND2_X1 U570 ( .A1(n680), .A2(n431), .ZN(n718) );
  NOR2_X1 U571 ( .A1(n681), .A2(n358), .ZN(n431) );
  XNOR2_X1 U572 ( .A(n432), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U573 ( .A1(n436), .A2(n434), .ZN(n432) );
  XNOR2_X1 U574 ( .A(n647), .B(n365), .ZN(n433) );
  XNOR2_X1 U575 ( .A(n643), .B(n360), .ZN(n435) );
  XNOR2_X1 U576 ( .A(n651), .B(n363), .ZN(n436) );
  INV_X1 U577 ( .A(n437), .ZN(n479) );
  INV_X1 U578 ( .A(n536), .ZN(n439) );
  XNOR2_X1 U579 ( .A(n649), .B(n361), .ZN(n441) );
  XNOR2_X2 U580 ( .A(n526), .B(n525), .ZN(n595) );
  NOR2_X1 U581 ( .A1(n650), .A2(G902), .ZN(n560) );
  XNOR2_X2 U582 ( .A(n443), .B(n442), .ZN(n752) );
  NAND2_X1 U583 ( .A1(n687), .A2(n444), .ZN(n446) );
  AND2_X1 U584 ( .A1(n597), .A2(n688), .ZN(n444) );
  INV_X1 U585 ( .A(KEYINPUT44), .ZN(n457) );
  XNOR2_X1 U586 ( .A(n465), .B(n463), .ZN(n642) );
  XNOR2_X1 U587 ( .A(n555), .B(n464), .ZN(n463) );
  INV_X1 U588 ( .A(n507), .ZN(n466) );
  XNOR2_X1 U589 ( .A(n470), .B(n551), .ZN(n471) );
  XNOR2_X1 U590 ( .A(n553), .B(n552), .ZN(n470) );
  NAND2_X1 U591 ( .A1(n615), .A2(n475), .ZN(n474) );
  AND2_X1 U592 ( .A1(n616), .A2(n613), .ZN(n475) );
  XNOR2_X1 U593 ( .A(KEYINPUT59), .B(KEYINPUT85), .ZN(n477) );
  XOR2_X1 U594 ( .A(n723), .B(n722), .Z(n478) );
  INV_X1 U595 ( .A(KEYINPUT64), .ZN(n624) );
  XNOR2_X1 U596 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U598 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U599 ( .A(KEYINPUT0), .ZN(n534) );
  INV_X1 U600 ( .A(G472), .ZN(n546) );
  INV_X1 U601 ( .A(n486), .ZN(n519) );
  XOR2_X1 U602 ( .A(G137), .B(G140), .Z(n554) );
  XOR2_X1 U603 ( .A(KEYINPUT68), .B(G110), .Z(n513) );
  NOR2_X1 U604 ( .A1(G902), .A2(n724), .ZN(n485) );
  XNOR2_X1 U605 ( .A(KEYINPUT67), .B(G469), .ZN(n484) );
  INV_X1 U606 ( .A(n626), .ZN(n687) );
  XOR2_X1 U607 ( .A(n486), .B(n509), .Z(n488) );
  NAND2_X1 U608 ( .A1(G217), .A2(n550), .ZN(n487) );
  XNOR2_X1 U609 ( .A(n488), .B(n487), .ZN(n492) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n490) );
  XNOR2_X1 U611 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U612 ( .A(n492), .B(n491), .Z(n494) );
  XNOR2_X1 U613 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n493) );
  XNOR2_X1 U614 ( .A(n494), .B(n493), .ZN(n727) );
  NOR2_X1 U615 ( .A1(G902), .A2(n727), .ZN(n495) );
  XNOR2_X1 U616 ( .A(G478), .B(n495), .ZN(n574) );
  XNOR2_X1 U617 ( .A(KEYINPUT10), .B(n512), .ZN(n555) );
  XOR2_X1 U618 ( .A(G122), .B(G104), .Z(n507) );
  XOR2_X1 U619 ( .A(G140), .B(KEYINPUT11), .Z(n498) );
  XNOR2_X1 U620 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U621 ( .A1(G214), .A2(n537), .ZN(n500) );
  NOR2_X1 U622 ( .A1(G902), .A2(n642), .ZN(n502) );
  XNOR2_X1 U623 ( .A(KEYINPUT92), .B(KEYINPUT13), .ZN(n501) );
  NAND2_X1 U624 ( .A1(G234), .A2(n637), .ZN(n503) );
  XNOR2_X1 U625 ( .A(KEYINPUT20), .B(n503), .ZN(n556) );
  NAND2_X1 U626 ( .A1(n556), .A2(G221), .ZN(n504) );
  XNOR2_X1 U627 ( .A(n504), .B(KEYINPUT21), .ZN(n683) );
  INV_X1 U628 ( .A(n683), .ZN(n505) );
  XOR2_X1 U629 ( .A(KEYINPUT16), .B(n507), .Z(n511) );
  XNOR2_X1 U630 ( .A(KEYINPUT3), .B(G119), .ZN(n508) );
  XNOR2_X1 U631 ( .A(n479), .B(n508), .ZN(n536) );
  XNOR2_X1 U632 ( .A(n536), .B(n509), .ZN(n510) );
  INV_X1 U633 ( .A(n512), .ZN(n514) );
  XNOR2_X1 U634 ( .A(n514), .B(n513), .ZN(n515) );
  NAND2_X1 U635 ( .A1(G224), .A2(n730), .ZN(n516) );
  XNOR2_X1 U636 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U637 ( .A(n518), .B(KEYINPUT73), .Z(n521) );
  XNOR2_X1 U638 ( .A(KEYINPUT4), .B(n519), .ZN(n520) );
  XNOR2_X1 U639 ( .A(n521), .B(n520), .ZN(n522) );
  NAND2_X1 U640 ( .A1(n644), .A2(n637), .ZN(n526) );
  NAND2_X1 U641 ( .A1(n523), .A2(G210), .ZN(n524) );
  NOR2_X1 U642 ( .A1(G898), .A2(n730), .ZN(n737) );
  XNOR2_X1 U643 ( .A(n528), .B(KEYINPUT14), .ZN(n530) );
  NAND2_X1 U644 ( .A1(G902), .A2(n530), .ZN(n584) );
  INV_X1 U645 ( .A(n584), .ZN(n529) );
  NAND2_X1 U646 ( .A1(n737), .A2(n529), .ZN(n532) );
  NAND2_X1 U647 ( .A1(G952), .A2(n530), .ZN(n531) );
  XOR2_X1 U648 ( .A(KEYINPUT86), .B(n531), .Z(n713) );
  NAND2_X1 U649 ( .A1(n730), .A2(n713), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n532), .A2(n587), .ZN(n533) );
  NAND2_X1 U651 ( .A1(n537), .A2(G210), .ZN(n538) );
  XNOR2_X1 U652 ( .A(n539), .B(n538), .ZN(n543) );
  NAND2_X1 U653 ( .A1(G221), .A2(n550), .ZN(n551) );
  XNOR2_X1 U654 ( .A(n555), .B(n554), .ZN(n740) );
  AND2_X1 U655 ( .A1(G217), .A2(n556), .ZN(n558) );
  XNOR2_X1 U656 ( .A(KEYINPUT88), .B(KEYINPUT25), .ZN(n557) );
  NAND2_X1 U657 ( .A1(n561), .A2(n684), .ZN(n562) );
  NOR2_X1 U658 ( .A1(n687), .A2(n562), .ZN(n660) );
  INV_X1 U659 ( .A(n684), .ZN(n583) );
  NOR2_X1 U660 ( .A1(n660), .A2(n755), .ZN(n564) );
  NOR2_X1 U661 ( .A1(n574), .A2(n572), .ZN(n565) );
  INV_X1 U662 ( .A(n566), .ZN(n577) );
  XOR2_X1 U663 ( .A(KEYINPUT96), .B(KEYINPUT33), .Z(n567) );
  XNOR2_X1 U664 ( .A(n568), .B(KEYINPUT34), .ZN(n569) );
  NOR2_X1 U665 ( .A1(n684), .A2(n570), .ZN(n571) );
  NAND2_X1 U666 ( .A1(n626), .A2(n571), .ZN(n652) );
  INV_X1 U667 ( .A(n572), .ZN(n573) );
  NAND2_X1 U668 ( .A1(n574), .A2(n573), .ZN(n618) );
  INV_X1 U669 ( .A(n618), .ZN(n668) );
  NOR2_X1 U670 ( .A1(n574), .A2(n573), .ZN(n670) );
  NOR2_X1 U671 ( .A1(n668), .A2(n670), .ZN(n704) );
  NAND2_X1 U672 ( .A1(n691), .A2(n575), .ZN(n694) );
  XOR2_X1 U673 ( .A(KEYINPUT31), .B(n576), .Z(n671) );
  NOR2_X1 U674 ( .A1(n577), .A2(n608), .ZN(n578) );
  INV_X1 U675 ( .A(KEYINPUT45), .ZN(n580) );
  NOR2_X1 U676 ( .A1(n704), .A2(KEYINPUT47), .ZN(n582) );
  XNOR2_X1 U677 ( .A(KEYINPUT70), .B(n582), .ZN(n594) );
  NOR2_X1 U678 ( .A1(n583), .A2(n683), .ZN(n588) );
  NOR2_X1 U679 ( .A1(G900), .A2(n584), .ZN(n585) );
  NAND2_X1 U680 ( .A1(G953), .A2(n585), .ZN(n586) );
  NAND2_X1 U681 ( .A1(n587), .A2(n586), .ZN(n609) );
  AND2_X1 U682 ( .A1(n588), .A2(n609), .ZN(n596) );
  NAND2_X1 U683 ( .A1(n596), .A2(n605), .ZN(n589) );
  INV_X1 U684 ( .A(n591), .ZN(n592) );
  XNOR2_X1 U685 ( .A(n593), .B(KEYINPUT74), .ZN(n603) );
  BUF_X2 U686 ( .A(n595), .Z(n613) );
  INV_X1 U687 ( .A(n613), .ZN(n629) );
  AND2_X1 U688 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U689 ( .A(KEYINPUT36), .B(KEYINPUT106), .ZN(n599) );
  XNOR2_X1 U690 ( .A(n600), .B(n599), .ZN(n601) );
  INV_X1 U691 ( .A(n704), .ZN(n602) );
  NAND2_X1 U692 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U693 ( .A1(n604), .A2(KEYINPUT47), .ZN(n612) );
  XOR2_X1 U694 ( .A(KEYINPUT30), .B(KEYINPUT101), .Z(n607) );
  XNOR2_X1 U695 ( .A(n607), .B(n606), .ZN(n616) );
  XOR2_X1 U696 ( .A(KEYINPUT82), .B(KEYINPUT39), .Z(n617) );
  INV_X1 U697 ( .A(KEYINPUT38), .ZN(n614) );
  XNOR2_X1 U698 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n619) );
  XNOR2_X1 U699 ( .A(n620), .B(n619), .ZN(n753) );
  NOR2_X1 U700 ( .A1(n698), .A2(n622), .ZN(n623) );
  XNOR2_X1 U701 ( .A(KEYINPUT99), .B(n625), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT43), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U705 ( .A(KEYINPUT100), .B(n631), .ZN(n754) );
  INV_X1 U706 ( .A(n670), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n676) );
  INV_X1 U708 ( .A(n676), .ZN(n634) );
  AND2_X1 U709 ( .A1(n754), .A2(n634), .ZN(n639) );
  INV_X1 U710 ( .A(KEYINPUT2), .ZN(n636) );
  XOR2_X1 U711 ( .A(KEYINPUT79), .B(n637), .Z(n635) );
  INV_X1 U712 ( .A(n637), .ZN(n638) );
  AND2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n721), .A2(G475), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n721), .A2(G210), .ZN(n647) );
  INV_X1 U716 ( .A(n644), .ZN(n646) );
  XOR2_X1 U717 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n645) );
  NAND2_X1 U718 ( .A1(n721), .A2(G472), .ZN(n649) );
  NAND2_X1 U719 ( .A1(G217), .A2(n721), .ZN(n651) );
  XNOR2_X1 U720 ( .A(G101), .B(n652), .ZN(G3) );
  NAND2_X1 U721 ( .A1(n657), .A2(n668), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(G104), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n655) );
  XNOR2_X1 U724 ( .A(G107), .B(KEYINPUT108), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U726 ( .A(KEYINPUT26), .B(n656), .Z(n659) );
  NAND2_X1 U727 ( .A1(n657), .A2(n670), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(G9) );
  XOR2_X1 U729 ( .A(G110), .B(n660), .Z(G12) );
  XOR2_X1 U730 ( .A(KEYINPUT29), .B(KEYINPUT110), .Z(n662) );
  NAND2_X1 U731 ( .A1(n670), .A2(n603), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U733 ( .A(G128), .B(n663), .ZN(G30) );
  XNOR2_X1 U734 ( .A(n664), .B(G143), .ZN(G45) );
  XOR2_X1 U735 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n666) );
  NAND2_X1 U736 ( .A1(n668), .A2(n603), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U738 ( .A(G146), .B(n667), .ZN(G48) );
  NAND2_X1 U739 ( .A1(n671), .A2(n668), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n669), .B(G113), .ZN(G15) );
  XOR2_X1 U741 ( .A(G116), .B(KEYINPUT113), .Z(n673) );
  NAND2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U743 ( .A(n673), .B(n672), .ZN(G18) );
  XOR2_X1 U744 ( .A(G125), .B(KEYINPUT37), .Z(n674) );
  XNOR2_X1 U745 ( .A(n675), .B(n674), .ZN(G27) );
  XOR2_X1 U746 ( .A(G134), .B(n676), .Z(G36) );
  XOR2_X1 U747 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n677) );
  XNOR2_X1 U748 ( .A(KEYINPUT53), .B(n677), .ZN(n720) );
  XNOR2_X1 U749 ( .A(n679), .B(KEYINPUT77), .ZN(n680) );
  NOR2_X1 U750 ( .A1(n709), .A2(n698), .ZN(n682) );
  NOR2_X1 U751 ( .A1(G953), .A2(n682), .ZN(n716) );
  NAND2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U753 ( .A(KEYINPUT49), .B(n685), .Z(n686) );
  XNOR2_X1 U754 ( .A(n686), .B(KEYINPUT114), .ZN(n693) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n689), .B(KEYINPUT50), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U760 ( .A(KEYINPUT51), .B(n696), .ZN(n697) );
  NOR2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n711) );
  NOR2_X1 U762 ( .A1(n621), .A2(n699), .ZN(n700) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U764 ( .A(KEYINPUT115), .B(n702), .Z(n707) );
  NOR2_X1 U765 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U766 ( .A(KEYINPUT116), .B(n705), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U768 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U770 ( .A(KEYINPUT52), .B(n712), .Z(n714) );
  NAND2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U772 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U773 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n720), .B(n719), .ZN(G75) );
  NAND2_X1 U775 ( .A1(n721), .A2(G469), .ZN(n725) );
  XOR2_X1 U776 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n723) );
  XNOR2_X1 U777 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n722) );
  NAND2_X1 U778 ( .A1(G478), .A2(n721), .ZN(n726) );
  XNOR2_X1 U779 ( .A(n726), .B(n727), .ZN(n728) );
  NOR2_X1 U780 ( .A1(n729), .A2(n728), .ZN(G63) );
  NAND2_X1 U781 ( .A1(n730), .A2(n371), .ZN(n734) );
  NAND2_X1 U782 ( .A1(G953), .A2(G224), .ZN(n731) );
  XNOR2_X1 U783 ( .A(KEYINPUT61), .B(n731), .ZN(n732) );
  NAND2_X1 U784 ( .A1(n732), .A2(G898), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n734), .A2(n733), .ZN(n739) );
  XNOR2_X1 U786 ( .A(n735), .B(G110), .ZN(n736) );
  NOR2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(G69) );
  XNOR2_X1 U789 ( .A(n741), .B(n740), .ZN(n746) );
  XNOR2_X1 U790 ( .A(n742), .B(KEYINPUT124), .ZN(n743) );
  XNOR2_X1 U791 ( .A(n746), .B(n743), .ZN(n744) );
  NOR2_X1 U792 ( .A1(G953), .A2(n744), .ZN(n745) );
  XNOR2_X1 U793 ( .A(KEYINPUT125), .B(n745), .ZN(n751) );
  XNOR2_X1 U794 ( .A(G227), .B(n746), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(G953), .ZN(n749) );
  XNOR2_X1 U797 ( .A(KEYINPUT126), .B(n749), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n751), .A2(n750), .ZN(G72) );
  XNOR2_X1 U799 ( .A(n752), .B(G122), .ZN(G24) );
  XOR2_X1 U800 ( .A(n753), .B(G131), .Z(G33) );
  XNOR2_X1 U801 ( .A(G140), .B(n754), .ZN(G42) );
  XOR2_X1 U802 ( .A(n755), .B(G119), .Z(G21) );
  XOR2_X1 U803 ( .A(G137), .B(n756), .Z(G39) );
endmodule

