

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739;

  NOR2_X1 U368 ( .A1(n624), .A2(n592), .ZN(n411) );
  XNOR2_X1 U369 ( .A(n397), .B(n385), .ZN(n602) );
  XNOR2_X1 U370 ( .A(n595), .B(n594), .ZN(n638) );
  NOR2_X1 U371 ( .A1(n659), .A2(n658), .ZN(n664) );
  NOR2_X1 U372 ( .A1(G902), .A2(n688), .ZN(n534) );
  NOR2_X1 U373 ( .A1(n374), .A2(n373), .ZN(n372) );
  NOR2_X1 U374 ( .A1(n382), .A2(n377), .ZN(n373) );
  AND2_X1 U375 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U376 ( .A(n531), .B(n346), .ZN(n532) );
  XNOR2_X1 U377 ( .A(n416), .B(KEYINPUT70), .ZN(n513) );
  INV_X1 U378 ( .A(G953), .ZN(n725) );
  INV_X1 U379 ( .A(n530), .ZN(n346) );
  XNOR2_X2 U380 ( .A(n722), .B(G101), .ZN(n531) );
  XNOR2_X2 U381 ( .A(n359), .B(n358), .ZN(n709) );
  XNOR2_X2 U382 ( .A(n531), .B(n704), .ZN(n465) );
  NOR2_X1 U383 ( .A1(n737), .A2(n736), .ZN(n406) );
  XNOR2_X2 U384 ( .A(KEYINPUT69), .B(G131), .ZN(n416) );
  XNOR2_X2 U385 ( .A(n504), .B(n450), .ZN(n722) );
  XNOR2_X1 U386 ( .A(n561), .B(n404), .ZN(n659) );
  XNOR2_X1 U387 ( .A(n499), .B(n498), .ZN(n641) );
  AND2_X1 U388 ( .A1(n412), .A2(n641), .ZN(n624) );
  XNOR2_X1 U389 ( .A(n388), .B(n387), .ZN(n737) );
  AND2_X1 U390 ( .A1(n553), .A2(n562), .ZN(n351) );
  NOR2_X1 U391 ( .A1(n562), .A2(n553), .ZN(n632) );
  OR2_X1 U392 ( .A1(n641), .A2(n574), .ZN(n648) );
  OR2_X1 U393 ( .A1(n679), .A2(n381), .ZN(n380) );
  XNOR2_X1 U394 ( .A(n528), .B(n529), .ZN(n719) );
  XNOR2_X1 U395 ( .A(n513), .B(n415), .ZN(n529) );
  BUF_X1 U396 ( .A(n581), .Z(n347) );
  XNOR2_X1 U397 ( .A(n348), .B(n719), .ZN(n533) );
  XOR2_X1 U398 ( .A(n527), .B(n526), .Z(n348) );
  NAND2_X1 U399 ( .A1(n366), .A2(n349), .ZN(n449) );
  XOR2_X1 U400 ( .A(n590), .B(KEYINPUT81), .Z(n349) );
  BUF_X2 U401 ( .A(n606), .Z(n397) );
  XNOR2_X1 U402 ( .A(n418), .B(G146), .ZN(n481) );
  INV_X1 U403 ( .A(G125), .ZN(n418) );
  OR2_X1 U404 ( .A1(n469), .A2(G902), .ZN(n431) );
  NAND2_X1 U405 ( .A1(n554), .A2(n378), .ZN(n377) );
  XNOR2_X1 U406 ( .A(KEYINPUT99), .B(n480), .ZN(n642) );
  INV_X1 U407 ( .A(KEYINPUT44), .ZN(n598) );
  NOR2_X1 U408 ( .A1(n561), .A2(n658), .ZN(n438) );
  OR2_X2 U409 ( .A1(n647), .A2(n648), .ZN(n414) );
  XOR2_X1 U410 ( .A(G116), .B(G122), .Z(n508) );
  XNOR2_X1 U411 ( .A(n516), .B(n421), .ZN(n691) );
  XNOR2_X1 U412 ( .A(n424), .B(n422), .ZN(n421) );
  XNOR2_X1 U413 ( .A(n519), .B(n423), .ZN(n422) );
  AND2_X1 U414 ( .A1(n355), .A2(n599), .ZN(n522) );
  NOR2_X1 U415 ( .A1(G902), .A2(G237), .ZN(n467) );
  INV_X1 U416 ( .A(KEYINPUT19), .ZN(n378) );
  NOR2_X1 U417 ( .A1(n351), .A2(n632), .ZN(n662) );
  INV_X1 U418 ( .A(KEYINPUT106), .ZN(n413) );
  XNOR2_X1 U419 ( .A(n478), .B(n477), .ZN(n494) );
  XNOR2_X1 U420 ( .A(KEYINPUT20), .B(KEYINPUT98), .ZN(n477) );
  NOR2_X1 U421 ( .A1(G953), .A2(G237), .ZN(n454) );
  XOR2_X1 U422 ( .A(G113), .B(G104), .Z(n517) );
  XNOR2_X1 U423 ( .A(KEYINPUT87), .B(KEYINPUT8), .ZN(n486) );
  XNOR2_X1 U424 ( .A(n460), .B(n402), .ZN(n530) );
  INV_X1 U425 ( .A(KEYINPUT78), .ZN(n402) );
  XNOR2_X1 U426 ( .A(G110), .B(G107), .ZN(n460) );
  XNOR2_X1 U427 ( .A(G110), .B(KEYINPUT96), .ZN(n488) );
  XNOR2_X1 U428 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n483) );
  XNOR2_X1 U429 ( .A(n481), .B(n417), .ZN(n718) );
  INV_X1 U430 ( .A(KEYINPUT10), .ZN(n417) );
  XNOR2_X1 U431 ( .A(G134), .B(G107), .ZN(n501) );
  XOR2_X1 U432 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n502) );
  XNOR2_X1 U433 ( .A(n465), .B(n464), .ZN(n679) );
  XNOR2_X1 U434 ( .A(n705), .B(n444), .ZN(n464) );
  XNOR2_X1 U435 ( .A(n462), .B(n463), .ZN(n444) );
  AND2_X1 U436 ( .A1(n393), .A2(n392), .ZN(n565) );
  XNOR2_X1 U437 ( .A(n564), .B(KEYINPUT41), .ZN(n656) );
  XNOR2_X1 U438 ( .A(n428), .B(n427), .ZN(n572) );
  INV_X1 U439 ( .A(KEYINPUT39), .ZN(n427) );
  NOR2_X1 U440 ( .A1(n566), .A2(n659), .ZN(n428) );
  AND2_X1 U441 ( .A1(n438), .A2(n439), .ZN(n437) );
  OR2_X1 U442 ( .A1(n525), .A2(n439), .ZN(n434) );
  NAND2_X1 U443 ( .A1(n436), .A2(KEYINPUT36), .ZN(n435) );
  BUF_X1 U444 ( .A(n645), .Z(n396) );
  XNOR2_X1 U445 ( .A(G478), .B(n510), .ZN(n553) );
  XNOR2_X1 U446 ( .A(n521), .B(n520), .ZN(n562) );
  XNOR2_X1 U447 ( .A(n497), .B(n496), .ZN(n498) );
  NOR2_X1 U448 ( .A1(G902), .A2(n701), .ZN(n499) );
  BUF_X1 U449 ( .A(n647), .Z(n386) );
  NAND2_X1 U450 ( .A1(n364), .A2(n362), .ZN(n611) );
  INV_X1 U451 ( .A(G472), .ZN(n363) );
  NOR2_X1 U452 ( .A1(G952), .A2(n725), .ZN(n703) );
  NOR2_X1 U453 ( .A1(n677), .A2(G953), .ZN(n678) );
  AND2_X1 U454 ( .A1(n551), .A2(n552), .ZN(n389) );
  NAND2_X1 U455 ( .A1(n662), .A2(KEYINPUT47), .ZN(n549) );
  XNOR2_X1 U456 ( .A(G116), .B(KEYINPUT5), .ZN(n443) );
  XNOR2_X1 U457 ( .A(G137), .B(G113), .ZN(n453) );
  INV_X1 U458 ( .A(KEYINPUT46), .ZN(n405) );
  NAND2_X1 U459 ( .A1(n379), .A2(n376), .ZN(n375) );
  XNOR2_X1 U460 ( .A(n442), .B(n440), .ZN(n455) );
  XNOR2_X1 U461 ( .A(n441), .B(G146), .ZN(n440) );
  XNOR2_X1 U462 ( .A(n453), .B(n443), .ZN(n442) );
  INV_X1 U463 ( .A(KEYINPUT101), .ZN(n441) );
  INV_X1 U464 ( .A(G134), .ZN(n415) );
  XOR2_X1 U465 ( .A(KEYINPUT65), .B(KEYINPUT4), .Z(n450) );
  XNOR2_X1 U466 ( .A(G137), .B(G140), .ZN(n528) );
  INV_X1 U467 ( .A(G140), .ZN(n423) );
  XNOR2_X1 U468 ( .A(n518), .B(n515), .ZN(n424) );
  XOR2_X1 U469 ( .A(G146), .B(G104), .Z(n527) );
  XNOR2_X1 U470 ( .A(n481), .B(n461), .ZN(n462) );
  OR2_X1 U471 ( .A1(n468), .A2(n466), .ZN(n381) );
  NAND2_X1 U472 ( .A1(n468), .A2(n466), .ZN(n383) );
  NAND2_X1 U473 ( .A1(n679), .A2(n468), .ZN(n384) );
  INV_X1 U474 ( .A(KEYINPUT38), .ZN(n404) );
  INV_X1 U475 ( .A(n557), .ZN(n395) );
  INV_X1 U476 ( .A(n438), .ZN(n436) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n593) );
  XNOR2_X1 U478 ( .A(KEYINPUT0), .B(KEYINPUT68), .ZN(n582) );
  NOR2_X1 U479 ( .A1(n563), .A2(n562), .ZN(n660) );
  XNOR2_X1 U480 ( .A(n495), .B(KEYINPUT97), .ZN(n497) );
  XOR2_X1 U481 ( .A(G119), .B(KEYINPUT3), .Z(n452) );
  XNOR2_X1 U482 ( .A(n445), .B(n458), .ZN(n705) );
  XNOR2_X1 U483 ( .A(n530), .B(n459), .ZN(n445) );
  XOR2_X1 U484 ( .A(KEYINPUT16), .B(KEYINPUT75), .Z(n459) );
  INV_X1 U485 ( .A(n414), .ZN(n605) );
  INV_X1 U486 ( .A(KEYINPUT94), .ZN(n385) );
  XNOR2_X1 U487 ( .A(n493), .B(n492), .ZN(n701) );
  XNOR2_X1 U488 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U489 ( .A(n507), .B(n390), .ZN(n509) );
  XNOR2_X1 U490 ( .A(n506), .B(KEYINPUT7), .ZN(n390) );
  XNOR2_X1 U491 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U492 ( .A(n679), .B(n680), .ZN(n681) );
  INV_X1 U493 ( .A(KEYINPUT42), .ZN(n387) );
  NAND2_X1 U494 ( .A1(n656), .A2(n565), .ZN(n388) );
  XNOR2_X1 U495 ( .A(n426), .B(n425), .ZN(n736) );
  INV_X1 U496 ( .A(KEYINPUT40), .ZN(n425) );
  AND2_X1 U497 ( .A1(n525), .A2(n437), .ZN(n432) );
  INV_X1 U498 ( .A(KEYINPUT35), .ZN(n407) );
  INV_X1 U499 ( .A(n597), .ZN(n409) );
  XNOR2_X1 U500 ( .A(KEYINPUT32), .B(KEYINPUT66), .ZN(n448) );
  NOR2_X1 U501 ( .A1(n597), .A2(n558), .ZN(n627) );
  XNOR2_X1 U502 ( .A(n369), .B(KEYINPUT67), .ZN(n412) );
  OR2_X1 U503 ( .A1(n591), .A2(n367), .ZN(n369) );
  NAND2_X1 U504 ( .A1(n386), .A2(n368), .ZN(n367) );
  NOR2_X1 U505 ( .A1(n613), .A2(n703), .ZN(n615) );
  XNOR2_X1 U506 ( .A(n686), .B(n400), .ZN(n689) );
  XNOR2_X1 U507 ( .A(n688), .B(n687), .ZN(n400) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(G75) );
  XNOR2_X1 U509 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n446) );
  NAND2_X1 U510 ( .A1(n640), .A2(n353), .ZN(n447) );
  OR2_X1 U511 ( .A1(n554), .A2(n378), .ZN(n350) );
  AND2_X1 U512 ( .A1(n366), .A2(n386), .ZN(n352) );
  AND2_X1 U513 ( .A1(n678), .A2(n639), .ZN(n353) );
  OR2_X1 U514 ( .A1(n662), .A2(n608), .ZN(n354) );
  AND2_X1 U515 ( .A1(n542), .A2(n351), .ZN(n355) );
  AND2_X1 U516 ( .A1(n546), .A2(n435), .ZN(n356) );
  INV_X1 U517 ( .A(KEYINPUT36), .ZN(n439) );
  XOR2_X1 U518 ( .A(KEYINPUT34), .B(KEYINPUT74), .Z(n357) );
  XOR2_X1 U519 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n358) );
  NAND2_X1 U520 ( .A1(n572), .A2(n351), .ZN(n426) );
  NAND2_X1 U521 ( .A1(n399), .A2(n556), .ZN(n566) );
  NOR2_X1 U522 ( .A1(n683), .A2(n703), .ZN(n685) );
  NOR2_X1 U523 ( .A1(n694), .A2(n703), .ZN(n696) );
  XNOR2_X1 U524 ( .A(n361), .B(n598), .ZN(n360) );
  NAND2_X1 U525 ( .A1(n360), .A2(n609), .ZN(n359) );
  NAND2_X1 U526 ( .A1(n411), .A2(n735), .ZN(n361) );
  NOR2_X4 U527 ( .A1(n637), .A2(n610), .ZN(n365) );
  NOR2_X1 U528 ( .A1(n610), .A2(n363), .ZN(n362) );
  INV_X1 U529 ( .A(n637), .ZN(n364) );
  NAND2_X1 U530 ( .A1(n365), .A2(G210), .ZN(n682) );
  NAND2_X1 U531 ( .A1(n365), .A2(G475), .ZN(n693) );
  NAND2_X1 U532 ( .A1(n365), .A2(G478), .ZN(n697) );
  NAND2_X1 U533 ( .A1(n365), .A2(G217), .ZN(n700) );
  NAND2_X1 U534 ( .A1(n365), .A2(G469), .ZN(n686) );
  INV_X1 U535 ( .A(n591), .ZN(n366) );
  INV_X1 U536 ( .A(n396), .ZN(n368) );
  NAND2_X1 U537 ( .A1(n382), .A2(n380), .ZN(n541) );
  NAND2_X1 U538 ( .A1(n372), .A2(n370), .ZN(n581) );
  NAND2_X1 U539 ( .A1(n371), .A2(n382), .ZN(n370) );
  AND2_X1 U540 ( .A1(n380), .A2(KEYINPUT19), .ZN(n371) );
  NAND2_X1 U541 ( .A1(n375), .A2(n350), .ZN(n374) );
  INV_X1 U542 ( .A(n377), .ZN(n376) );
  INV_X1 U543 ( .A(n380), .ZN(n379) );
  NOR2_X1 U544 ( .A1(n647), .A2(n586), .ZN(n587) );
  XNOR2_X2 U545 ( .A(n555), .B(KEYINPUT1), .ZN(n647) );
  XNOR2_X1 U546 ( .A(n543), .B(KEYINPUT28), .ZN(n393) );
  NOR2_X1 U547 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U548 ( .A(n641), .ZN(n586) );
  NAND2_X1 U549 ( .A1(n394), .A2(n641), .ZN(n500) );
  NAND2_X1 U550 ( .A1(n420), .A2(n389), .ZN(n391) );
  XNOR2_X1 U551 ( .A(n401), .B(KEYINPUT22), .ZN(n591) );
  NAND2_X1 U552 ( .A1(n638), .A2(n602), .ZN(n596) );
  XNOR2_X1 U553 ( .A(n583), .B(n582), .ZN(n606) );
  AND2_X1 U554 ( .A1(n603), .A2(n557), .ZN(n399) );
  XNOR2_X1 U555 ( .A(n391), .B(KEYINPUT84), .ZN(n419) );
  INV_X1 U556 ( .A(n555), .ZN(n392) );
  NOR2_X1 U557 ( .A1(n642), .A2(n395), .ZN(n394) );
  NAND2_X1 U558 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U559 ( .A1(n584), .A2(n585), .ZN(n401) );
  NOR2_X2 U560 ( .A1(n709), .A2(n717), .ZN(n403) );
  XNOR2_X2 U561 ( .A(n398), .B(G143), .ZN(n504) );
  XNOR2_X2 U562 ( .A(G128), .B(KEYINPUT83), .ZN(n398) );
  XNOR2_X2 U563 ( .A(n403), .B(KEYINPUT2), .ZN(n637) );
  XNOR2_X1 U564 ( .A(n406), .B(n405), .ZN(n567) );
  XNOR2_X2 U565 ( .A(n408), .B(n407), .ZN(n735) );
  NAND2_X1 U566 ( .A1(n410), .A2(n409), .ZN(n408) );
  XNOR2_X1 U567 ( .A(n596), .B(n357), .ZN(n410) );
  XNOR2_X2 U568 ( .A(n534), .B(n535), .ZN(n555) );
  NOR2_X1 U569 ( .A1(n732), .A2(n419), .ZN(n559) );
  INV_X1 U570 ( .A(n627), .ZN(n420) );
  AND2_X1 U571 ( .A1(n660), .A2(n575), .ZN(n585) );
  XNOR2_X1 U572 ( .A(n430), .B(n429), .ZN(n556) );
  INV_X1 U573 ( .A(KEYINPUT30), .ZN(n429) );
  NAND2_X1 U574 ( .A1(n645), .A2(n554), .ZN(n430) );
  XNOR2_X2 U575 ( .A(n431), .B(G472), .ZN(n645) );
  NOR2_X2 U576 ( .A1(n433), .A2(n432), .ZN(n547) );
  NAND2_X1 U577 ( .A1(n434), .A2(n356), .ZN(n433) );
  NAND2_X1 U578 ( .A1(n525), .A2(n554), .ZN(n545) );
  XNOR2_X2 U579 ( .A(n449), .B(n448), .ZN(n734) );
  INV_X1 U580 ( .A(n541), .ZN(n561) );
  XNOR2_X1 U581 ( .A(n682), .B(n681), .ZN(n683) );
  INV_X1 U582 ( .A(n606), .ZN(n584) );
  AND2_X1 U583 ( .A1(G210), .A2(n514), .ZN(n451) );
  INV_X1 U584 ( .A(KEYINPUT48), .ZN(n569) );
  INV_X1 U585 ( .A(n574), .ZN(n575) );
  XNOR2_X1 U586 ( .A(n455), .B(n451), .ZN(n456) );
  XNOR2_X1 U587 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U588 ( .A(KEYINPUT90), .B(KEYINPUT33), .ZN(n594) );
  XNOR2_X1 U589 ( .A(n456), .B(n529), .ZN(n457) );
  XNOR2_X1 U590 ( .A(n485), .B(n718), .ZN(n493) );
  XNOR2_X1 U591 ( .A(n693), .B(n692), .ZN(n694) );
  INV_X1 U592 ( .A(KEYINPUT63), .ZN(n614) );
  XNOR2_X1 U593 ( .A(KEYINPUT73), .B(n452), .ZN(n704) );
  XOR2_X1 U594 ( .A(KEYINPUT79), .B(n454), .Z(n514) );
  XNOR2_X1 U595 ( .A(n465), .B(n457), .ZN(n469) );
  XNOR2_X1 U596 ( .A(n469), .B(KEYINPUT62), .ZN(n612) );
  XNOR2_X2 U597 ( .A(G902), .B(KEYINPUT15), .ZN(n610) );
  INV_X1 U598 ( .A(n610), .ZN(n466) );
  XNOR2_X1 U599 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n463) );
  XNOR2_X1 U600 ( .A(n508), .B(n517), .ZN(n458) );
  AND2_X1 U601 ( .A1(G224), .A2(n725), .ZN(n461) );
  XNOR2_X1 U602 ( .A(n467), .B(KEYINPUT77), .ZN(n523) );
  AND2_X1 U603 ( .A1(G210), .A2(n523), .ZN(n468) );
  XOR2_X2 U604 ( .A(KEYINPUT6), .B(n645), .Z(n599) );
  NAND2_X1 U605 ( .A1(G234), .A2(G237), .ZN(n470) );
  XNOR2_X1 U606 ( .A(n470), .B(KEYINPUT14), .ZN(n473) );
  NAND2_X1 U607 ( .A1(G902), .A2(n473), .ZN(n576) );
  NOR2_X1 U608 ( .A1(G900), .A2(n576), .ZN(n471) );
  NAND2_X1 U609 ( .A1(G953), .A2(n471), .ZN(n472) );
  XOR2_X1 U610 ( .A(KEYINPUT107), .B(n472), .Z(n476) );
  NAND2_X1 U611 ( .A1(G952), .A2(n473), .ZN(n474) );
  XNOR2_X1 U612 ( .A(KEYINPUT92), .B(n474), .ZN(n675) );
  NOR2_X1 U613 ( .A1(n675), .A2(G953), .ZN(n475) );
  XNOR2_X1 U614 ( .A(n475), .B(KEYINPUT93), .ZN(n578) );
  NAND2_X1 U615 ( .A1(n476), .A2(n578), .ZN(n557) );
  NAND2_X1 U616 ( .A1(n610), .A2(G234), .ZN(n478) );
  NAND2_X1 U617 ( .A1(n494), .A2(G221), .ZN(n479) );
  XOR2_X1 U618 ( .A(KEYINPUT21), .B(n479), .Z(n480) );
  XNOR2_X1 U619 ( .A(G128), .B(G119), .ZN(n482) );
  XNOR2_X1 U620 ( .A(n528), .B(n482), .ZN(n484) );
  XNOR2_X1 U621 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U622 ( .A1(n725), .A2(G234), .ZN(n487) );
  XNOR2_X1 U623 ( .A(n487), .B(n486), .ZN(n505) );
  NAND2_X1 U624 ( .A1(n505), .A2(G221), .ZN(n491) );
  XOR2_X1 U625 ( .A(KEYINPUT86), .B(KEYINPUT95), .Z(n489) );
  XNOR2_X1 U626 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U627 ( .A1(n494), .A2(G217), .ZN(n495) );
  XNOR2_X1 U628 ( .A(KEYINPUT25), .B(KEYINPUT80), .ZN(n496) );
  XNOR2_X1 U629 ( .A(KEYINPUT71), .B(n500), .ZN(n542) );
  XNOR2_X1 U630 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U631 ( .A(n504), .B(n503), .Z(n507) );
  NAND2_X1 U632 ( .A1(G217), .A2(n505), .ZN(n506) );
  XOR2_X1 U633 ( .A(n509), .B(n508), .Z(n698) );
  NOR2_X1 U634 ( .A1(G902), .A2(n698), .ZN(n510) );
  XOR2_X1 U635 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n512) );
  XNOR2_X1 U636 ( .A(G122), .B(KEYINPUT102), .ZN(n511) );
  XNOR2_X1 U637 ( .A(n512), .B(n511), .ZN(n519) );
  XOR2_X1 U638 ( .A(n513), .B(n718), .Z(n516) );
  NAND2_X1 U639 ( .A1(G214), .A2(n514), .ZN(n515) );
  XNOR2_X1 U640 ( .A(G143), .B(n517), .ZN(n518) );
  NOR2_X1 U641 ( .A1(G902), .A2(n691), .ZN(n521) );
  XNOR2_X1 U642 ( .A(KEYINPUT13), .B(G475), .ZN(n520) );
  XNOR2_X1 U643 ( .A(n522), .B(KEYINPUT108), .ZN(n525) );
  NAND2_X1 U644 ( .A1(n523), .A2(G214), .ZN(n524) );
  XNOR2_X1 U645 ( .A(KEYINPUT91), .B(n524), .ZN(n658) );
  INV_X1 U646 ( .A(n658), .ZN(n554) );
  XNOR2_X1 U647 ( .A(n545), .B(KEYINPUT109), .ZN(n536) );
  XNOR2_X1 U648 ( .A(KEYINPUT72), .B(G469), .ZN(n535) );
  NAND2_X1 U649 ( .A1(G227), .A2(n725), .ZN(n526) );
  XNOR2_X1 U650 ( .A(n532), .B(n533), .ZN(n688) );
  NAND2_X1 U651 ( .A1(n536), .A2(n386), .ZN(n537) );
  XNOR2_X1 U652 ( .A(n537), .B(KEYINPUT110), .ZN(n538) );
  XOR2_X1 U653 ( .A(KEYINPUT43), .B(n538), .Z(n539) );
  NOR2_X1 U654 ( .A1(n541), .A2(n539), .ZN(n636) );
  NOR2_X1 U655 ( .A1(n662), .A2(KEYINPUT47), .ZN(n540) );
  XNOR2_X1 U656 ( .A(KEYINPUT76), .B(n540), .ZN(n544) );
  AND2_X1 U657 ( .A1(n542), .A2(n645), .ZN(n543) );
  NAND2_X1 U658 ( .A1(n347), .A2(n565), .ZN(n550) );
  INV_X1 U659 ( .A(n550), .ZN(n628) );
  NAND2_X1 U660 ( .A1(n544), .A2(n628), .ZN(n560) );
  INV_X1 U661 ( .A(KEYINPUT111), .ZN(n548) );
  INV_X1 U662 ( .A(n386), .ZN(n546) );
  XNOR2_X1 U663 ( .A(n548), .B(n547), .ZN(n732) );
  XOR2_X1 U664 ( .A(n549), .B(KEYINPUT85), .Z(n552) );
  NAND2_X1 U665 ( .A1(n550), .A2(KEYINPUT47), .ZN(n551) );
  INV_X1 U666 ( .A(n553), .ZN(n563) );
  NAND2_X1 U667 ( .A1(n563), .A2(n562), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n642), .B(KEYINPUT100), .ZN(n574) );
  NOR2_X1 U669 ( .A1(n555), .A2(n648), .ZN(n603) );
  OR2_X1 U670 ( .A1(n561), .A2(n566), .ZN(n558) );
  NAND2_X1 U671 ( .A1(n560), .A2(n559), .ZN(n568) );
  NAND2_X1 U672 ( .A1(n664), .A2(n660), .ZN(n564) );
  NOR2_X1 U673 ( .A1(n568), .A2(n567), .ZN(n570) );
  NOR2_X1 U674 ( .A1(n636), .A2(n571), .ZN(n573) );
  NAND2_X1 U675 ( .A1(n572), .A2(n632), .ZN(n635) );
  NAND2_X1 U676 ( .A1(n573), .A2(n635), .ZN(n717) );
  NOR2_X1 U677 ( .A1(G898), .A2(n725), .ZN(n708) );
  INV_X1 U678 ( .A(n576), .ZN(n577) );
  NAND2_X1 U679 ( .A1(n708), .A2(n577), .ZN(n579) );
  NAND2_X1 U680 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U681 ( .A(n599), .B(KEYINPUT82), .ZN(n589) );
  XNOR2_X1 U682 ( .A(n587), .B(KEYINPUT105), .ZN(n588) );
  INV_X1 U683 ( .A(n734), .ZN(n592) );
  NAND2_X1 U684 ( .A1(n593), .A2(n599), .ZN(n595) );
  NOR2_X1 U685 ( .A1(n641), .A2(n599), .ZN(n600) );
  NAND2_X1 U686 ( .A1(n352), .A2(n600), .ZN(n601) );
  XNOR2_X1 U687 ( .A(KEYINPUT104), .B(n601), .ZN(n739) );
  NAND2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U689 ( .A1(n396), .A2(n604), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n396), .A2(n605), .ZN(n653) );
  NOR2_X1 U691 ( .A1(n397), .A2(n653), .ZN(n607) );
  XOR2_X1 U692 ( .A(KEYINPUT31), .B(n607), .Z(n633) );
  NOR2_X1 U693 ( .A1(n619), .A2(n633), .ZN(n608) );
  AND2_X1 U694 ( .A1(n739), .A2(n354), .ZN(n609) );
  XNOR2_X1 U695 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U696 ( .A(n615), .B(n614), .ZN(G57) );
  XOR2_X1 U697 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n617) );
  NAND2_X1 U698 ( .A1(n619), .A2(n351), .ZN(n616) );
  XNOR2_X1 U699 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U700 ( .A(G104), .B(n618), .ZN(G6) );
  XNOR2_X1 U701 ( .A(G107), .B(KEYINPUT26), .ZN(n623) );
  XOR2_X1 U702 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n621) );
  NAND2_X1 U703 ( .A1(n619), .A2(n632), .ZN(n620) );
  XNOR2_X1 U704 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U705 ( .A(n623), .B(n622), .ZN(G9) );
  XOR2_X1 U706 ( .A(n624), .B(G110), .Z(G12) );
  XOR2_X1 U707 ( .A(G128), .B(KEYINPUT29), .Z(n626) );
  NAND2_X1 U708 ( .A1(n628), .A2(n632), .ZN(n625) );
  XNOR2_X1 U709 ( .A(n626), .B(n625), .ZN(G30) );
  XOR2_X1 U710 ( .A(n627), .B(G143), .Z(G45) );
  XOR2_X1 U711 ( .A(G146), .B(KEYINPUT115), .Z(n630) );
  NAND2_X1 U712 ( .A1(n628), .A2(n351), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n630), .B(n629), .ZN(G48) );
  NAND2_X1 U714 ( .A1(n633), .A2(n351), .ZN(n631) );
  XNOR2_X1 U715 ( .A(n631), .B(G113), .ZN(G15) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U717 ( .A(n634), .B(G116), .ZN(G18) );
  XNOR2_X1 U718 ( .A(G134), .B(n635), .ZN(G36) );
  XOR2_X1 U719 ( .A(G140), .B(n636), .Z(G42) );
  XNOR2_X1 U720 ( .A(n637), .B(KEYINPUT88), .ZN(n640) );
  BUF_X1 U721 ( .A(n638), .Z(n668) );
  NAND2_X1 U722 ( .A1(n668), .A2(n656), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U724 ( .A(KEYINPUT49), .B(n643), .ZN(n644) );
  NOR2_X1 U725 ( .A1(n396), .A2(n644), .ZN(n646) );
  XNOR2_X1 U726 ( .A(n646), .B(KEYINPUT116), .ZN(n652) );
  XOR2_X1 U727 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n650) );
  NAND2_X1 U728 ( .A1(n648), .A2(n386), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U732 ( .A(KEYINPUT51), .B(n655), .Z(n657) );
  NAND2_X1 U733 ( .A1(n657), .A2(n656), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n661) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n666) );
  INV_X1 U736 ( .A(n662), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n667), .B(KEYINPUT118), .ZN(n669) );
  NAND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n672), .B(KEYINPUT119), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n673), .B(KEYINPUT52), .ZN(n674) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n676), .B(KEYINPUT120), .ZN(n677) );
  XOR2_X1 U746 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n680) );
  XOR2_X1 U747 ( .A(KEYINPUT89), .B(KEYINPUT56), .Z(n684) );
  XNOR2_X1 U748 ( .A(n685), .B(n684), .ZN(G51) );
  XOR2_X1 U749 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n687) );
  NOR2_X1 U750 ( .A1(n703), .A2(n689), .ZN(G54) );
  XOR2_X1 U751 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n690) );
  XOR2_X1 U752 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n695) );
  XNOR2_X1 U753 ( .A(n696), .B(n695), .ZN(G60) );
  XNOR2_X1 U754 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U755 ( .A1(n703), .A2(n699), .ZN(G63) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U757 ( .A1(n703), .A2(n702), .ZN(G66) );
  XNOR2_X1 U758 ( .A(n705), .B(n704), .ZN(n706) );
  XOR2_X1 U759 ( .A(G101), .B(n706), .Z(n707) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(n716) );
  OR2_X1 U761 ( .A1(n709), .A2(G953), .ZN(n714) );
  NAND2_X1 U762 ( .A1(G224), .A2(G953), .ZN(n710) );
  XNOR2_X1 U763 ( .A(n710), .B(KEYINPUT124), .ZN(n711) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n711), .ZN(n712) );
  NAND2_X1 U765 ( .A1(G898), .A2(n712), .ZN(n713) );
  NAND2_X1 U766 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U767 ( .A(n716), .B(n715), .ZN(G69) );
  XOR2_X1 U768 ( .A(KEYINPUT126), .B(n717), .Z(n724) );
  XOR2_X1 U769 ( .A(n719), .B(n718), .Z(n720) );
  XNOR2_X1 U770 ( .A(KEYINPUT125), .B(n720), .ZN(n721) );
  XOR2_X1 U771 ( .A(n722), .B(n721), .Z(n727) );
  INV_X1 U772 ( .A(n727), .ZN(n723) );
  XOR2_X1 U773 ( .A(n724), .B(n723), .Z(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n731) );
  XOR2_X1 U775 ( .A(G227), .B(n727), .Z(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G72) );
  XNOR2_X1 U779 ( .A(n732), .B(G125), .ZN(n733) );
  XNOR2_X1 U780 ( .A(n733), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U781 ( .A(n734), .B(G119), .ZN(G21) );
  XNOR2_X1 U782 ( .A(n735), .B(G122), .ZN(G24) );
  XOR2_X1 U783 ( .A(G131), .B(n736), .Z(G33) );
  XNOR2_X1 U784 ( .A(G137), .B(KEYINPUT127), .ZN(n738) );
  XNOR2_X1 U785 ( .A(n738), .B(n737), .ZN(G39) );
  XNOR2_X1 U786 ( .A(G101), .B(n739), .ZN(G3) );
endmodule

