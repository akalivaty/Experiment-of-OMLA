//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT4), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT78), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT78), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G141gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n207), .A3(G148gat), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n204), .A2(G148gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND3_X1   g020(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n222), .A2(new_n223), .A3(new_n212), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G127gat), .ZN(new_n228));
  INV_X1    g027(.A(G127gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G134gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n233));
  INV_X1    g032(.A(G120gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G113gat), .ZN(new_n235));
  INV_X1    g034(.A(G113gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G120gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n203), .B1(new_n226), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n242), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n211), .A2(new_n216), .B1(new_n221), .B2(new_n224), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT4), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n210), .A2(new_n218), .B1(KEYINPUT77), .B2(KEYINPUT2), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT77), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n215), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G155gat), .ZN(new_n252));
  INV_X1    g051(.A(G162gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n249), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n208), .A2(new_n210), .B1(new_n215), .B2(new_n214), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT3), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n217), .A2(new_n260), .A3(new_n225), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n261), .A3(new_n242), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n247), .A2(KEYINPUT5), .A3(new_n248), .A4(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n248), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n242), .A2(new_n258), .A3(new_n257), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n217), .A2(new_n225), .B1(new_n241), .B2(new_n233), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n262), .A2(new_n243), .A3(new_n248), .A4(new_n246), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G1gat), .B(G29gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT0), .ZN(new_n272));
  XNOR2_X1  g071(.A(G57gat), .B(G85gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n263), .A2(new_n270), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n263), .B2(new_n270), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n202), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n276), .A2(new_n277), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n270), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n274), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n283), .A2(KEYINPUT83), .A3(new_n277), .A4(new_n276), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n280), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G226gat), .A2(G233gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT27), .B(G183gat), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(KEYINPUT28), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT70), .A2(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(KEYINPUT70), .A2(G183gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT27), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(G190gat), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n290), .B1(new_n297), .B2(KEYINPUT28), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(G169gat), .ZN(new_n300));
  INV_X1    g099(.A(G176gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT67), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n300), .A2(new_n301), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(KEYINPUT26), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n299), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OR2_X1    g115(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n317), .A2(KEYINPUT23), .A3(new_n300), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n321), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n319), .A2(KEYINPUT65), .A3(new_n320), .A4(new_n322), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT25), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n329), .A2(new_n322), .A3(KEYINPUT25), .A4(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n302), .A2(new_n304), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(KEYINPUT23), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT24), .B1(new_n299), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n334), .B2(new_n299), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n312), .A2(KEYINPUT69), .ZN(new_n337));
  INV_X1    g136(.A(new_n293), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(new_n289), .A3(new_n291), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n312), .A2(KEYINPUT69), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n336), .A2(new_n337), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n333), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n311), .B1(new_n327), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n287), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n310), .A2(new_n299), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT70), .B(G183gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n295), .B1(new_n349), .B2(KEYINPUT27), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n350), .B2(G190gat), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n347), .B1(new_n351), .B2(new_n290), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n300), .A2(KEYINPUT23), .ZN(new_n353));
  AND2_X1   g152(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n322), .A2(new_n320), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n324), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n316), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n326), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n352), .B1(new_n362), .B2(new_n342), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n286), .ZN(new_n364));
  XNOR2_X1  g163(.A(G197gat), .B(G204gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366));
  INV_X1    g165(.A(G211gat), .ZN(new_n367));
  INV_X1    g166(.A(G218gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT74), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G218gat), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n365), .B(new_n366), .C1(new_n372), .C2(KEYINPUT22), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT22), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT74), .B(G218gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n367), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n366), .B1(new_n377), .B2(new_n365), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n346), .A2(new_n364), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n366), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n369), .A2(new_n371), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT22), .B1(new_n382), .B2(G211gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n365), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n373), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n286), .B1(new_n363), .B2(KEYINPUT29), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n344), .A2(new_n287), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT37), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n379), .B1(new_n346), .B2(new_n364), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n386), .A3(new_n388), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT37), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(G8gat), .B(G36gat), .Z(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n390), .A2(new_n394), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT38), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT38), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n390), .A2(new_n403), .A3(new_n394), .A4(new_n400), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n391), .A2(new_n392), .A3(new_n399), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n285), .A2(new_n402), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n265), .A2(new_n266), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT39), .B1(new_n407), .B2(new_n264), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n262), .A2(new_n243), .A3(new_n246), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n264), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n264), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n274), .B1(new_n411), .B2(KEYINPUT39), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n276), .B1(new_n413), .B2(KEYINPUT40), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(KEYINPUT40), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT82), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n417), .A3(KEYINPUT40), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT30), .A4(new_n399), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n400), .B1(new_n380), .B2(new_n389), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G78gat), .B(G106gat), .ZN(new_n426));
  INV_X1    g225(.A(G50gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G22gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT29), .B1(new_n245), .B2(new_n260), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(new_n431), .B2(new_n386), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n385), .B2(new_n373), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n226), .B1(new_n433), .B2(KEYINPUT3), .ZN(new_n434));
  INV_X1    g233(.A(G228gat), .ZN(new_n435));
  INV_X1    g234(.A(G233gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n261), .A2(new_n345), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n379), .A3(KEYINPUT80), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n432), .A2(new_n434), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n441));
  INV_X1    g240(.A(new_n437), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n345), .B1(new_n374), .B2(new_n378), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n260), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n444), .B2(new_n226), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n439), .A4(new_n432), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n438), .A2(new_n379), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n437), .B1(new_n434), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n429), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  AOI211_X1 g251(.A(G22gat), .B(new_n450), .C1(new_n441), .C2(new_n447), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n428), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n431), .A2(new_n430), .A3(new_n386), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT80), .B1(new_n438), .B2(new_n379), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n446), .B1(new_n457), .B2(new_n445), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n451), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(G22gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n448), .A2(new_n429), .A3(new_n451), .ZN(new_n462));
  INV_X1    g261(.A(new_n428), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n454), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n454), .B2(new_n464), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n406), .B(new_n425), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n454), .A2(new_n464), .ZN(new_n469));
  INV_X1    g268(.A(new_n465), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n464), .A3(new_n465), .ZN(new_n472));
  INV_X1    g271(.A(new_n424), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n283), .A2(new_n277), .A3(new_n276), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n281), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n471), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n468), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n360), .A2(new_n361), .B1(new_n341), .B2(new_n333), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n242), .B1(new_n480), .B2(new_n352), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n311), .B(new_n244), .C1(new_n327), .C2(new_n343), .ZN(new_n482));
  NAND2_X1  g281(.A1(G227gat), .A2(G233gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT34), .ZN(new_n485));
  XNOR2_X1  g284(.A(G71gat), .B(G99gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT71), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G15gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n486), .B(KEYINPUT71), .ZN(new_n490));
  INV_X1    g289(.A(G15gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G43gat), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n483), .B1(new_n481), .B2(new_n482), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(KEYINPUT33), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT32), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n482), .ZN(new_n500));
  INV_X1    g299(.A(new_n483), .ZN(new_n501));
  AOI221_X4 g300(.A(new_n497), .B1(new_n494), .B2(KEYINPUT33), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n485), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n362), .A2(new_n342), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n244), .B1(new_n504), .B2(new_n311), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n480), .A2(new_n242), .A3(new_n352), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT32), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n510), .A3(new_n494), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT34), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n484), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n503), .A2(new_n515), .A3(KEYINPUT72), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT72), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n518), .B(new_n485), .C1(new_n499), .C2(new_n502), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n503), .A2(new_n515), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n516), .A2(KEYINPUT73), .A3(new_n517), .A4(new_n519), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n475), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(new_n424), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n528), .B(new_n523), .C1(new_n466), .C2(new_n467), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT35), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n285), .A2(KEYINPUT35), .A3(new_n424), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n519), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n471), .A2(new_n472), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n479), .A2(new_n526), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  OR2_X1    g336(.A1(G43gat), .A2(G50gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(G43gat), .A2(G50gat), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(G29gat), .A2(G36gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT14), .ZN(new_n542));
  INV_X1    g341(.A(G29gat), .ZN(new_n543));
  INV_X1    g342(.A(G36gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n540), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT85), .B(G43gat), .Z(new_n547));
  OAI211_X1 g346(.A(new_n537), .B(new_n539), .C1(new_n547), .C2(G50gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(KEYINPUT86), .B2(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n540), .A2(new_n545), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n546), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT17), .ZN(new_n554));
  XNOR2_X1  g353(.A(G15gat), .B(G22gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT16), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(G1gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(G1gat), .B2(new_n555), .ZN(new_n558));
  INV_X1    g357(.A(G8gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n560), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n553), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n566), .A2(KEYINPUT87), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n567), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n560), .B(new_n553), .Z(new_n570));
  XOR2_X1   g369(.A(new_n562), .B(KEYINPUT13), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G169gat), .B(G197gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT12), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n568), .A2(new_n569), .A3(new_n572), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n536), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT92), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(new_n592), .B2(new_n591), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n590), .ZN(new_n597));
  NAND2_X1  g396(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n591), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n594), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n595), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n589), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G99gat), .B(G106gat), .Z(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  XNOR2_X1  g404(.A(G57gat), .B(G64gat), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G71gat), .B(G78gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  OR2_X1    g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n605), .A2(new_n610), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT10), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n610), .B(KEYINPUT90), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n605), .A3(KEYINPUT10), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G230gat), .ZN(new_n617));
  OAI22_X1  g416(.A1(new_n613), .A2(new_n616), .B1(new_n617), .B2(new_n436), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n611), .A2(new_n612), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n617), .A2(new_n436), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G120gat), .B(G148gat), .Z(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n618), .A2(new_n621), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT99), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(KEYINPUT99), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n610), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(KEYINPUT21), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n563), .B1(new_n614), .B2(KEYINPUT21), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT20), .ZN(new_n642));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT88), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G183gat), .B(G211gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT91), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n645), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n640), .B(new_n648), .Z(new_n649));
  OR2_X1    g448(.A1(new_n605), .A2(KEYINPUT95), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n605), .A2(KEYINPUT95), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n554), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(G232gat), .A2(G233gat), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n605), .A2(new_n553), .B1(KEYINPUT41), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n652), .A2(new_n658), .A3(new_n654), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n653), .A2(KEYINPUT41), .ZN(new_n660));
  XNOR2_X1  g459(.A(G134gat), .B(G162gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n657), .A2(KEYINPUT96), .A3(new_n659), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT96), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n666), .A2(new_n662), .B1(new_n657), .B2(new_n659), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n634), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n585), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n527), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n424), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT100), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(G8gat), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n675), .A2(new_n674), .A3(new_n677), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(G1325gat));
  NAND4_X1  g480(.A1(new_n585), .A2(new_n491), .A3(new_n532), .A4(new_n670), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n671), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n682), .B1(new_n684), .B2(new_n491), .ZN(G1326gat));
  INV_X1    g484(.A(new_n534), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  NOR3_X1   g488(.A1(new_n634), .A2(new_n668), .A3(new_n649), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n585), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(new_n543), .A3(new_n527), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT101), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n535), .A2(new_n530), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n526), .A2(new_n468), .A3(new_n477), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n664), .B2(new_n667), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n666), .A2(new_n662), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n657), .A2(new_n659), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(KEYINPUT102), .A3(new_n663), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n536), .A2(new_n668), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n634), .ZN(new_n711));
  INV_X1    g510(.A(new_n649), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n583), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n527), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n543), .B1(new_n715), .B2(KEYINPUT103), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(KEYINPUT103), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n694), .A2(new_n717), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n691), .A2(new_n544), .A3(new_n424), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT46), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n544), .B1(new_n714), .B2(new_n424), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT104), .ZN(G1329gat));
  NAND2_X1  g522(.A1(new_n714), .A2(new_n683), .ZN(new_n724));
  INV_X1    g523(.A(new_n532), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n547), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n724), .A2(new_n547), .B1(new_n691), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1330gat));
  NAND3_X1  g532(.A1(new_n714), .A2(G50gat), .A3(new_n686), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n691), .A2(new_n686), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(G50gat), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g536(.A1(new_n536), .A2(new_n711), .A3(new_n583), .A4(new_n669), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n527), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n424), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT49), .B(G64gat), .Z(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(G1333gat));
  NAND2_X1  g543(.A1(new_n738), .A2(new_n683), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n725), .A2(G71gat), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n745), .A2(G71gat), .B1(new_n738), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n738), .A2(new_n686), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n649), .A2(new_n583), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n634), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n710), .A2(KEYINPUT107), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n755));
  INV_X1    g554(.A(new_n752), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n709), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n475), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  INV_X1    g560(.A(new_n668), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n683), .A2(new_n478), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n534), .A2(new_n533), .B1(new_n529), .B2(KEYINPUT35), .ZN(new_n764));
  OAI211_X1 g563(.A(KEYINPUT108), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n751), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT108), .B1(new_n697), .B2(new_n762), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n761), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n536), .B2(new_n668), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(KEYINPUT51), .A3(new_n751), .A4(new_n765), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(KEYINPUT109), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n773), .B(new_n761), .C1(new_n766), .C2(new_n767), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n634), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n527), .A2(new_n587), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n760), .B1(new_n775), .B2(new_n776), .ZN(G1336gat));
  NAND2_X1  g576(.A1(new_n768), .A2(new_n771), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n634), .A2(new_n588), .A3(new_n424), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT110), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n753), .A2(new_n473), .A3(new_n757), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n782), .B2(new_n588), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n772), .A2(new_n774), .A3(new_n780), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT111), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n787), .A3(new_n774), .A4(new_n780), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n709), .A2(new_n424), .A3(new_n756), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G92gat), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT112), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  AOI211_X1 g595(.A(new_n796), .B(new_n793), .C1(new_n786), .C2(new_n788), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n784), .B1(new_n795), .B2(new_n797), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n759), .B2(new_n526), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n725), .A2(G99gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n775), .B2(new_n800), .ZN(G1338gat));
  NAND3_X1  g600(.A1(new_n754), .A2(new_n686), .A3(new_n758), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(G106gat), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n711), .A2(G106gat), .A3(new_n534), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n802), .A2(new_n803), .B1(new_n778), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n775), .A2(G106gat), .A3(new_n534), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n709), .A2(new_n686), .A3(new_n756), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n803), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n806), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n805), .A2(new_n806), .B1(new_n807), .B2(new_n810), .ZN(G1339gat));
  NAND2_X1  g610(.A1(new_n670), .A2(new_n584), .ZN(new_n812));
  INV_X1    g611(.A(new_n704), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n620), .B(new_n615), .C1(new_n619), .C2(KEYINPUT10), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n618), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  OAI221_X1 g615(.A(new_n816), .B1(new_n617), .B2(new_n436), .C1(new_n613), .C2(new_n616), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n627), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n627), .A4(new_n817), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n820), .A2(new_n630), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n562), .B1(new_n561), .B2(new_n564), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n570), .A2(new_n571), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n578), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n828), .A2(new_n582), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n813), .A2(new_n822), .A3(new_n823), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n699), .A2(new_n703), .A3(new_n830), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n820), .A2(new_n630), .A3(new_n821), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT115), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n633), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n830), .B1(new_n835), .B2(new_n631), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n583), .A3(new_n630), .A4(new_n821), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n831), .A2(new_n834), .B1(new_n704), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n812), .B1(new_n839), .B2(new_n649), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n686), .A2(new_n725), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n424), .A2(new_n475), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(KEYINPUT116), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(new_n843), .A3(new_n841), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(new_n236), .A3(new_n584), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n840), .A2(new_n527), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n534), .A2(new_n523), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n424), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n583), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n849), .A2(new_n855), .ZN(G1340gat));
  NAND3_X1  g655(.A1(new_n844), .A2(new_n634), .A3(new_n847), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n711), .A2(G120gat), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n857), .A2(G120gat), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT117), .ZN(G1341gat));
  OAI21_X1  g659(.A(G127gat), .B1(new_n848), .B2(new_n712), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n854), .A2(new_n229), .A3(new_n649), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1342gat));
  NOR3_X1   g662(.A1(new_n853), .A2(G134gat), .A3(new_n668), .ZN(new_n864));
  XNOR2_X1  g663(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n848), .B2(new_n668), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1343gat));
  AND2_X1   g667(.A1(new_n205), .A2(new_n207), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n526), .A2(new_n843), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(new_n840), .B2(new_n686), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n686), .A2(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n831), .A2(new_n834), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n838), .A2(new_n668), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n712), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n878), .B2(new_n812), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n871), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n870), .B1(new_n880), .B2(new_n584), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n683), .A2(new_n534), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n850), .A2(new_n473), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n583), .A2(new_n204), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT121), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g685(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n887));
  NAND3_X1  g686(.A1(new_n881), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT120), .B(new_n871), .C1(new_n873), .C2(new_n879), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n583), .A3(new_n891), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n892), .A2(new_n870), .B1(new_n883), .B2(new_n885), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n888), .B1(new_n893), .B2(new_n894), .ZN(G1344gat));
  NAND3_X1  g694(.A1(new_n890), .A2(new_n634), .A3(new_n891), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n209), .A2(KEYINPUT59), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n833), .B2(new_n668), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n821), .A2(new_n630), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n901), .A2(new_n762), .A3(KEYINPUT124), .A4(new_n820), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n902), .A3(new_n830), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n649), .B1(new_n903), .B2(new_n876), .ZN(new_n904));
  INV_X1    g703(.A(new_n812), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n686), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n840), .A2(new_n686), .A3(new_n872), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n910), .A2(new_n634), .A3(new_n871), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT59), .B1(new_n911), .B2(new_n209), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n898), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n883), .A2(new_n209), .A3(new_n634), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT123), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1345gat));
  NAND2_X1  g715(.A1(new_n890), .A2(new_n891), .ZN(new_n917));
  OAI21_X1  g716(.A(G155gat), .B1(new_n917), .B2(new_n712), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n883), .A2(new_n252), .A3(new_n649), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1346gat));
  NOR3_X1   g719(.A1(new_n917), .A2(new_n253), .A3(new_n704), .ZN(new_n921));
  AOI21_X1  g720(.A(G162gat), .B1(new_n883), .B2(new_n762), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n473), .A2(new_n527), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n842), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n300), .A3(new_n584), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n840), .A2(new_n475), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n473), .A3(new_n851), .ZN(new_n928));
  AOI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n583), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n926), .A2(new_n929), .ZN(G1348gat));
  AOI21_X1  g729(.A(G176gat), .B1(new_n928), .B2(new_n634), .ZN(new_n931));
  INV_X1    g730(.A(new_n925), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n711), .B1(new_n317), .B2(new_n318), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(G1349gat));
  OAI21_X1  g733(.A(new_n349), .B1(new_n925), .B2(new_n712), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n928), .A2(new_n288), .A3(new_n649), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n928), .A2(new_n289), .A3(new_n813), .ZN(new_n939));
  OAI21_X1  g738(.A(G190gat), .B1(new_n925), .B2(new_n668), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n683), .A2(new_n534), .A3(new_n473), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n927), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n583), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n526), .A2(new_n924), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n949), .B1(new_n908), .B2(new_n909), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n583), .A2(G197gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  INV_X1    g751(.A(G204gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n947), .A2(new_n953), .A3(new_n634), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n955));
  INV_X1    g754(.A(new_n950), .ZN(new_n956));
  OAI21_X1  g755(.A(G204gat), .B1(new_n956), .B2(new_n711), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n947), .A2(new_n367), .A3(new_n649), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961));
  INV_X1    g760(.A(new_n949), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n910), .A2(new_n961), .A3(new_n649), .A4(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n950), .B2(new_n649), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n963), .A2(G211gat), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n968), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n960), .B1(new_n967), .B2(new_n970), .ZN(G1354gat));
  AOI21_X1  g770(.A(G218gat), .B1(new_n947), .B2(new_n813), .ZN(new_n972));
  AOI211_X1 g771(.A(new_n376), .B(new_n668), .C1(new_n950), .C2(KEYINPUT127), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G1355gat));
endmodule


