//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  INV_X1    g0005(.A(KEYINPUT64), .ZN(new_n206));
  NAND3_X1  g0006(.A1(new_n201), .A2(new_n206), .A3(new_n202), .ZN(new_n207));
  AND3_X1   g0007(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n210), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n221), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XOR2_X1   g0033(.A(G226), .B(G232), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT67), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n224), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n225), .A2(new_n254), .ZN(new_n255));
  OAI22_X1  g0055(.A1(new_n255), .A2(new_n202), .B1(new_n225), .B2(G68), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n225), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n205), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n253), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT11), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT71), .A2(G1), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT71), .A2(G1), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n253), .B1(new_n263), .B2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G68), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT12), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT71), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT71), .A2(G1), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n269), .A2(G13), .A3(G20), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G68), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n271), .A2(KEYINPUT12), .A3(G68), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n260), .B(new_n265), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT69), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT69), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n268), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT70), .ZN(new_n284));
  AND2_X1   g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n224), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT70), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(new_n289), .A3(new_n268), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n284), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n285), .A2(new_n224), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n281), .A2(new_n277), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT72), .B1(new_n263), .B2(new_n293), .ZN(new_n294));
  AND4_X1   g0094(.A1(KEYINPUT72), .A2(new_n269), .A3(new_n293), .A4(new_n270), .ZN(new_n295));
  OAI211_X1 g0095(.A(G238), .B(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT13), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n213), .A2(G1698), .ZN(new_n298));
  AND2_X1   g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NOR2_X1   g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n298), .B1(G226), .B2(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G97), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n286), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n291), .A2(new_n296), .A3(new_n297), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT75), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n292), .B1(new_n301), .B2(new_n302), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n269), .A2(new_n293), .A3(new_n270), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT72), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n269), .A2(new_n293), .A3(KEYINPUT72), .A4(new_n270), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n286), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n307), .B1(new_n312), .B2(G238), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT75), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n297), .A4(new_n291), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n291), .A2(new_n296), .A3(new_n304), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT13), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n306), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(G179), .A3(new_n305), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n319), .B1(new_n318), .B2(G169), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n276), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n317), .A2(G190), .A3(new_n305), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n317), .A2(KEYINPUT76), .A3(G190), .A4(new_n305), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n276), .B1(new_n318), .B2(G200), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n329), .A2(KEYINPUT77), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT77), .B1(new_n329), .B2(new_n330), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n324), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(G244), .B(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n291), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G1698), .ZN(new_n336));
  OAI211_X1 g0136(.A(G232), .B(new_n336), .C1(new_n299), .C2(new_n300), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT73), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n254), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n343), .A2(KEYINPUT73), .A3(G232), .A4(new_n336), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(G238), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n341), .A2(G107), .A3(new_n342), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n286), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n335), .A2(G190), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n351), .A2(new_n257), .B1(new_n225), .B2(new_n205), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(new_n255), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n253), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n272), .A2(new_n205), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n264), .A2(G77), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n348), .B1(new_n339), .B2(new_n344), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n291), .B(new_n334), .C1(new_n359), .C2(new_n292), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n360), .B2(G200), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT74), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n350), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI211_X1 g0163(.A(KEYINPUT74), .B(new_n358), .C1(new_n360), .C2(G200), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n349), .A2(new_n368), .A3(new_n291), .A4(new_n334), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n369), .A3(new_n358), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(G232), .B(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n373));
  OR2_X1    g0173(.A1(G223), .A2(G1698), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(G226), .B2(new_n336), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n299), .A2(new_n300), .ZN(new_n376));
  INV_X1    g0176(.A(G87), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n375), .A2(new_n376), .B1(new_n254), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n286), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n291), .A2(new_n373), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G200), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n291), .A2(new_n373), .A3(G190), .A4(new_n379), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n384));
  INV_X1    g0184(.A(G159), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n255), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n212), .A2(new_n273), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n201), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT79), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT79), .B(G20), .C1(new_n387), .C2(new_n201), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g0192(.A(KEYINPUT78), .B(KEYINPUT7), .Z(new_n393));
  NAND3_X1  g0193(.A1(new_n341), .A2(new_n225), .A3(new_n342), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n376), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n273), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n384), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n225), .A3(new_n376), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n394), .A2(KEYINPUT7), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(G68), .A3(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n401), .A2(KEYINPUT16), .A3(new_n391), .A4(new_n390), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n402), .A3(new_n253), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n271), .A2(new_n353), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n264), .B2(new_n353), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n383), .A2(KEYINPUT17), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n403), .A2(new_n381), .A3(new_n405), .A4(new_n382), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n343), .A2(G223), .A3(G1698), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n343), .A2(G222), .A3(new_n336), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n412), .C1(new_n205), .C2(new_n343), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n286), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n312), .A2(G226), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(new_n291), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n366), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n225), .B1(new_n204), .B2(new_n207), .ZN(new_n418));
  INV_X1    g0218(.A(G150), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n353), .A2(new_n257), .B1(new_n419), .B2(new_n255), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n253), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n271), .A2(G50), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(G50), .B2(new_n264), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n414), .A2(new_n415), .A3(new_n368), .A4(new_n291), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n417), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n416), .A2(G200), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT9), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n414), .A2(new_n415), .A3(G190), .A4(new_n291), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT9), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT10), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n430), .A2(new_n432), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT10), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n427), .A4(new_n431), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n426), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n380), .A2(G169), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n368), .B2(new_n380), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n403), .A2(new_n405), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n442), .B1(new_n440), .B2(new_n441), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n372), .A2(new_n410), .A3(new_n438), .A4(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n333), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT19), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n225), .B1(new_n302), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(G97), .A2(G107), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n377), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n225), .B(G68), .C1(new_n299), .C2(new_n300), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n448), .B1(new_n257), .B2(new_n214), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT84), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT84), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n452), .A2(new_n453), .A3(new_n457), .A4(new_n454), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n253), .A3(new_n458), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n252), .A2(new_n224), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n269), .A2(G33), .A3(new_n270), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n271), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT82), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n271), .A2(new_n461), .A3(new_n460), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n351), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n272), .A2(new_n351), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n459), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(G238), .B(new_n336), .C1(new_n299), .C2(new_n300), .ZN(new_n470));
  OAI211_X1 g0270(.A(G244), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G116), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n286), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n269), .A2(G45), .A3(new_n270), .ZN(new_n475));
  INV_X1    g0275(.A(G250), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n286), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n263), .A2(G45), .A3(new_n287), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n366), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n286), .A2(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n368), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n469), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT6), .ZN(new_n485));
  AND2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(new_n450), .ZN(new_n487));
  INV_X1    g0287(.A(G107), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(G97), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT81), .ZN(new_n490));
  NAND2_X1  g0290(.A1(KEYINPUT6), .A2(G97), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(G107), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G20), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n225), .A2(new_n254), .A3(G77), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n488), .B1(new_n395), .B2(new_n396), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n253), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n272), .A2(new_n214), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n463), .A2(G97), .A3(new_n465), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g0301(.A1(KEYINPUT4), .A2(G244), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n336), .B(new_n502), .C1(new_n299), .C2(new_n300), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  INV_X1    g0304(.A(G244), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n341), .B2(new_n342), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n503), .B(new_n504), .C1(new_n506), .C2(KEYINPUT4), .ZN(new_n507));
  OAI21_X1  g0307(.A(G250), .B1(new_n299), .B2(new_n300), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n336), .B1(new_n508), .B2(KEYINPUT4), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n286), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(G45), .B1(new_n281), .B2(KEYINPUT5), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n511), .A2(new_n262), .A3(new_n261), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n286), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G257), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n269), .A2(new_n270), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT83), .B1(new_n516), .B2(new_n511), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n513), .B(G274), .C1(new_n285), .C2(new_n224), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT83), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT5), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n277), .B1(new_n521), .B2(G41), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n263), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n517), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n510), .A2(new_n515), .A3(new_n368), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n510), .A2(new_n515), .A3(new_n524), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n366), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n501), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(G200), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n500), .A2(new_n499), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n510), .A2(new_n515), .A3(G190), .A4(new_n524), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n529), .A2(new_n498), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n474), .A2(G190), .A3(new_n479), .ZN(new_n533));
  INV_X1    g0333(.A(G200), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n474), .B2(new_n479), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n463), .A2(G87), .A3(new_n465), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT85), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n463), .A2(KEYINPUT85), .A3(G87), .A4(new_n465), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n459), .A2(new_n468), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n536), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND4_X1   g0343(.A1(new_n484), .A2(new_n528), .A3(new_n532), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n476), .A2(new_n336), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n215), .A2(G1698), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(new_n546), .C1(new_n299), .C2(new_n300), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G294), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n286), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n522), .A2(new_n269), .A3(new_n270), .ZN(new_n551));
  INV_X1    g0351(.A(new_n513), .ZN(new_n552));
  OAI211_X1 g0352(.A(G264), .B(new_n292), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n524), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n534), .ZN(new_n555));
  INV_X1    g0355(.A(G190), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n524), .A2(new_n550), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(KEYINPUT86), .A2(G87), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n225), .B(new_n559), .C1(new_n299), .C2(new_n300), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT22), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT22), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n343), .A2(new_n562), .A3(new_n225), .A4(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT24), .ZN(new_n565));
  INV_X1    g0365(.A(new_n257), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n225), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n488), .A2(KEYINPUT23), .A3(G20), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n566), .A2(G116), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n564), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n565), .B1(new_n564), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n253), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n463), .A2(G107), .A3(new_n465), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n272), .A2(KEYINPUT25), .A3(new_n488), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT25), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n271), .B2(G107), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n558), .A2(new_n573), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n564), .A2(new_n570), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT24), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n564), .A2(new_n565), .A3(new_n570), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n579), .B1(new_n585), .B2(new_n253), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n554), .A2(new_n366), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G179), .B2(new_n554), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n581), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G270), .B(new_n292), .C1(new_n551), .C2(new_n552), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G257), .A2(G1698), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n336), .A2(G264), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n343), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n376), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n286), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n524), .A2(new_n590), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(G116), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n272), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n271), .A2(new_n461), .A3(new_n460), .A4(G116), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n252), .A2(new_n224), .B1(G20), .B2(new_n598), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n504), .B(new_n225), .C1(G33), .C2(new_n214), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n601), .A2(KEYINPUT20), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT20), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n599), .B(new_n600), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n597), .A2(new_n605), .A3(G169), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(G179), .A2(new_n524), .A3(new_n590), .A4(new_n596), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n606), .A2(new_n607), .B1(new_n609), .B2(new_n605), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n605), .B1(new_n597), .B2(G200), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n556), .B2(new_n597), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n589), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n447), .A2(new_n544), .A3(new_n614), .ZN(G372));
  NAND2_X1  g0415(.A1(new_n434), .A2(new_n437), .ZN(new_n616));
  INV_X1    g0416(.A(new_n410), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n371), .B1(new_n331), .B2(new_n332), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n324), .ZN(new_n619));
  INV_X1    g0419(.A(new_n445), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n426), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n528), .A2(new_n532), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n543), .A2(new_n484), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n608), .B(new_n610), .C1(new_n586), .C2(new_n588), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .A4(new_n581), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n501), .A2(new_n525), .A3(new_n527), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n484), .A4(new_n543), .ZN(new_n630));
  INV_X1    g0430(.A(new_n484), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n530), .A2(new_n498), .B1(new_n526), .B2(new_n366), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n543), .A2(new_n632), .A3(new_n484), .A4(new_n525), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n633), .B2(KEYINPUT26), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n627), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n447), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n623), .A2(new_n636), .ZN(G369));
  INV_X1    g0437(.A(new_n589), .ZN(new_n638));
  INV_X1    g0438(.A(G13), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n263), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n638), .B1(new_n586), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n586), .A2(new_n588), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n650), .B2(new_n647), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n608), .A2(new_n610), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(new_n605), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n613), .B2(new_n654), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n646), .B1(new_n608), .B2(new_n610), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n638), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n649), .A2(new_n647), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n658), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n229), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n451), .A2(G116), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n222), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT28), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n614), .A2(new_n544), .A3(new_n647), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n524), .A2(new_n590), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n292), .B1(new_n547), .B2(new_n548), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n514), .B2(G264), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n292), .B1(new_n376), .B2(new_n594), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n368), .B1(new_n676), .B2(new_n593), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n673), .A2(new_n482), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n672), .B1(new_n678), .B2(new_n526), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n524), .A2(new_n590), .A3(new_n596), .A4(G179), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n550), .A2(new_n553), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n680), .A2(new_n480), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n510), .A2(new_n515), .A3(KEYINPUT30), .A4(new_n524), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(new_n684), .A3(KEYINPUT87), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT87), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n678), .B2(new_n683), .ZN(new_n687));
  AOI21_X1  g0487(.A(G179), .B1(new_n675), .B2(new_n524), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(new_n480), .A3(new_n526), .A4(new_n597), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n679), .A2(new_n685), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n646), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n671), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n635), .A2(new_n697), .A3(new_n647), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n635), .B2(new_n647), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n670), .B1(new_n700), .B2(G1), .ZN(G364));
  AOI21_X1  g0501(.A(new_n268), .B1(new_n640), .B2(G45), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n665), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n657), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(G330), .B2(new_n656), .ZN(new_n706));
  INV_X1    g0506(.A(new_n704), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n224), .B1(G20), .B2(new_n366), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n225), .A2(G179), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(G190), .A3(G200), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G87), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n343), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n225), .A2(new_n368), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G200), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n556), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G190), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n710), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G159), .ZN(new_n723));
  XOR2_X1   g0523(.A(KEYINPUT89), .B(KEYINPUT32), .Z(new_n724));
  OAI22_X1  g0524(.A1(new_n719), .A2(new_n202), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n556), .A2(G179), .A3(G200), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n225), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n725), .B1(G97), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n716), .A2(G190), .A3(new_n534), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n716), .A2(new_n720), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n212), .B1(new_n731), .B2(new_n205), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n723), .B2(new_n724), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n710), .A2(new_n556), .A3(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n488), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n717), .A2(G190), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(G68), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n715), .A2(new_n729), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G322), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G311), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n376), .B1(new_n731), .B2(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n740), .B(new_n742), .C1(G329), .C2(new_n722), .ZN(new_n743));
  INV_X1    g0543(.A(new_n734), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G283), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT33), .B(G317), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G294), .A2(new_n728), .B1(new_n736), .B2(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n718), .A2(G326), .B1(new_n712), .B2(G303), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n743), .A2(new_n745), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n709), .B1(new_n738), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n708), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n343), .A2(G355), .A3(new_n229), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G116), .B2(new_n229), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT88), .Z(new_n757));
  NOR2_X1   g0557(.A1(new_n250), .A2(new_n277), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n664), .A2(new_n343), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n278), .A2(new_n280), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n223), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n757), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n707), .B(new_n750), .C1(new_n754), .C2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n753), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n656), .B2(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n706), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(G396));
  NAND2_X1  g0567(.A1(new_n646), .A2(new_n358), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n363), .B2(new_n364), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT93), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n370), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n358), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n360), .B2(new_n366), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(KEYINPUT93), .A3(new_n369), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(KEYINPUT94), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  AND4_X1   g0576(.A1(KEYINPUT93), .A2(new_n367), .A3(new_n369), .A4(new_n358), .ZN(new_n777));
  AOI21_X1  g0577(.A(KEYINPUT93), .B1(new_n773), .B2(new_n369), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT94), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n534), .B1(new_n335), .B2(new_n349), .ZN(new_n781));
  OAI21_X1  g0581(.A(KEYINPUT74), .B1(new_n781), .B2(new_n358), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n361), .A2(new_n362), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n782), .A2(new_n783), .A3(new_n350), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n779), .A2(new_n780), .A3(new_n784), .A4(new_n768), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n776), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(new_n635), .A3(new_n647), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n633), .A2(KEYINPUT26), .ZN(new_n788));
  AND3_X1   g0588(.A1(new_n788), .A2(new_n484), .A3(new_n630), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n646), .B1(new_n789), .B2(new_n627), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n776), .B(new_n785), .C1(new_n370), .C2(new_n647), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n696), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n704), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n793), .B2(new_n792), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n709), .A2(new_n752), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n704), .B1(G77), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  INV_X1    g0598(.A(new_n736), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n798), .A2(new_n799), .B1(new_n719), .B2(new_n594), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G87), .B2(new_n744), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n343), .B1(new_n722), .B2(G311), .ZN(new_n802));
  INV_X1    g0602(.A(new_n730), .ZN(new_n803));
  INV_X1    g0603(.A(new_n731), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n803), .A2(G294), .B1(new_n804), .B2(G116), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n728), .A2(G97), .B1(new_n712), .B2(G107), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n801), .A2(new_n802), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G137), .A2(new_n718), .B1(new_n736), .B2(G150), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT91), .Z(new_n809));
  INV_X1    g0609(.A(G143), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n810), .B2(new_n730), .C1(new_n385), .C2(new_n731), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT92), .B(KEYINPUT34), .Z(new_n812));
  XOR2_X1   g0612(.A(new_n811), .B(new_n812), .Z(new_n813));
  AOI22_X1  g0613(.A1(new_n728), .A2(G58), .B1(new_n712), .B2(G50), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n744), .A2(G68), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n376), .B1(new_n722), .B2(G132), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n807), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n797), .B1(new_n818), .B2(new_n708), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n752), .B2(new_n791), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n795), .A2(KEYINPUT95), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(KEYINPUT95), .B1(new_n795), .B2(new_n820), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G384));
  NOR2_X1   g0624(.A1(new_n263), .A2(new_n640), .ZN(new_n825));
  INV_X1    g0625(.A(G330), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n276), .A2(new_n646), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n329), .A2(new_n330), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT77), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n329), .A2(KEYINPUT77), .A3(new_n330), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n827), .B1(new_n832), .B2(new_n324), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n324), .B(new_n827), .C1(new_n331), .C2(new_n332), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT97), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n695), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n671), .A2(new_n693), .A3(KEYINPUT97), .A4(new_n694), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(new_n791), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n440), .A2(new_n441), .ZN(new_n843));
  INV_X1    g0643(.A(new_n644), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n441), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n845), .A3(new_n407), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(KEYINPUT37), .ZN(new_n847));
  INV_X1    g0647(.A(new_n384), .ZN(new_n848));
  INV_X1    g0648(.A(new_n392), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n401), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n402), .A2(new_n253), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n405), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT96), .B1(new_n852), .B2(new_n844), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(KEYINPUT96), .A3(new_n844), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n852), .A2(new_n440), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n854), .A2(new_n407), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n847), .B1(new_n857), .B2(KEYINPUT37), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n852), .A2(KEYINPUT96), .A3(new_n844), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n853), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n410), .B2(new_n445), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n842), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n843), .A2(KEYINPUT18), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n863), .A2(new_n406), .A3(new_n864), .A4(new_n409), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n854), .A2(new_n855), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n856), .A2(new_n407), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n860), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n867), .B(KEYINPUT38), .C1(new_n870), .C2(new_n847), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n862), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT40), .B1(new_n841), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT40), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n846), .B(new_n868), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n845), .B1(new_n410), .B2(new_n445), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n842), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n877), .B2(new_n871), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n873), .B1(new_n841), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n447), .A2(new_n838), .A3(new_n839), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n826), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n862), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT39), .B1(new_n877), .B2(new_n871), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n324), .A2(new_n646), .ZN(new_n885));
  OR3_X1    g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n620), .A2(new_n644), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n779), .A2(new_n646), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n827), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n333), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n787), .A2(new_n889), .B1(new_n891), .B2(new_n834), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n872), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n886), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n447), .B1(new_n698), .B2(new_n699), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n623), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n894), .B(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n825), .B1(new_n882), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n897), .B2(new_n882), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n598), .B(new_n227), .C1(new_n493), .C2(KEYINPUT35), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(KEYINPUT35), .B2(new_n493), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT36), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n387), .A2(new_n222), .A3(new_n205), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n273), .A2(G50), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n639), .B(new_n516), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n899), .A2(new_n902), .A3(new_n905), .ZN(G367));
  NAND2_X1  g0706(.A1(new_n242), .A2(new_n759), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n907), .B(new_n754), .C1(new_n229), .C2(new_n351), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT103), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n707), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n909), .B2(new_n908), .ZN(new_n911));
  INV_X1    g0711(.A(G317), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n730), .A2(new_n594), .B1(new_n721), .B2(new_n912), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n343), .B(new_n913), .C1(G283), .C2(new_n804), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n712), .A2(G116), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT46), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n734), .A2(new_n214), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(G107), .B2(new_n728), .ZN(new_n918));
  AOI22_X1  g0718(.A1(G294), .A2(new_n736), .B1(new_n718), .B2(G311), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n914), .A2(new_n916), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT104), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n727), .A2(new_n273), .B1(new_n730), .B2(new_n419), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT105), .ZN(new_n923));
  INV_X1    g0723(.A(G137), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n343), .B1(new_n721), .B2(new_n924), .C1(new_n202), .C2(new_n731), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n810), .A2(new_n719), .B1(new_n799), .B2(new_n385), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n212), .A2(new_n711), .B1(new_n734), .B2(new_n205), .ZN(new_n927));
  OR4_X1    g0727(.A1(new_n923), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n920), .A2(KEYINPUT104), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT47), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n911), .B1(new_n931), .B2(new_n708), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n541), .A2(new_n542), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n646), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n625), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n484), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n932), .B1(new_n764), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n660), .B1(new_n651), .B2(new_n659), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(new_n657), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n700), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT102), .Z(new_n941));
  NOR2_X1   g0741(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n501), .A2(new_n646), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n624), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n628), .A2(new_n646), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n942), .B1(new_n662), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n944), .A2(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n660), .A2(new_n661), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(KEYINPUT100), .C2(KEYINPUT44), .ZN(new_n950));
  NAND2_X1  g0750(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT99), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n662), .A2(new_n953), .A3(new_n946), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT99), .B1(new_n948), .B2(new_n949), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT45), .B1(new_n954), .B2(new_n955), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n658), .A2(KEYINPUT101), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n941), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n700), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n665), .B(KEYINPUT41), .Z(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n703), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n658), .A2(new_n948), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT98), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n948), .A2(new_n660), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(KEYINPUT42), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n528), .B1(new_n944), .B2(new_n650), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n973), .A2(KEYINPUT42), .B1(new_n647), .B2(new_n976), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n975), .A2(new_n977), .B1(KEYINPUT43), .B2(new_n936), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n970), .A2(new_n971), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n970), .B2(new_n971), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n937), .B1(new_n966), .B2(new_n982), .ZN(G387));
  NOR2_X1   g0783(.A1(new_n651), .A2(new_n764), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n667), .A2(new_n664), .A3(new_n376), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n488), .B2(new_n664), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT106), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n239), .B1(new_n278), .B2(new_n280), .ZN(new_n988));
  INV_X1    g0788(.A(new_n353), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n202), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT50), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n667), .B(new_n277), .C1(new_n273), .C2(new_n205), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n759), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n987), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n754), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n704), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n730), .A2(new_n202), .B1(new_n731), .B2(new_n273), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n376), .B(new_n997), .C1(G150), .C2(new_n722), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n736), .A2(new_n989), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n466), .A2(new_n728), .B1(new_n718), .B2(G159), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n917), .B1(G77), .B2(new_n712), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n803), .A2(G317), .B1(new_n804), .B2(G303), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n719), .B2(new_n739), .C1(new_n741), .C2(new_n799), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT48), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n728), .A2(G283), .B1(new_n712), .B2(G294), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n343), .B1(new_n722), .B2(G326), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(new_n598), .C2(new_n734), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1002), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n984), .B(new_n996), .C1(new_n1015), .C2(new_n708), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n703), .B2(new_n939), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n939), .A2(new_n700), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n940), .A2(new_n665), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(G393));
  INV_X1    g0820(.A(new_n958), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1021), .A2(new_n952), .A3(new_n658), .A4(new_n956), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT108), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT108), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(new_n658), .C2(new_n959), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(new_n702), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n948), .A2(new_n753), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n247), .A2(new_n664), .A3(new_n343), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n754), .B1(new_n214), .B2(new_n229), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n704), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n719), .A2(new_n912), .B1(new_n741), .B2(new_n730), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT52), .ZN(new_n1032));
  INV_X1    g0832(.A(G294), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n376), .B1(new_n731), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G322), .B2(new_n722), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n735), .B1(G116), .B2(new_n728), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n736), .A2(G303), .B1(new_n712), .B2(G283), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(KEYINPUT110), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n719), .A2(new_n419), .B1(new_n385), .B2(new_n730), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n711), .A2(new_n273), .B1(new_n721), .B2(new_n810), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT109), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT109), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n727), .A2(new_n205), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n343), .B1(new_n731), .B2(new_n353), .C1(new_n377), .C2(new_n734), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(G50), .C2(new_n736), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1038), .A2(KEYINPUT110), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1039), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1030), .B1(new_n1050), .B2(new_n708), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1026), .B1(new_n1027), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n666), .B1(new_n941), .B2(new_n961), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1025), .A2(new_n940), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(KEYINPUT111), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT111), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1052), .B1(new_n1056), .B2(new_n1057), .ZN(G390));
  INV_X1    g0858(.A(KEYINPUT113), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n447), .A2(new_n838), .A3(G330), .A4(new_n839), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n621), .A2(new_n895), .A3(new_n1060), .A4(new_n622), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n787), .A2(new_n889), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n891), .A2(new_n834), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n696), .A2(new_n791), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n787), .A2(new_n891), .A3(new_n834), .A4(new_n889), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AND4_X1   g0867(.A1(G330), .A2(new_n838), .A3(new_n791), .A4(new_n839), .ZN(new_n1068));
  AND4_X1   g0868(.A1(new_n787), .A2(new_n891), .A3(new_n834), .A4(new_n889), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n892), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1059), .B(new_n1061), .C1(new_n1067), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1067), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1061), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT113), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n877), .A2(new_n871), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n888), .B1(new_n790), .B2(new_n786), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n885), .B(new_n1076), .C1(new_n836), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT112), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT112), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1064), .A2(new_n1080), .A3(new_n885), .A4(new_n1076), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n885), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n883), .A2(new_n884), .B1(new_n892), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n836), .A2(new_n840), .A3(new_n826), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1063), .A2(new_n696), .A3(new_n791), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1079), .A2(new_n1087), .A3(new_n1083), .A4(new_n1081), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n666), .B1(new_n1075), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1088), .B(new_n1086), .C1(new_n1071), .C2(new_n1074), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n751), .B1(new_n883), .B2(new_n884), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n704), .B1(new_n989), .B2(new_n796), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n730), .A2(new_n598), .B1(new_n721), .B2(new_n1033), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n343), .B(new_n1095), .C1(G97), .C2(new_n804), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n713), .A3(new_n815), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1045), .B1(G283), .B2(new_n718), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n488), .B2(new_n799), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G159), .A2(new_n728), .B1(new_n718), .B2(G128), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n202), .B2(new_n734), .C1(new_n924), .C2(new_n799), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1102));
  OR3_X1    g0902(.A1(new_n1102), .A2(new_n711), .A3(new_n419), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT54), .B(G143), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n804), .A2(new_n1105), .B1(new_n722), .B2(G125), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n376), .B1(new_n803), .B2(G132), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1102), .B1(new_n711), .B2(new_n419), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1097), .A2(new_n1099), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1110), .A2(KEYINPUT115), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n709), .B1(new_n1110), .B2(KEYINPUT115), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1094), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1093), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1089), .B2(new_n702), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1092), .A2(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(KEYINPUT118), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1063), .A2(new_n791), .A3(new_n838), .A4(new_n839), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1076), .A2(KEYINPUT40), .ZN(new_n1120));
  OAI21_X1  g0920(.A(G330), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1118), .B1(new_n873), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n826), .B1(new_n841), .B2(new_n878), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n872), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n874), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(KEYINPUT118), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n844), .A2(new_n424), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n438), .B(new_n1127), .Z(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1128), .B(new_n1129), .Z(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1122), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1123), .A2(new_n1125), .A3(KEYINPUT118), .A4(new_n1130), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n894), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n894), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1136), .A3(new_n1133), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n703), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1130), .A2(new_n751), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n704), .B1(G50), .B2(new_n796), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT116), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n799), .A2(new_n214), .B1(new_n734), .B2(new_n212), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G116), .B2(new_n718), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n376), .A2(new_n281), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G283), .B2(new_n722), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n803), .A2(G107), .B1(new_n804), .B2(new_n466), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n728), .A2(G68), .B1(new_n712), .B2(G77), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT58), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1144), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n718), .A2(G125), .ZN(new_n1153));
  INV_X1    g0953(.A(G132), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n799), .B2(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n803), .A2(G128), .B1(new_n804), .B2(G137), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n711), .B2(new_n1104), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G150), .C2(new_n728), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n744), .A2(G159), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G33), .B(G41), .C1(new_n722), .C2(G124), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1152), .B1(new_n1149), .B2(new_n1148), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1141), .B1(new_n1165), .B2(new_n708), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1139), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT117), .Z(new_n1168));
  NAND2_X1  g0968(.A1(new_n1138), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1091), .A2(new_n1073), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n1137), .A3(new_n1135), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n666), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1132), .A2(new_n1136), .A3(new_n1133), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1136), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(KEYINPUT57), .A3(new_n1170), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1169), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(G375));
  NAND3_X1  g0979(.A1(new_n1070), .A2(new_n1061), .A3(new_n1067), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1075), .A2(new_n965), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1072), .A2(new_n703), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n704), .B1(G68), .B2(new_n796), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n730), .A2(new_n924), .B1(new_n731), .B2(new_n419), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n376), .B(new_n1184), .C1(G128), .C2(new_n722), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n712), .A2(G159), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G132), .A2(new_n718), .B1(new_n736), .B2(new_n1105), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n728), .A2(G50), .B1(new_n744), .B2(G58), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n719), .A2(new_n1033), .B1(new_n734), .B2(new_n205), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n799), .A2(new_n598), .B1(new_n711), .B2(new_n214), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n376), .B1(new_n721), .B2(new_n594), .C1(new_n488), .C2(new_n731), .ZN(new_n1192));
  OR3_X1    g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n727), .A2(new_n351), .B1(new_n730), .B2(new_n798), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT119), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1189), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1183), .B1(new_n1196), .B2(new_n708), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n1063), .B2(new_n752), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1182), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1181), .A2(new_n1200), .ZN(G381));
  INV_X1    g1001(.A(new_n1057), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1055), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n964), .B1(new_n962), .B2(new_n700), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n980), .B(new_n981), .C1(new_n1204), .C2(new_n703), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1203), .A2(new_n1205), .A3(new_n937), .A4(new_n1052), .ZN(new_n1206));
  OR3_X1    g1006(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1206), .A2(G381), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT120), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(G375), .A2(G378), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(G407));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n645), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(G407), .A2(G213), .A3(new_n1212), .ZN(G409));
  NAND2_X1  g1013(.A1(new_n645), .A2(G213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1176), .A2(new_n703), .B1(new_n1139), .B2(new_n1166), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1176), .A2(new_n965), .A3(new_n1170), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G378), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1178), .B2(G378), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1214), .B1(new_n1218), .B2(KEYINPUT121), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1115), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1169), .B(new_n1220), .C1(new_n1173), .C2(new_n1177), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT121), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n1217), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT125), .B1(new_n1219), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1075), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1225), .A2(new_n1180), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT122), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1180), .A2(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n665), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT123), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1225), .A2(new_n1180), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1229), .A2(new_n665), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT123), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1230), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1199), .B1(new_n1232), .B2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(G384), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1199), .B(new_n823), .C1(new_n1232), .C2(new_n1236), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G2897), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1214), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1238), .A2(new_n1239), .B1(new_n1241), .B2(new_n1214), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1218), .A2(KEYINPUT121), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1222), .B1(new_n1221), .B2(new_n1217), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT125), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1214), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1224), .A2(new_n1245), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT126), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1224), .A2(new_n1252), .A3(new_n1245), .A4(new_n1249), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(new_n766), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT127), .B1(G390), .B2(G387), .ZN(new_n1255));
  AND2_X1   g1055(.A1(G390), .A2(G387), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G390), .A2(G387), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1254), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1206), .A2(new_n1259), .A3(KEYINPUT127), .A4(new_n1260), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1257), .A2(new_n1258), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1169), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(G378), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1217), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1240), .A2(new_n1267), .A3(KEYINPUT63), .A4(new_n1214), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1262), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1246), .A2(new_n1247), .A3(new_n1240), .A4(new_n1214), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1251), .A2(new_n1253), .A3(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1267), .A2(new_n1214), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1245), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1240), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT62), .B1(new_n1278), .B2(new_n1276), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1279), .A3(new_n1258), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1270), .A2(KEYINPUT62), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1275), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1273), .A2(new_n1282), .ZN(G405));
  XNOR2_X1  g1083(.A(new_n1178), .B(G378), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1240), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1275), .ZN(G402));
endmodule


