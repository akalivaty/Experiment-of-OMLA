//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(G224), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT89), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  OR2_X1    g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT0), .A3(G128), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n205), .B1(G143), .B2(new_n190), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n194), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n198), .A2(new_n205), .A3(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n201), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n204), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  OAI211_X1 g028(.A(KEYINPUT7), .B(new_n189), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n214), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n189), .A2(KEYINPUT7), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n216), .A2(new_n212), .A3(new_n204), .A4(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT2), .B(G113), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT69), .A2(G116), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT69), .A2(G116), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n221), .A2(KEYINPUT70), .A3(G119), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G116), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n224), .B2(G119), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(G116), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT69), .A2(G116), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT69), .A2(G116), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT70), .B1(new_n233), .B2(G119), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n221), .A2(G119), .A3(new_n222), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n238), .A2(KEYINPUT5), .A3(new_n229), .A4(new_n223), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n224), .A2(KEYINPUT5), .A3(G119), .ZN(new_n240));
  INV_X1    g054(.A(G113), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n220), .A2(new_n235), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G104), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT3), .B1(new_n244), .B2(G107), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT79), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(KEYINPUT79), .B(KEYINPUT3), .C1(new_n244), .C2(G107), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT80), .A2(G107), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT80), .A2(G107), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n247), .A2(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G107), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT81), .B1(new_n254), .B2(G104), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n244), .A3(G107), .ZN(new_n257));
  AOI21_X1  g071(.A(G101), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(G104), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n251), .B2(G104), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n253), .A2(new_n258), .B1(new_n260), .B2(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n243), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G110), .B(G122), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT8), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n215), .A2(new_n218), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT91), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n250), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT80), .A2(G107), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n252), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n255), .A2(new_n257), .ZN(new_n271));
  INV_X1    g085(.A(new_n248), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT79), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n270), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G101), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT82), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n279), .A3(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n275), .B1(new_n253), .B2(new_n258), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(G101), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n219), .B1(new_n230), .B2(new_n234), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n238), .A2(new_n220), .A3(new_n229), .A4(new_n223), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n282), .A2(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n243), .A2(new_n261), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n263), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n291), .B1(new_n265), .B2(new_n266), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n267), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT87), .A2(KEYINPUT6), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n281), .A2(new_n286), .B1(new_n261), .B2(new_n243), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n290), .B1(new_n295), .B2(KEYINPUT86), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n287), .A2(KEYINPUT86), .A3(new_n288), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT86), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n294), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n295), .A2(KEYINPUT86), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .A4(new_n290), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n291), .A2(KEYINPUT6), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n298), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n213), .A2(new_n214), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(new_n189), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n305), .A2(KEYINPUT90), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT90), .B1(new_n305), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n293), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n311), .B(new_n293), .C1(new_n308), .C2(new_n309), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n201), .A2(G140), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT75), .ZN(new_n319));
  OR3_X1    g133(.A1(new_n316), .A2(KEYINPUT75), .A3(G125), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT16), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G146), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n317), .A2(new_n318), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n190), .ZN(new_n327));
  XOR2_X1   g141(.A(KEYINPUT24), .B(G110), .Z(new_n328));
  NAND2_X1  g142(.A1(new_n227), .A2(G128), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n207), .A2(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n328), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n227), .A2(G128), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n329), .B(new_n336), .C1(new_n337), .C2(KEYINPUT23), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G110), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n325), .B(new_n327), .C1(new_n335), .C2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n332), .A2(new_n334), .A3(new_n328), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(G110), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n321), .A2(new_n190), .A3(new_n323), .ZN(new_n344));
  AOI211_X1 g158(.A(KEYINPUT76), .B(new_n343), .C1(new_n344), .C2(new_n325), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n325), .A2(new_n344), .ZN(new_n347));
  INV_X1    g161(.A(new_n343), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n340), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G137), .ZN(new_n351));
  INV_X1    g165(.A(G221), .ZN(new_n352));
  INV_X1    g166(.A(G234), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n352), .A2(new_n353), .A3(G953), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n351), .B(new_n354), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n340), .B(new_n355), .C1(new_n345), .C2(new_n349), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G217), .B1(new_n353), .B2(G902), .ZN(new_n360));
  INV_X1    g174(.A(G902), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n357), .A2(new_n364), .A3(new_n361), .A4(new_n358), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n357), .A2(new_n361), .A3(new_n358), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT77), .B1(new_n366), .B2(KEYINPUT25), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n360), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n363), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n284), .A2(new_n285), .ZN(new_n376));
  INV_X1    g190(.A(G137), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT66), .B1(new_n377), .B2(G134), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT66), .ZN(new_n379));
  INV_X1    g193(.A(G134), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G137), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT65), .B(G131), .Z(new_n383));
  OAI21_X1  g197(.A(KEYINPUT11), .B1(new_n380), .B2(G137), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT11), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n377), .A3(G134), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n382), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G131), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n382), .B2(new_n387), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n200), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n382), .A2(new_n383), .A3(new_n387), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n380), .A2(G137), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n377), .A2(G134), .ZN(new_n394));
  OAI21_X1  g208(.A(G131), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n210), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(KEYINPUT30), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n396), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n391), .A2(KEYINPUT67), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n197), .A2(new_n199), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n387), .A2(new_n378), .A3(new_n381), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G131), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n402), .B2(new_n392), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT67), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n398), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n407));
  OAI211_X1 g221(.A(new_n376), .B(new_n397), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n409));
  INV_X1    g223(.A(G237), .ZN(new_n410));
  INV_X1    g224(.A(G953), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(G210), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n409), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT26), .B(G101), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n413), .B(new_n414), .Z(new_n415));
  NAND4_X1  g229(.A1(new_n391), .A2(new_n284), .A3(new_n285), .A4(new_n396), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n408), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT31), .ZN(new_n418));
  INV_X1    g232(.A(new_n415), .ZN(new_n419));
  INV_X1    g233(.A(new_n376), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n406), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT28), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n420), .A2(KEYINPUT28), .A3(new_n396), .A4(new_n391), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n419), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT31), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n408), .A2(new_n427), .A3(new_n415), .A4(new_n416), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n418), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(G472), .A2(G902), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT32), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT32), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n408), .A2(new_n416), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT72), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(KEYINPUT29), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n419), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT72), .B1(new_n421), .B2(new_n425), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n391), .A2(KEYINPUT67), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n402), .A2(new_n392), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n404), .B1(new_n442), .B2(new_n200), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n396), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n376), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n445), .A2(new_n437), .A3(new_n424), .A4(new_n423), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n440), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n423), .A2(KEYINPUT73), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n376), .B1(new_n398), .B2(new_n403), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n422), .B1(new_n450), .B2(new_n416), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n423), .A2(KEYINPUT73), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n449), .B(KEYINPUT29), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n415), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n361), .B(new_n439), .C1(new_n448), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G472), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n375), .B1(new_n435), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT9), .B(G234), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n352), .B1(new_n459), .B2(new_n361), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n282), .A2(new_n283), .ZN(new_n462));
  INV_X1    g276(.A(new_n280), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n279), .B1(new_n274), .B2(new_n276), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n462), .B(new_n200), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n258), .B(new_n270), .C1(new_n273), .C2(new_n272), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n260), .A2(G101), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT83), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n207), .B1(new_n206), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT83), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n198), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n209), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n466), .B(new_n467), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT10), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n208), .B2(new_n209), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n474), .A2(new_n475), .B1(new_n261), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n388), .A2(new_n390), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n465), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G110), .B(G140), .ZN(new_n480));
  INV_X1    g294(.A(G227), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(G953), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n480), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n466), .A2(new_n467), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n211), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n474), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT12), .B1(new_n487), .B2(new_n442), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n489), .B(new_n478), .C1(new_n486), .C2(new_n474), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n479), .B(new_n484), .C1(new_n488), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n465), .A2(new_n477), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n442), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n484), .B1(new_n493), .B2(new_n479), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n491), .B1(new_n494), .B2(KEYINPUT84), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n491), .A2(KEYINPUT84), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AOI211_X1 g311(.A(G469), .B(G902), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n479), .B1(new_n488), .B2(new_n490), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n483), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n493), .A2(new_n484), .A3(new_n479), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(G469), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G469), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(new_n361), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n461), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n459), .A2(G217), .A3(new_n411), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n207), .B2(G143), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n192), .A2(KEYINPUT96), .A3(G128), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT13), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n512), .A2(new_n513), .B1(new_n207), .B2(G143), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n514), .A2(KEYINPUT97), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n512), .A2(new_n513), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n514), .B2(KEYINPUT97), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n380), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n207), .A2(G143), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n512), .A2(new_n380), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G122), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G116), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT95), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n231), .A2(new_n232), .A3(new_n521), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n525), .A3(new_n251), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n251), .B1(new_n523), .B2(new_n525), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n518), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n512), .A2(new_n519), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G134), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n520), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n526), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n525), .A2(new_n535), .A3(KEYINPUT14), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT98), .B1(new_n524), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n524), .A2(new_n537), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n523), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n534), .B1(new_n541), .B2(G107), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n508), .B1(new_n530), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n523), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n538), .B2(new_n536), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n526), .B(new_n533), .C1(new_n545), .C2(new_n254), .ZN(new_n546));
  INV_X1    g360(.A(new_n508), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n546), .B(new_n547), .C1(new_n518), .C2(new_n529), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n361), .ZN(new_n550));
  INV_X1    g364(.A(G478), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(KEYINPUT15), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n550), .A2(new_n552), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n410), .A2(new_n411), .A3(G214), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(G143), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n383), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n383), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n326), .A2(KEYINPUT19), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n319), .A2(new_n320), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(KEYINPUT19), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n562), .B(new_n325), .C1(G146), .C2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(G113), .B(G122), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G104), .ZN(new_n568));
  OR3_X1    g382(.A1(new_n564), .A2(KEYINPUT92), .A3(new_n190), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n327), .B(KEYINPUT92), .C1(new_n564), .C2(new_n190), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n557), .A2(KEYINPUT18), .A3(G131), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n557), .B1(KEYINPUT18), .B2(G131), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n560), .A2(new_n561), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n558), .A2(KEYINPUT17), .A3(new_n559), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n344), .A4(new_n325), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n568), .B1(new_n579), .B2(new_n573), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n573), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n574), .B1(new_n584), .B2(new_n568), .ZN(new_n585));
  NOR2_X1   g399(.A1(G475), .A2(G902), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI22_X1  g401(.A1(new_n582), .A2(KEYINPUT20), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n575), .A2(new_n580), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT20), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n589), .A2(new_n581), .A3(new_n590), .A4(new_n586), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n568), .ZN(new_n593));
  OR3_X1    g407(.A1(new_n583), .A2(KEYINPUT94), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n583), .B1(KEYINPUT94), .B2(new_n593), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n361), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G475), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n411), .A2(G952), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(G234), .B2(G237), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n361), .B(new_n411), .C1(G234), .C2(G237), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT21), .B(G898), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n555), .A2(new_n592), .A3(new_n597), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n507), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G214), .B1(G237), .B2(G902), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n606), .B(KEYINPUT85), .Z(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n315), .A2(new_n457), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n374), .B(new_n461), .C1(new_n498), .C2(new_n506), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n429), .A2(new_n361), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G472), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n431), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n611), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n495), .B2(new_n497), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n503), .ZN(new_n618));
  INV_X1    g432(.A(new_n506), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n460), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n613), .A2(G472), .B1(new_n429), .B2(new_n430), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(KEYINPUT99), .A3(new_n374), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n550), .A2(new_n551), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n550), .A2(KEYINPUT101), .A3(new_n551), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n548), .B2(KEYINPUT100), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n549), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n551), .A2(G902), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n592), .A2(new_n597), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n634), .A2(new_n635), .A3(new_n602), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n315), .A2(new_n606), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n623), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  INV_X1    g454(.A(new_n606), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n313), .B2(new_n314), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n585), .A2(new_n587), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n590), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n553), .A2(new_n554), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n597), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n623), .A2(new_n643), .A3(new_n602), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT102), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT103), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  AOI21_X1  g466(.A(new_n607), .B1(new_n313), .B2(new_n314), .ZN(new_n653));
  INV_X1    g467(.A(new_n362), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n356), .A2(KEYINPUT36), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n350), .B(new_n655), .Z(new_n656));
  AOI22_X1  g470(.A1(new_n369), .A2(new_n373), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n615), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n653), .A2(new_n605), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT37), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n600), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n599), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n647), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n642), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT106), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n429), .A2(new_n433), .A3(new_n430), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n433), .B1(new_n429), .B2(new_n430), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n456), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n657), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n674), .A2(new_n620), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n315), .A2(new_n677), .A3(new_n606), .A4(new_n669), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n671), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XNOR2_X1  g494(.A(new_n667), .B(KEYINPUT39), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n620), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n682), .B(KEYINPUT40), .Z(new_n683));
  NOR2_X1   g497(.A1(new_n436), .A2(new_n419), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n450), .A2(new_n416), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n361), .B1(new_n685), .B2(new_n415), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n435), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n592), .A2(new_n597), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n646), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n675), .A2(new_n690), .A3(new_n641), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n683), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n315), .B(KEYINPUT38), .Z(new_n693));
  OR2_X1    g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT107), .B(G143), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G45));
  NOR3_X1   g510(.A1(new_n634), .A2(new_n635), .A3(new_n668), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n676), .A2(new_n642), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n617), .B2(new_n503), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n617), .B2(KEYINPUT108), .ZN(new_n702));
  INV_X1    g516(.A(new_n479), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n478), .B1(new_n465), .B2(new_n477), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n483), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT84), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n496), .B1(new_n707), .B2(new_n491), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(G902), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n701), .B1(new_n702), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n617), .A2(KEYINPUT108), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n709), .B1(new_n708), .B2(G902), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n700), .A4(G469), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n457), .A3(new_n461), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n637), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT41), .B(G113), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  AOI21_X1  g533(.A(new_n460), .B1(new_n711), .B2(new_n714), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n647), .A2(new_n602), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n642), .A3(new_n457), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  AOI21_X1  g537(.A(new_n657), .B1(new_n435), .B2(new_n456), .ZN(new_n724));
  INV_X1    g538(.A(new_n604), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n720), .A2(new_n642), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n418), .B(new_n428), .C1(new_n415), .C2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n430), .B(KEYINPUT110), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND4_X1   g546(.A1(new_n374), .A2(new_n614), .A3(new_n603), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n715), .A2(new_n461), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n690), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n315), .A2(new_n606), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n728), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n641), .B(new_n690), .C1(new_n313), .C2(new_n314), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(KEYINPUT111), .A3(new_n720), .A4(new_n733), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  AND2_X1   g555(.A1(new_n614), .A2(new_n732), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n675), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n720), .A2(new_n743), .A3(new_n642), .A4(new_n697), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  AND3_X1   g559(.A1(new_n313), .A2(new_n314), .A3(new_n606), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n502), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n500), .A2(KEYINPUT112), .A3(new_n501), .A4(G469), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n748), .A2(new_n505), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n460), .B1(new_n750), .B2(new_n618), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n746), .A2(new_n697), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n674), .A2(new_n374), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT113), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n674), .A2(new_n755), .A3(new_n374), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT42), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n313), .A2(new_n751), .A3(new_n314), .A4(new_n606), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n753), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n697), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n389), .ZN(G33));
  NAND4_X1  g578(.A1(new_n746), .A2(new_n457), .A3(new_n669), .A4(new_n751), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  AND2_X1   g580(.A1(new_n500), .A2(new_n501), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n767), .A2(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(KEYINPUT45), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(G469), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n504), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(KEYINPUT46), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n618), .B1(new_n773), .B2(KEYINPUT46), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n461), .B(new_n681), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT43), .B1(new_n635), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n628), .A2(new_n633), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n635), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n779), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n621), .A2(new_n657), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n782), .A2(KEYINPUT44), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT44), .B1(new_n782), .B2(new_n783), .ZN(new_n785));
  INV_X1    g599(.A(new_n746), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n777), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  OAI21_X1  g603(.A(new_n461), .B1(new_n774), .B2(new_n775), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT47), .B(new_n461), .C1(new_n774), .C2(new_n775), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n634), .A2(new_n635), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n667), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n674), .A3(new_n374), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(new_n746), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  XOR2_X1   g613(.A(new_n715), .B(KEYINPUT116), .Z(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT49), .Z(new_n801));
  INV_X1    g615(.A(new_n688), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n781), .A2(new_n375), .A3(new_n607), .A4(new_n460), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n801), .A2(new_n693), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n782), .A2(new_n599), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n742), .A2(new_n374), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n786), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n800), .A2(new_n461), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n808), .B1(new_n794), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n720), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n786), .A2(new_n811), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n374), .A2(new_n812), .A3(new_n599), .A4(new_n802), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n635), .A3(new_n634), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n805), .A2(new_n812), .A3(new_n743), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n807), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n641), .A3(new_n693), .A4(new_n720), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n810), .B(new_n816), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT119), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n678), .A2(new_n676), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n677), .B1(new_n642), .B2(new_n669), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n698), .B(new_n744), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n688), .A2(new_n657), .A3(new_n667), .A4(new_n751), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n736), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT52), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n744), .A2(new_n698), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  INV_X1    g647(.A(new_n830), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n832), .A2(new_n679), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n722), .A2(new_n726), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n609), .B1(new_n716), .B2(new_n637), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n653), .A2(new_n616), .A3(new_n622), .A4(new_n636), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n740), .A2(new_n837), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n597), .A2(new_n645), .A3(new_n555), .A4(new_n667), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n674), .A2(new_n842), .A3(new_n620), .A4(new_n675), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n760), .A2(new_n669), .B1(new_n843), .B2(new_n746), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n746), .A2(new_n743), .A3(new_n697), .A4(new_n751), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n758), .A2(new_n844), .A3(new_n762), .A4(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n689), .A2(new_n602), .A3(new_n555), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n653), .A2(new_n616), .A3(new_n622), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n659), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT117), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n848), .A2(new_n851), .A3(new_n659), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n841), .A2(new_n846), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n836), .A2(new_n854), .A3(KEYINPUT53), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n843), .A2(new_n746), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n765), .A2(new_n845), .A3(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n674), .A2(new_n755), .A3(new_n374), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n755), .B1(new_n674), .B2(new_n374), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n759), .A2(new_n796), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n761), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n759), .A2(new_n796), .A3(new_n753), .A4(KEYINPUT42), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n858), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n722), .A2(new_n726), .ZN(new_n866));
  INV_X1    g680(.A(new_n840), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n866), .A2(new_n838), .A3(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n848), .A2(new_n851), .A3(new_n659), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n851), .B1(new_n848), .B2(new_n659), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(new_n740), .A3(new_n868), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n831), .A2(new_n835), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n856), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n855), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n836), .A2(new_n854), .A3(KEYINPUT118), .A4(KEYINPUT53), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n855), .A2(new_n874), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n805), .A2(new_n812), .A3(new_n861), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT48), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n807), .A2(new_n643), .A3(new_n811), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n598), .B(new_n885), .C1(new_n795), .C2(new_n813), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n884), .B(new_n886), .C1(new_n822), .C2(new_n823), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n825), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n804), .B1(new_n888), .B2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n411), .A2(G952), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n305), .B(new_n307), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT55), .Z(new_n893));
  NAND4_X1  g707(.A1(new_n876), .A2(G210), .A3(G902), .A4(new_n877), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n876), .A2(G902), .A3(new_n877), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n876), .A2(KEYINPUT120), .A3(G902), .A4(new_n877), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n312), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n893), .A2(new_n895), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n891), .B(new_n896), .C1(new_n901), .C2(new_n902), .ZN(G51));
  NAND3_X1  g717(.A1(new_n876), .A2(KEYINPUT54), .A3(new_n877), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n876), .A2(KEYINPUT121), .A3(KEYINPUT54), .A4(new_n877), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n880), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n504), .B(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n708), .B(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n899), .A2(new_n900), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n772), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n891), .B1(new_n912), .B2(new_n914), .ZN(G54));
  AND2_X1   g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n913), .A2(KEYINPUT123), .A3(new_n589), .A4(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n899), .A2(new_n900), .A3(new_n916), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n585), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n891), .B1(new_n919), .B2(new_n585), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(G60));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT59), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n908), .A2(new_n631), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n881), .A2(new_n879), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT54), .B1(new_n876), .B2(new_n877), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n631), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n891), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n925), .A2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n359), .B1(new_n878), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n891), .ZN(new_n935));
  INV_X1    g749(.A(new_n933), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n876), .A2(new_n656), .A3(new_n877), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT61), .B1(new_n937), .B2(KEYINPUT124), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G66));
  OAI21_X1  g754(.A(G953), .B1(new_n601), .B2(new_n187), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n841), .A2(new_n853), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(G953), .ZN(new_n943));
  INV_X1    g757(.A(new_n305), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(G898), .B2(new_n411), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT125), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n943), .B(new_n946), .ZN(G69));
  OAI21_X1  g761(.A(new_n397), .B1(new_n406), .B2(new_n407), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n565), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n795), .B1(new_n635), .B2(new_n646), .ZN(new_n950));
  OR4_X1    g764(.A1(new_n753), .A2(new_n786), .A3(new_n682), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n788), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n694), .A2(new_n679), .A3(new_n832), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n954), .A2(new_n798), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n949), .B1(new_n958), .B2(new_n411), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n949), .B1(new_n664), .B2(new_n411), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n777), .A2(new_n738), .A3(new_n861), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n798), .A2(new_n765), .A3(new_n788), .A4(new_n961), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n962), .A2(new_n763), .A3(new_n828), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n963), .B2(new_n411), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n411), .B1(G227), .B2(G900), .ZN(new_n965));
  OR3_X1    g779(.A1(new_n959), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n959), .B2(new_n964), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G72));
  INV_X1    g782(.A(new_n684), .ZN(new_n969));
  INV_X1    g783(.A(new_n942), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n958), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  AOI21_X1  g787(.A(new_n969), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n436), .A2(new_n419), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n969), .A2(new_n975), .A3(new_n973), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n881), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n973), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n963), .B2(new_n942), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n975), .B(KEYINPUT127), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n935), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n974), .A2(new_n977), .A3(new_n981), .ZN(G57));
endmodule


