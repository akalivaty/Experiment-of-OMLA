//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  INV_X1    g033(.A(new_n452), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n463), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n467), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(new_n465), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n469), .A2(new_n470), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n467), .A2(new_n468), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NOR2_X1   g061(.A1(new_n482), .A2(new_n479), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n479), .A2(G2105), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n487), .A2(G124), .B1(new_n488), .B2(G136), .ZN(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n482), .C2(G112), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OR2_X1    g067(.A1(new_n463), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n479), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n469), .A2(new_n470), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n482), .A2(new_n499), .A3(new_n500), .A4(G138), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT4), .B1(new_n471), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n506), .A2(new_n509), .A3(G62), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n505), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT5), .B(G543), .Z(new_n513));
  AND3_X1   g088(.A1(KEYINPUT69), .A2(KEYINPUT6), .A3(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT6), .B1(KEYINPUT69), .B2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(G543), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n517), .A2(G88), .B1(new_n519), .B2(G50), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n520), .B1(new_n511), .B2(KEYINPUT71), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n512), .A2(new_n521), .ZN(G166));
  AND2_X1   g097(.A1(new_n517), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n525), .B(new_n526), .C1(new_n518), .C2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n523), .A2(new_n528), .ZN(G168));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  INV_X1    g105(.A(G77), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n513), .A2(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI221_X1 g110(.A(KEYINPUT72), .B1(new_n531), .B2(new_n532), .C1(new_n513), .C2(new_n530), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(G651), .A3(new_n536), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT73), .B(G52), .Z(new_n538));
  AOI22_X1  g113(.A1(new_n517), .A2(G90), .B1(new_n519), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n505), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n519), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n517), .A2(G81), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT75), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  AOI22_X1  g130(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n505), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT76), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n518), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n518), .B2(new_n559), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n560), .A2(new_n561), .B1(G91), .B2(new_n517), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n517), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n519), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n519), .A2(G48), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n513), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(G651), .A2(new_n575), .B1(new_n517), .B2(G86), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(G72), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G60), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n513), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n505), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n582), .B1(new_n581), .B2(new_n580), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n517), .A2(G85), .B1(new_n519), .B2(G47), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(new_n517), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n513), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n519), .B2(G54), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(G868), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g169(.A(new_n593), .B1(G171), .B2(G868), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  AND2_X1   g174(.A1(new_n587), .A2(new_n591), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT79), .B(G559), .Z(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(G860), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT80), .ZN(G148));
  NOR2_X1   g178(.A1(new_n548), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n601), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT81), .Z(new_n606));
  AOI21_X1  g181(.A(new_n604), .B1(new_n606), .B2(G868), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n499), .A2(new_n464), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  OAI221_X1 g189(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n482), .C2(G111), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n487), .A2(G123), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n488), .A2(G135), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2096), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n626), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2443), .B(G2446), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT82), .ZN(new_n634));
  OAI21_X1  g209(.A(G14), .B1(new_n631), .B2(new_n632), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(G401));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT83), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2072), .B(G2078), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT84), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT86), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT85), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(KEYINPUT18), .ZN(new_n647));
  OAI21_X1  g222(.A(KEYINPUT17), .B1(new_n638), .B2(new_n639), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(new_n642), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n642), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n640), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2096), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT20), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n656), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n656), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT87), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G229));
  NOR2_X1   g248(.A1(G16), .A2(G19), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n549), .B2(G16), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1341), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G4), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n600), .B2(new_n678), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n680), .A2(G1348), .ZN(new_n681));
  INV_X1    g256(.A(G29), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G26), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT28), .Z(new_n684));
  AOI22_X1  g259(.A1(new_n487), .A2(G128), .B1(new_n488), .B2(G140), .ZN(new_n685));
  NOR2_X1   g260(.A1(G104), .A2(G2105), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT93), .ZN(new_n687));
  OAI21_X1  g262(.A(G2104), .B1(new_n482), .B2(G116), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n684), .B1(new_n689), .B2(G29), .ZN(new_n690));
  INV_X1    g265(.A(G2067), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n680), .A2(G1348), .ZN(new_n693));
  NOR4_X1   g268(.A1(new_n677), .A2(new_n681), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT94), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n678), .A2(G20), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT23), .Z(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G299), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1956), .ZN(new_n699));
  NOR2_X1   g274(.A1(G171), .A2(new_n678), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G5), .B2(new_n678), .ZN(new_n701));
  INV_X1    g276(.A(G1961), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n702), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT31), .B(G11), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT30), .B(G28), .Z(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n618), .A2(G29), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(KEYINPUT99), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n678), .A2(G21), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G168), .B2(new_n678), .ZN(new_n711));
  OAI221_X1 g286(.A(new_n709), .B1(KEYINPUT99), .B2(new_n708), .C1(new_n711), .C2(G1966), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n682), .A2(G32), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n487), .A2(G129), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT96), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT97), .B(KEYINPUT26), .ZN(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n716), .B(new_n717), .Z(new_n718));
  AND2_X1   g293(.A1(new_n464), .A2(G105), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n488), .B2(G141), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n715), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n713), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT27), .B(G1996), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n712), .B(new_n724), .C1(G1966), .C2(new_n711), .ZN(new_n725));
  INV_X1    g300(.A(G2090), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n682), .A2(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n682), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT29), .Z(new_n729));
  OAI21_X1  g304(.A(new_n725), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n726), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g307(.A1(KEYINPUT24), .A2(G34), .ZN(new_n733));
  NOR2_X1   g308(.A1(KEYINPUT24), .A2(G34), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n485), .A2(G29), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT100), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n682), .A2(G27), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G164), .B2(new_n682), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT101), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G2078), .Z(new_n743));
  NOR4_X1   g318(.A1(new_n730), .A2(new_n732), .A3(new_n739), .A4(new_n743), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n682), .A2(G33), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT25), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n488), .A2(G139), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n747), .B(new_n748), .C1(new_n482), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n745), .B1(new_n750), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G2072), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT95), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n722), .A2(new_n723), .B1(new_n751), .B2(new_n752), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n754), .B(new_n755), .C1(new_n737), .C2(new_n736), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT98), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n695), .A2(new_n704), .A3(new_n744), .A4(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G305), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G16), .ZN(new_n760));
  OR2_X1    g335(.A1(G6), .A2(G16), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(KEYINPUT32), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n760), .A2(new_n764), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G1981), .ZN(new_n767));
  INV_X1    g342(.A(G1981), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n763), .A2(new_n768), .A3(new_n765), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(G166), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G16), .B2(G22), .ZN(new_n772));
  INV_X1    g347(.A(G1971), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n678), .A2(G23), .ZN(new_n775));
  INV_X1    g350(.A(G288), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n678), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT33), .B(G1976), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n777), .B(new_n778), .Z(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n773), .B2(new_n772), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n770), .A2(new_n774), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n770), .A2(KEYINPUT89), .A3(new_n774), .A4(new_n780), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n783), .A2(KEYINPUT34), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n783), .A2(KEYINPUT90), .A3(KEYINPUT34), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(KEYINPUT34), .B1(new_n783), .B2(new_n784), .ZN(new_n790));
  INV_X1    g365(.A(G290), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(new_n678), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n678), .B2(G24), .ZN(new_n793));
  INV_X1    g368(.A(G1986), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n487), .A2(G119), .B1(new_n488), .B2(G131), .ZN(new_n797));
  OAI221_X1 g372(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n482), .C2(G107), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G25), .B(new_n799), .S(G29), .Z(new_n800));
  XOR2_X1   g375(.A(KEYINPUT35), .B(G1991), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n795), .A2(new_n796), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n790), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n789), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT91), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n808), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n789), .A2(new_n810), .A3(new_n804), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n758), .B1(new_n809), .B2(new_n811), .ZN(G311));
  INV_X1    g387(.A(new_n758), .ZN(new_n813));
  INV_X1    g388(.A(new_n811), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n810), .B1(new_n789), .B2(new_n804), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(G150));
  NAND2_X1  g391(.A1(new_n517), .A2(G93), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n519), .A2(G55), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n817), .B(new_n818), .C1(new_n505), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G860), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n600), .A2(G559), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT103), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n548), .B(new_n820), .Z(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n828), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n822), .B1(new_n837), .B2(new_n838), .ZN(G145));
  NAND2_X1  g414(.A1(new_n501), .A2(new_n503), .ZN(new_n840));
  INV_X1    g415(.A(new_n498), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n689), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n721), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n750), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n487), .A2(G130), .B1(new_n488), .B2(G142), .ZN(new_n846));
  OAI221_X1 g421(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n482), .C2(G118), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n610), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n799), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT105), .B1(new_n845), .B2(new_n850), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n485), .B(new_n618), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n491), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(KEYINPUT106), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n856), .A2(KEYINPUT106), .ZN(new_n860));
  AOI211_X1 g435(.A(new_n859), .B(new_n860), .C1(new_n850), .C2(new_n845), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n852), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT40), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n854), .A2(new_n857), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT40), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n867), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(G395));
  NAND2_X1  g445(.A1(new_n600), .A2(new_n597), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n592), .A2(G299), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT41), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT107), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n873), .B(KEYINPUT41), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(KEYINPUT107), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n606), .B(new_n827), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n873), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n881), .B2(new_n879), .ZN(new_n882));
  NAND2_X1  g457(.A1(G303), .A2(G305), .ZN(new_n883));
  NAND2_X1  g458(.A1(G166), .A2(new_n759), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(new_n776), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n883), .B(new_n884), .C1(KEYINPUT108), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(KEYINPUT108), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT42), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n882), .B(new_n889), .ZN(new_n890));
  MUX2_X1   g465(.A(new_n820), .B(new_n890), .S(G868), .Z(G295));
  MUX2_X1   g466(.A(new_n820), .B(new_n890), .S(G868), .Z(G331));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n893));
  XNOR2_X1  g468(.A(G301), .B(G168), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n894), .A2(new_n826), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n826), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(new_n876), .C1(KEYINPUT107), .C2(new_n877), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n881), .A3(new_n896), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n888), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n863), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n888), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n893), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n877), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT109), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n905), .A3(new_n899), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n899), .A2(new_n905), .ZN(new_n907));
  INV_X1    g482(.A(new_n888), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(KEYINPUT43), .A3(new_n863), .A4(new_n900), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT44), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n901), .B2(new_n902), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n909), .A2(new_n893), .A3(new_n863), .A4(new_n900), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n912), .A2(new_n917), .ZN(G397));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(G164), .B2(G1384), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n474), .A2(G40), .A3(new_n484), .A4(new_n476), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n721), .B(G1996), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n689), .B(G2067), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n799), .B(new_n801), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n925), .B(new_n926), .C1(new_n794), .C2(new_n791), .ZN(new_n927));
  NOR2_X1   g502(.A1(G290), .A2(G1986), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT110), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT62), .ZN(new_n931));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n842), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AND4_X1   g509(.A1(G40), .A2(new_n474), .A3(new_n484), .A4(new_n476), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n936));
  AND4_X1   g511(.A1(new_n737), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n919), .A2(G1384), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n840), .B2(new_n841), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(new_n921), .ZN(new_n941));
  AOI21_X1  g516(.A(G1966), .B1(new_n941), .B2(new_n920), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT123), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(KEYINPUT116), .B(G8), .ZN(new_n944));
  NOR2_X1   g519(.A1(G168), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n842), .A2(new_n938), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n935), .A2(new_n920), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1966), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT123), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n737), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n943), .A2(new_n945), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n943), .A2(G8), .A3(new_n952), .ZN(new_n955));
  INV_X1    g530(.A(new_n945), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n949), .A2(new_n951), .ZN(new_n958));
  INV_X1    g533(.A(new_n944), .ZN(new_n959));
  AOI211_X1 g534(.A(KEYINPUT51), .B(new_n945), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n931), .B(new_n953), .C1(new_n957), .C2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT53), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(G164), .B2(new_n939), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n920), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n842), .A2(KEYINPUT111), .A3(new_n938), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n935), .A4(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n935), .A3(new_n920), .A4(new_n964), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT112), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n962), .B1(new_n971), .B2(G2078), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n702), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n962), .A2(G2078), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n947), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT124), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n974), .B(new_n979), .C1(new_n947), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G301), .B1(new_n972), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n961), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n842), .A2(new_n932), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(new_n921), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(new_n944), .ZN(new_n986));
  INV_X1    g561(.A(G1976), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(new_n987), .B2(G288), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT52), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT49), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n572), .A2(new_n768), .A3(new_n576), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n768), .B1(new_n572), .B2(new_n576), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n993), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(KEYINPUT49), .A3(new_n991), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n996), .A3(new_n986), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(G288), .B2(new_n987), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n986), .B(new_n998), .C1(new_n987), .C2(G288), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n989), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n968), .A2(new_n773), .A3(new_n970), .ZN(new_n1001));
  INV_X1    g576(.A(new_n933), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(G164), .B2(G1384), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n935), .B(new_n1003), .C1(new_n984), .C2(KEYINPUT50), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(G2090), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n959), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(G166), .B2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(KEYINPUT55), .B(G8), .C1(new_n512), .C2(new_n521), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1000), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n973), .A2(G2090), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1001), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT114), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1010), .A2(KEYINPUT115), .A3(new_n1011), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT115), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1001), .A2(new_n1020), .A3(new_n1014), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1016), .A2(new_n1019), .A3(G8), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT126), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1013), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n1013), .B2(new_n1022), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n983), .B(KEYINPUT127), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n953), .B1(new_n957), .B2(new_n960), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1013), .A2(new_n1022), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT126), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1013), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT127), .B1(new_n1033), .B2(new_n983), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1016), .A2(G8), .A3(new_n1021), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1012), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n958), .A2(G168), .A3(new_n959), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1000), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1036), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1039), .A2(KEYINPUT63), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1000), .B1(new_n1044), .B2(new_n1022), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n986), .B(KEYINPUT117), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n997), .A2(new_n987), .A3(new_n776), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n991), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1041), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT119), .B1(new_n560), .B2(new_n561), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(KEYINPUT57), .ZN(new_n1051));
  XNOR2_X1  g626(.A(G299), .B(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT56), .B(G2072), .Z(new_n1053));
  OR2_X1    g628(.A1(new_n969), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1956), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1004), .A2(KEYINPUT118), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT118), .B1(new_n1004), .B2(new_n1055), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1052), .B(new_n1054), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G164), .A2(G1384), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n935), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT120), .B1(new_n1061), .B2(G2067), .ZN(new_n1062));
  INV_X1    g637(.A(G1348), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n973), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n985), .A2(new_n1065), .A3(new_n691), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n600), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1059), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1004), .A2(new_n1055), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1004), .A2(KEYINPUT118), .A3(new_n1055), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1052), .B1(new_n1074), .B2(new_n1054), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n592), .A2(KEYINPUT60), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1077), .A2(new_n1062), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND2_X1  g654(.A1(new_n1061), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n969), .B2(G1996), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n549), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1081), .B2(new_n549), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1078), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .A4(new_n592), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1068), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1075), .B2(new_n1059), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1058), .B1(new_n1075), .B2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1074), .A2(KEYINPUT121), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(KEYINPUT61), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1092), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1095), .A2(new_n1096), .A3(KEYINPUT122), .A4(KEYINPUT61), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1076), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n965), .A2(new_n967), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n482), .B1(new_n481), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1103), .B2(new_n481), .ZN(new_n1105));
  AND4_X1   g680(.A1(G40), .A2(new_n477), .A3(new_n975), .A4(new_n1105), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1102), .A2(new_n1106), .B1(new_n973), .B2(new_n702), .ZN(new_n1107));
  AOI21_X1  g682(.A(G2078), .B1(new_n968), .B2(new_n970), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(KEYINPUT53), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1101), .B1(new_n1109), .B2(G171), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n972), .A2(G301), .A3(new_n981), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1112), .A2(new_n1027), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n972), .A2(G301), .A3(new_n1107), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1101), .B1(new_n1115), .B2(new_n982), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1113), .B(new_n1116), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1049), .B1(new_n1100), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n930), .B1(new_n1035), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n925), .A2(new_n926), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n929), .A2(new_n922), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1120), .A2(new_n922), .B1(KEYINPUT48), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(KEYINPUT48), .B2(new_n1122), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n925), .A2(new_n801), .A3(new_n798), .A4(new_n797), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(G2067), .B2(new_n689), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n922), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n922), .B1(new_n924), .B2(new_n721), .ZN(new_n1128));
  NOR4_X1   g703(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT46), .A4(G1996), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT46), .ZN(new_n1130));
  INV_X1    g705(.A(G1996), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1130), .B1(new_n922), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1128), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT47), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1124), .A2(new_n1127), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1119), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g711(.A1(new_n858), .A2(new_n865), .ZN(new_n1138));
  NOR4_X1   g712(.A1(G401), .A2(G227), .A3(G229), .A4(new_n461), .ZN(new_n1139));
  AND3_X1   g713(.A1(new_n1138), .A2(new_n915), .A3(new_n1139), .ZN(G308));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n915), .A3(new_n1139), .ZN(G225));
endmodule


