

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779;

  OR2_X1 U376 ( .A1(n531), .A2(n557), .ZN(n565) );
  XNOR2_X1 U377 ( .A(n406), .B(KEYINPUT64), .ZN(n405) );
  INV_X1 U378 ( .A(G953), .ZN(n772) );
  XNOR2_X2 U379 ( .A(n409), .B(KEYINPUT40), .ZN(n533) );
  NAND2_X2 U380 ( .A1(n373), .A2(n371), .ZN(n556) );
  NOR2_X1 U381 ( .A1(n537), .A2(n589), .ZN(n549) );
  NAND2_X1 U382 ( .A1(n395), .A2(n392), .ZN(n632) );
  AND2_X1 U383 ( .A1(n396), .A2(n631), .ZN(n395) );
  XNOR2_X1 U384 ( .A(n603), .B(n602), .ZN(n628) );
  OR2_X1 U385 ( .A1(n529), .A2(n566), .ZN(n701) );
  XNOR2_X1 U386 ( .A(n376), .B(n536), .ZN(n589) );
  AND2_X1 U387 ( .A1(n375), .A2(n374), .ZN(n373) );
  OR2_X1 U388 ( .A1(n667), .A2(G902), .ZN(n519) );
  XNOR2_X2 U389 ( .A(n469), .B(n419), .ZN(n516) );
  XNOR2_X2 U390 ( .A(n590), .B(KEYINPUT0), .ZN(n591) );
  NOR2_X1 U391 ( .A1(n369), .A2(n564), .ZN(n576) );
  XNOR2_X1 U392 ( .A(n370), .B(KEYINPUT39), .ZN(n583) );
  NOR2_X1 U393 ( .A1(n577), .A2(KEYINPUT48), .ZN(n389) );
  NAND2_X1 U394 ( .A1(n615), .A2(KEYINPUT86), .ZN(n397) );
  OR2_X1 U395 ( .A1(n432), .A2(n634), .ZN(n372) );
  OR2_X1 U396 ( .A1(n681), .A2(n682), .ZN(n685) );
  XNOR2_X1 U397 ( .A(n469), .B(n477), .ZN(n649) );
  INV_X1 U398 ( .A(G110), .ZN(n417) );
  XNOR2_X1 U399 ( .A(n463), .B(n462), .ZN(n464) );
  NAND2_X1 U400 ( .A1(n362), .A2(n354), .ZN(n377) );
  XNOR2_X1 U401 ( .A(n468), .B(KEYINPUT41), .ZN(n713) );
  NOR2_X1 U402 ( .A1(n701), .A2(n700), .ZN(n468) );
  AND2_X1 U403 ( .A1(n620), .A2(n528), .ZN(n561) );
  AND2_X1 U404 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U405 ( .A(n639), .B(KEYINPUT89), .ZN(n677) );
  XNOR2_X1 U406 ( .A(n391), .B(KEYINPUT83), .ZN(n584) );
  NAND2_X1 U407 ( .A1(n386), .A2(n385), .ZN(n391) );
  AND2_X1 U408 ( .A1(n388), .A2(n358), .ZN(n386) );
  NAND2_X1 U409 ( .A1(n401), .A2(n366), .ZN(n381) );
  NAND2_X1 U410 ( .A1(n432), .A2(n634), .ZN(n374) );
  XNOR2_X1 U411 ( .A(G137), .B(KEYINPUT5), .ZN(n471) );
  XNOR2_X1 U412 ( .A(KEYINPUT3), .B(G119), .ZN(n420) );
  XOR2_X1 U413 ( .A(G113), .B(G116), .Z(n421) );
  XNOR2_X1 U414 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U415 ( .A(G116), .B(G134), .ZN(n451) );
  NOR2_X1 U416 ( .A1(G953), .A2(G237), .ZN(n470) );
  XOR2_X1 U417 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n437) );
  NAND2_X1 U418 ( .A1(G234), .A2(G237), .ZN(n485) );
  OR2_X1 U419 ( .A1(n619), .A2(n566), .ZN(n525) );
  INV_X1 U420 ( .A(n410), .ZN(n771) );
  XNOR2_X1 U421 ( .A(G119), .B(G110), .ZN(n491) );
  XNOR2_X1 U422 ( .A(G128), .B(G146), .ZN(n493) );
  XNOR2_X1 U423 ( .A(G122), .B(G104), .ZN(n443) );
  XNOR2_X1 U424 ( .A(G125), .B(G140), .ZN(n439) );
  XNOR2_X1 U425 ( .A(G143), .B(G146), .ZN(n441) );
  XOR2_X1 U426 ( .A(G131), .B(G113), .Z(n442) );
  INV_X1 U427 ( .A(G134), .ZN(n473) );
  XNOR2_X1 U428 ( .A(KEYINPUT73), .B(G137), .ZN(n512) );
  XNOR2_X1 U429 ( .A(G104), .B(G140), .ZN(n511) );
  NOR2_X1 U430 ( .A1(n685), .A2(n572), .ZN(n523) );
  XNOR2_X1 U431 ( .A(n591), .B(KEYINPUT92), .ZN(n622) );
  XNOR2_X1 U432 ( .A(n384), .B(n364), .ZN(n534) );
  OR2_X1 U433 ( .A1(n713), .A2(n537), .ZN(n384) );
  AND2_X1 U434 ( .A1(n574), .A2(n605), .ZN(n646) );
  INV_X1 U435 ( .A(n693), .ZN(n399) );
  AND2_X1 U436 ( .A1(n628), .A2(n402), .ZN(n736) );
  NOR2_X1 U437 ( .A1(n359), .A2(n403), .ZN(n402) );
  INV_X1 U438 ( .A(n681), .ZN(n403) );
  XNOR2_X1 U439 ( .A(n565), .B(KEYINPUT107), .ZN(n745) );
  INV_X1 U440 ( .A(n677), .ZN(n640) );
  XNOR2_X1 U441 ( .A(n637), .B(n365), .ZN(n641) );
  INV_X1 U442 ( .A(G122), .ZN(n408) );
  AND2_X1 U443 ( .A1(n584), .A2(n363), .ZN(n353) );
  AND2_X1 U444 ( .A1(n411), .A2(n367), .ZN(n354) );
  AND2_X1 U445 ( .A1(n634), .A2(n633), .ZN(n355) );
  AND2_X1 U446 ( .A1(n745), .A2(n413), .ZN(n356) );
  XOR2_X1 U447 ( .A(KEYINPUT72), .B(KEYINPUT10), .Z(n357) );
  AND2_X1 U448 ( .A1(n387), .A2(n644), .ZN(n358) );
  NAND2_X1 U449 ( .A1(n686), .A2(n619), .ZN(n359) );
  AND2_X1 U450 ( .A1(n381), .A2(n411), .ZN(n360) );
  NOR2_X1 U451 ( .A1(n700), .A2(n682), .ZN(n361) );
  AND2_X1 U452 ( .A1(n382), .A2(n381), .ZN(n362) );
  AND2_X1 U453 ( .A1(n643), .A2(n412), .ZN(n363) );
  XOR2_X1 U454 ( .A(n522), .B(KEYINPUT42), .Z(n364) );
  XNOR2_X1 U455 ( .A(n609), .B(n608), .ZN(n648) );
  XOR2_X1 U456 ( .A(n636), .B(n635), .Z(n365) );
  XNOR2_X1 U457 ( .A(n516), .B(n429), .ZN(n672) );
  INV_X1 U458 ( .A(KEYINPUT66), .ZN(n400) );
  NAND2_X1 U459 ( .A1(n720), .A2(KEYINPUT2), .ZN(n366) );
  AND2_X1 U460 ( .A1(n355), .A2(KEYINPUT66), .ZN(n367) );
  NAND2_X1 U461 ( .A1(G898), .A2(KEYINPUT61), .ZN(n368) );
  NAND2_X1 U462 ( .A1(n533), .A2(n534), .ZN(n535) );
  NAND2_X1 U463 ( .A1(n563), .A2(n741), .ZN(n369) );
  XNOR2_X1 U464 ( .A(n508), .B(KEYINPUT28), .ZN(n521) );
  NAND2_X1 U465 ( .A1(n561), .A2(n698), .ZN(n370) );
  OR2_X1 U466 ( .A1(n672), .A2(n372), .ZN(n371) );
  NAND2_X1 U467 ( .A1(n672), .A2(n432), .ZN(n375) );
  NAND2_X1 U468 ( .A1(n556), .A2(n697), .ZN(n376) );
  NAND2_X2 U469 ( .A1(n378), .A2(n377), .ZN(n671) );
  NAND2_X1 U470 ( .A1(n379), .A2(n400), .ZN(n378) );
  NAND2_X1 U471 ( .A1(n360), .A2(n380), .ZN(n379) );
  AND2_X1 U472 ( .A1(n382), .A2(n355), .ZN(n380) );
  NAND2_X1 U473 ( .A1(n410), .A2(n366), .ZN(n382) );
  INV_X1 U474 ( .A(n383), .ZN(n401) );
  NAND2_X1 U475 ( .A1(n353), .A2(n383), .ZN(n411) );
  XNOR2_X2 U476 ( .A(n632), .B(KEYINPUT45), .ZN(n383) );
  AND2_X1 U477 ( .A1(n401), .A2(n368), .ZN(n750) );
  AND2_X1 U478 ( .A1(n771), .A2(n383), .ZN(n717) );
  INV_X1 U479 ( .A(n534), .ZN(n779) );
  NAND2_X1 U480 ( .A1(n578), .A2(KEYINPUT48), .ZN(n385) );
  NAND2_X1 U481 ( .A1(n577), .A2(KEYINPUT48), .ZN(n387) );
  NAND2_X1 U482 ( .A1(n390), .A2(n389), .ZN(n388) );
  INV_X1 U483 ( .A(n578), .ZN(n390) );
  NAND2_X1 U484 ( .A1(n393), .A2(n613), .ZN(n392) );
  NAND2_X1 U485 ( .A1(n394), .A2(n611), .ZN(n393) );
  NAND2_X1 U486 ( .A1(n601), .A2(KEYINPUT86), .ZN(n394) );
  NAND2_X1 U487 ( .A1(n398), .A2(n397), .ZN(n396) );
  INV_X1 U488 ( .A(n601), .ZN(n398) );
  NAND2_X1 U489 ( .A1(n591), .A2(n361), .ZN(n603) );
  NAND2_X1 U490 ( .A1(n591), .A2(n399), .ZN(n618) );
  NAND2_X1 U491 ( .A1(n628), .A2(n404), .ZN(n609) );
  AND2_X1 U492 ( .A1(n606), .A2(n681), .ZN(n404) );
  XNOR2_X2 U493 ( .A(n459), .B(n405), .ZN(n770) );
  XNOR2_X2 U494 ( .A(KEYINPUT4), .B(G146), .ZN(n406) );
  XNOR2_X2 U495 ( .A(n407), .B(G128), .ZN(n459) );
  XNOR2_X2 U496 ( .A(G143), .B(KEYINPUT65), .ZN(n407) );
  XNOR2_X1 U497 ( .A(n601), .B(n408), .ZN(G24) );
  XNOR2_X2 U498 ( .A(n600), .B(KEYINPUT35), .ZN(n601) );
  INV_X1 U499 ( .A(n533), .ZN(n647) );
  NAND2_X1 U500 ( .A1(n583), .A2(n532), .ZN(n409) );
  NAND2_X1 U501 ( .A1(n584), .A2(n643), .ZN(n410) );
  INV_X1 U502 ( .A(n366), .ZN(n412) );
  AND2_X1 U503 ( .A1(n568), .A2(n625), .ZN(n413) );
  XOR2_X1 U504 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n414) );
  AND2_X1 U505 ( .A1(G214), .A2(n470), .ZN(n415) );
  INV_X1 U506 ( .A(n697), .ZN(n566) );
  NOR2_X1 U507 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U508 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U509 ( .A(n438), .B(n415), .ZN(n440) );
  XNOR2_X1 U510 ( .A(n440), .B(n499), .ZN(n447) );
  BUF_X1 U511 ( .A(n556), .Z(n580) );
  XNOR2_X1 U512 ( .A(KEYINPUT70), .B(G101), .ZN(n416) );
  XNOR2_X2 U513 ( .A(n770), .B(n416), .ZN(n469) );
  XNOR2_X1 U514 ( .A(n417), .B(G107), .ZN(n757) );
  XNOR2_X1 U515 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n418) );
  XNOR2_X1 U516 ( .A(n757), .B(n418), .ZN(n419) );
  XNOR2_X1 U517 ( .A(n421), .B(n420), .ZN(n476) );
  XNOR2_X1 U518 ( .A(n443), .B(KEYINPUT16), .ZN(n422) );
  XNOR2_X1 U519 ( .A(n476), .B(n422), .ZN(n758) );
  XOR2_X1 U520 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n424) );
  XNOR2_X1 U521 ( .A(G125), .B(KEYINPUT17), .ZN(n423) );
  XNOR2_X1 U522 ( .A(n424), .B(n423), .ZN(n427) );
  NAND2_X1 U523 ( .A1(n772), .A2(G224), .ZN(n425) );
  XNOR2_X1 U524 ( .A(n425), .B(KEYINPUT90), .ZN(n426) );
  XNOR2_X1 U525 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U526 ( .A(n758), .B(n428), .ZN(n429) );
  XNOR2_X1 U527 ( .A(G902), .B(KEYINPUT15), .ZN(n480) );
  INV_X1 U528 ( .A(n480), .ZN(n634) );
  NOR2_X1 U529 ( .A1(G237), .A2(G902), .ZN(n431) );
  INV_X1 U530 ( .A(KEYINPUT78), .ZN(n430) );
  XNOR2_X1 U531 ( .A(n431), .B(n430), .ZN(n433) );
  AND2_X1 U532 ( .A1(n433), .A2(G210), .ZN(n432) );
  XNOR2_X1 U533 ( .A(n556), .B(KEYINPUT38), .ZN(n529) );
  INV_X1 U534 ( .A(n433), .ZN(n435) );
  INV_X1 U535 ( .A(G214), .ZN(n434) );
  OR2_X1 U536 ( .A1(n435), .A2(n434), .ZN(n697) );
  XNOR2_X1 U537 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n449) );
  XNOR2_X1 U538 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n436) );
  XNOR2_X1 U539 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U540 ( .A(n357), .B(n439), .ZN(n499) );
  XNOR2_X1 U541 ( .A(n442), .B(n441), .ZN(n445) );
  XNOR2_X1 U542 ( .A(n443), .B(KEYINPUT100), .ZN(n444) );
  XNOR2_X1 U543 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U544 ( .A(n447), .B(n446), .ZN(n660) );
  NOR2_X1 U545 ( .A1(G902), .A2(n660), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U547 ( .A(n450), .B(G475), .ZN(n531) );
  XOR2_X1 U548 ( .A(G122), .B(G107), .Z(n452) );
  XNOR2_X1 U549 ( .A(n452), .B(n451), .ZN(n456) );
  XOR2_X1 U550 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n454) );
  XNOR2_X1 U551 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n453) );
  XNOR2_X1 U552 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U553 ( .A(n456), .B(n455), .ZN(n465) );
  NAND2_X1 U554 ( .A1(n772), .A2(G234), .ZN(n458) );
  XNOR2_X1 U555 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n457) );
  XNOR2_X1 U556 ( .A(n458), .B(n457), .ZN(n496) );
  NAND2_X1 U557 ( .A1(n496), .A2(G217), .ZN(n463) );
  INV_X1 U558 ( .A(n459), .ZN(n461) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n460) );
  XNOR2_X1 U560 ( .A(n465), .B(n464), .ZN(n636) );
  INV_X1 U561 ( .A(G902), .ZN(n501) );
  NAND2_X1 U562 ( .A1(n636), .A2(n501), .ZN(n467) );
  INV_X1 U563 ( .A(G478), .ZN(n466) );
  XNOR2_X1 U564 ( .A(n467), .B(n466), .ZN(n530) );
  NAND2_X1 U565 ( .A1(n531), .A2(n530), .ZN(n700) );
  NAND2_X1 U566 ( .A1(n470), .A2(G210), .ZN(n472) );
  XNOR2_X1 U567 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U568 ( .A(n473), .B(G131), .ZN(n766) );
  XNOR2_X1 U569 ( .A(n474), .B(n766), .ZN(n475) );
  XNOR2_X1 U570 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U571 ( .A1(n649), .A2(n501), .ZN(n479) );
  XNOR2_X1 U572 ( .A(G472), .B(KEYINPUT97), .ZN(n478) );
  XNOR2_X2 U573 ( .A(n479), .B(n478), .ZN(n619) );
  NAND2_X1 U574 ( .A1(G234), .A2(n480), .ZN(n481) );
  XNOR2_X1 U575 ( .A(KEYINPUT20), .B(n481), .ZN(n502) );
  NAND2_X1 U576 ( .A1(G221), .A2(n502), .ZN(n484) );
  INV_X1 U577 ( .A(KEYINPUT95), .ZN(n482) );
  XNOR2_X1 U578 ( .A(n482), .B(KEYINPUT21), .ZN(n483) );
  XNOR2_X1 U579 ( .A(n484), .B(n483), .ZN(n682) );
  XNOR2_X1 U580 ( .A(n485), .B(KEYINPUT14), .ZN(n488) );
  AND2_X1 U581 ( .A1(G953), .A2(G902), .ZN(n486) );
  NAND2_X1 U582 ( .A1(n488), .A2(n486), .ZN(n585) );
  XNOR2_X1 U583 ( .A(KEYINPUT108), .B(n585), .ZN(n487) );
  NOR2_X1 U584 ( .A1(G900), .A2(n487), .ZN(n489) );
  NAND2_X1 U585 ( .A1(G952), .A2(n488), .ZN(n709) );
  NOR2_X1 U586 ( .A1(n709), .A2(G953), .ZN(n587) );
  OR2_X1 U587 ( .A1(n489), .A2(n587), .ZN(n526) );
  INV_X1 U588 ( .A(n526), .ZN(n490) );
  NOR2_X1 U589 ( .A1(n682), .A2(n490), .ZN(n507) );
  XNOR2_X1 U590 ( .A(n414), .B(n491), .ZN(n495) );
  INV_X1 U591 ( .A(KEYINPUT24), .ZN(n492) );
  XNOR2_X1 U592 ( .A(n495), .B(n494), .ZN(n498) );
  NAND2_X1 U593 ( .A1(n496), .A2(G221), .ZN(n497) );
  XNOR2_X1 U594 ( .A(n498), .B(n497), .ZN(n500) );
  XNOR2_X1 U595 ( .A(n499), .B(n512), .ZN(n765) );
  XNOR2_X1 U596 ( .A(n500), .B(n765), .ZN(n655) );
  NAND2_X1 U597 ( .A1(n655), .A2(n501), .ZN(n506) );
  NAND2_X1 U598 ( .A1(G217), .A2(n502), .ZN(n504) );
  XNOR2_X1 U599 ( .A(KEYINPUT94), .B(KEYINPUT25), .ZN(n503) );
  XNOR2_X1 U600 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X2 U601 ( .A(n506), .B(n505), .ZN(n681) );
  NAND2_X1 U602 ( .A1(n507), .A2(n681), .ZN(n567) );
  NOR2_X1 U603 ( .A1(n619), .A2(n567), .ZN(n508) );
  NAND2_X1 U604 ( .A1(n772), .A2(G227), .ZN(n509) );
  XNOR2_X1 U605 ( .A(n509), .B(KEYINPUT80), .ZN(n510) );
  XNOR2_X1 U606 ( .A(n766), .B(n510), .ZN(n514) );
  XNOR2_X1 U607 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U608 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U609 ( .A(n516), .B(n515), .ZN(n667) );
  INV_X1 U610 ( .A(KEYINPUT74), .ZN(n517) );
  XNOR2_X1 U611 ( .A(n517), .B(G469), .ZN(n518) );
  XNOR2_X2 U612 ( .A(n519), .B(n518), .ZN(n572) );
  XNOR2_X1 U613 ( .A(n572), .B(KEYINPUT109), .ZN(n520) );
  NAND2_X1 U614 ( .A1(n521), .A2(n520), .ZN(n537) );
  INV_X1 U615 ( .A(KEYINPUT110), .ZN(n522) );
  XNOR2_X1 U616 ( .A(n523), .B(KEYINPUT96), .ZN(n620) );
  INV_X1 U617 ( .A(KEYINPUT30), .ZN(n524) );
  XNOR2_X1 U618 ( .A(n525), .B(n524), .ZN(n527) );
  INV_X1 U619 ( .A(n529), .ZN(n698) );
  INV_X1 U620 ( .A(n530), .ZN(n557) );
  INV_X1 U621 ( .A(n565), .ZN(n532) );
  XNOR2_X1 U622 ( .A(n535), .B(KEYINPUT46), .ZN(n578) );
  INV_X1 U623 ( .A(KEYINPUT19), .ZN(n536) );
  INV_X1 U624 ( .A(n549), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n538), .A2(KEYINPUT82), .ZN(n544) );
  AND2_X1 U626 ( .A1(n531), .A2(n557), .ZN(n747) );
  INV_X1 U627 ( .A(n747), .ZN(n539) );
  AND2_X1 U628 ( .A1(n539), .A2(n565), .ZN(n702) );
  NOR2_X1 U629 ( .A1(n702), .A2(KEYINPUT77), .ZN(n542) );
  INV_X1 U630 ( .A(KEYINPUT47), .ZN(n541) );
  INV_X1 U631 ( .A(KEYINPUT82), .ZN(n540) );
  NAND2_X1 U632 ( .A1(n541), .A2(n540), .ZN(n545) );
  AND2_X1 U633 ( .A1(n542), .A2(n545), .ZN(n543) );
  NAND2_X1 U634 ( .A1(n544), .A2(n543), .ZN(n548) );
  INV_X1 U635 ( .A(n545), .ZN(n546) );
  OR2_X1 U636 ( .A1(n546), .A2(KEYINPUT47), .ZN(n547) );
  NAND2_X1 U637 ( .A1(n548), .A2(n547), .ZN(n554) );
  INV_X1 U638 ( .A(n702), .ZN(n623) );
  NOR2_X1 U639 ( .A1(KEYINPUT77), .A2(KEYINPUT47), .ZN(n550) );
  NAND2_X1 U640 ( .A1(n623), .A2(n550), .ZN(n551) );
  NAND2_X1 U641 ( .A1(n551), .A2(KEYINPUT82), .ZN(n552) );
  NAND2_X1 U642 ( .A1(n549), .A2(n552), .ZN(n553) );
  NAND2_X1 U643 ( .A1(n554), .A2(n553), .ZN(n564) );
  NAND2_X1 U644 ( .A1(n549), .A2(n623), .ZN(n555) );
  NAND2_X1 U645 ( .A1(n555), .A2(KEYINPUT77), .ZN(n563) );
  INV_X1 U646 ( .A(n531), .ZN(n558) );
  NAND2_X1 U647 ( .A1(n558), .A2(n557), .ZN(n560) );
  INV_X1 U648 ( .A(KEYINPUT106), .ZN(n559) );
  XNOR2_X1 U649 ( .A(n560), .B(n559), .ZN(n598) );
  AND2_X1 U650 ( .A1(n580), .A2(n598), .ZN(n562) );
  NAND2_X1 U651 ( .A1(n562), .A2(n561), .ZN(n741) );
  XNOR2_X1 U652 ( .A(n619), .B(KEYINPUT6), .ZN(n625) );
  NAND2_X1 U653 ( .A1(n356), .A2(n580), .ZN(n570) );
  INV_X1 U654 ( .A(KEYINPUT36), .ZN(n569) );
  XNOR2_X1 U655 ( .A(n570), .B(n569), .ZN(n574) );
  XNOR2_X1 U656 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n571) );
  XNOR2_X1 U657 ( .A(n572), .B(n571), .ZN(n686) );
  INV_X1 U658 ( .A(n686), .ZN(n573) );
  XNOR2_X1 U659 ( .A(n573), .B(KEYINPUT88), .ZN(n605) );
  XNOR2_X1 U660 ( .A(n646), .B(KEYINPUT85), .ZN(n575) );
  NAND2_X1 U661 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U662 ( .A1(n356), .A2(n686), .ZN(n579) );
  XNOR2_X1 U663 ( .A(n579), .B(KEYINPUT43), .ZN(n582) );
  INV_X1 U664 ( .A(n580), .ZN(n581) );
  NAND2_X1 U665 ( .A1(n582), .A2(n581), .ZN(n644) );
  NAND2_X1 U666 ( .A1(n583), .A2(n747), .ZN(n643) );
  NOR2_X1 U667 ( .A1(n585), .A2(G898), .ZN(n586) );
  NOR2_X1 U668 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X2 U669 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U670 ( .A(n685), .ZN(n616) );
  NAND2_X1 U671 ( .A1(n625), .A2(n616), .ZN(n592) );
  OR2_X1 U672 ( .A1(n686), .A2(n592), .ZN(n594) );
  INV_X1 U673 ( .A(KEYINPUT33), .ZN(n593) );
  XNOR2_X1 U674 ( .A(n594), .B(n593), .ZN(n712) );
  INV_X1 U675 ( .A(n712), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n622), .A2(n595), .ZN(n597) );
  INV_X1 U677 ( .A(KEYINPUT34), .ZN(n596) );
  XNOR2_X1 U678 ( .A(n597), .B(n596), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n600) );
  INV_X1 U680 ( .A(KEYINPUT22), .ZN(n602) );
  INV_X1 U681 ( .A(n625), .ZN(n604) );
  AND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U683 ( .A(KEYINPUT67), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT32), .ZN(n608) );
  INV_X1 U685 ( .A(KEYINPUT44), .ZN(n612) );
  NOR2_X1 U686 ( .A1(n736), .A2(n612), .ZN(n610) );
  AND2_X1 U687 ( .A1(n648), .A2(n610), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(KEYINPUT86), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n736), .A2(KEYINPUT44), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n648), .A2(n614), .ZN(n615) );
  INV_X1 U691 ( .A(n619), .ZN(n690) );
  NAND2_X1 U692 ( .A1(n616), .A2(n690), .ZN(n617) );
  OR2_X1 U693 ( .A1(n686), .A2(n617), .ZN(n693) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT31), .ZN(n748) );
  AND2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n732) );
  OR2_X1 U697 ( .A1(n748), .A2(n732), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n630) );
  NOR2_X1 U699 ( .A1(n625), .A2(n681), .ZN(n626) );
  AND2_X1 U700 ( .A1(n686), .A2(n626), .ZN(n627) );
  AND2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n729) );
  INV_X1 U702 ( .A(n729), .ZN(n629) );
  AND2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n631) );
  INV_X1 U704 ( .A(KEYINPUT79), .ZN(n720) );
  INV_X1 U705 ( .A(KEYINPUT2), .ZN(n718) );
  NAND2_X1 U706 ( .A1(n718), .A2(KEYINPUT79), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n671), .A2(G478), .ZN(n637) );
  XNOR2_X1 U708 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n635) );
  INV_X1 U709 ( .A(G952), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n638), .A2(G953), .ZN(n639) );
  NAND2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n642), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X1 U713 ( .A(n643), .B(G134), .ZN(G36) );
  XNOR2_X1 U714 ( .A(n644), .B(G140), .ZN(G42) );
  XNOR2_X1 U715 ( .A(G125), .B(KEYINPUT37), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(G27) );
  XOR2_X1 U717 ( .A(G131), .B(n647), .Z(G33) );
  XNOR2_X1 U718 ( .A(n648), .B(G119), .ZN(G21) );
  NAND2_X1 U719 ( .A1(n671), .A2(G472), .ZN(n651) );
  XOR2_X1 U720 ( .A(KEYINPUT62), .B(n649), .Z(n650) );
  XNOR2_X1 U721 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X2 U722 ( .A1(n652), .A2(n677), .ZN(n654) );
  XNOR2_X1 U723 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n654), .B(n653), .ZN(G57) );
  BUF_X1 U725 ( .A(n671), .Z(n665) );
  NAND2_X1 U726 ( .A1(n665), .A2(G217), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT124), .B(n655), .Z(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n658), .A2(n677), .ZN(G66) );
  NAND2_X1 U730 ( .A1(n671), .A2(G475), .ZN(n662) );
  XNOR2_X1 U731 ( .A(KEYINPUT69), .B(KEYINPUT59), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X2 U734 ( .A1(n663), .A2(n677), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n664), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U736 ( .A1(n665), .A2(G469), .ZN(n669) );
  XOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n666) );
  XNOR2_X1 U738 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U739 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U740 ( .A1(n670), .A2(n677), .ZN(G54) );
  NAND2_X1 U741 ( .A1(n671), .A2(G210), .ZN(n676) );
  XOR2_X1 U742 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n673) );
  XNOR2_X1 U743 ( .A(n673), .B(KEYINPUT55), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n672), .B(n674), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n676), .B(n675), .ZN(n678) );
  NOR2_X2 U746 ( .A1(n678), .A2(n677), .ZN(n680) );
  XNOR2_X1 U747 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n680), .B(n679), .ZN(G51) );
  XOR2_X1 U749 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n684) );
  NAND2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(n684), .B(n683), .ZN(n692) );
  NAND2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U753 ( .A(n687), .B(KEYINPUT117), .ZN(n688) );
  XNOR2_X1 U754 ( .A(KEYINPUT50), .B(n688), .ZN(n689) );
  NOR2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U758 ( .A(KEYINPUT51), .B(n695), .ZN(n696) );
  NOR2_X1 U759 ( .A1(n696), .A2(n713), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n704) );
  NOR2_X1 U762 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U764 ( .A1(n705), .A2(n712), .ZN(n706) );
  NOR2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U766 ( .A(n708), .B(KEYINPUT52), .ZN(n710) );
  NOR2_X1 U767 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n711), .B(KEYINPUT118), .ZN(n716) );
  OR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U770 ( .A1(n714), .A2(n772), .ZN(n715) );
  NOR2_X1 U771 ( .A1(n716), .A2(n715), .ZN(n726) );
  NOR2_X1 U772 ( .A1(n717), .A2(KEYINPUT81), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n719), .B(n718), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U775 ( .A1(n717), .A2(KEYINPUT2), .ZN(n722) );
  NAND2_X1 U776 ( .A1(n722), .A2(KEYINPUT79), .ZN(n723) );
  NAND2_X1 U777 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U779 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n728), .B(n727), .ZN(G75) );
  XOR2_X1 U781 ( .A(G101), .B(n729), .Z(G3) );
  XOR2_X1 U782 ( .A(G104), .B(KEYINPUT111), .Z(n731) );
  NAND2_X1 U783 ( .A1(n732), .A2(n745), .ZN(n730) );
  XNOR2_X1 U784 ( .A(n731), .B(n730), .ZN(G6) );
  XOR2_X1 U785 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n734) );
  NAND2_X1 U786 ( .A1(n732), .A2(n747), .ZN(n733) );
  XNOR2_X1 U787 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U788 ( .A(G107), .B(n735), .ZN(G9) );
  XOR2_X1 U789 ( .A(G110), .B(n736), .Z(n737) );
  XNOR2_X1 U790 ( .A(KEYINPUT112), .B(n737), .ZN(G12) );
  XOR2_X1 U791 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n739) );
  NAND2_X1 U792 ( .A1(n549), .A2(n747), .ZN(n738) );
  XNOR2_X1 U793 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U794 ( .A(G128), .B(n740), .Z(G30) );
  XNOR2_X1 U795 ( .A(n741), .B(G143), .ZN(n742) );
  XNOR2_X1 U796 ( .A(KEYINPUT114), .B(n742), .ZN(G45) );
  XOR2_X1 U797 ( .A(G146), .B(KEYINPUT115), .Z(n744) );
  NAND2_X1 U798 ( .A1(n549), .A2(n745), .ZN(n743) );
  XNOR2_X1 U799 ( .A(n744), .B(n743), .ZN(G48) );
  NAND2_X1 U800 ( .A1(n748), .A2(n745), .ZN(n746) );
  XNOR2_X1 U801 ( .A(n746), .B(G113), .ZN(G15) );
  NAND2_X1 U802 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U803 ( .A(n749), .B(G116), .ZN(G18) );
  NOR2_X1 U804 ( .A1(n750), .A2(G953), .ZN(n756) );
  NAND2_X1 U805 ( .A1(G224), .A2(KEYINPUT61), .ZN(n751) );
  NAND2_X1 U806 ( .A1(G898), .A2(n751), .ZN(n754) );
  AND2_X1 U807 ( .A1(G953), .A2(G224), .ZN(n752) );
  NOR2_X1 U808 ( .A1(KEYINPUT61), .A2(n752), .ZN(n753) );
  NOR2_X1 U809 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n763) );
  XNOR2_X1 U811 ( .A(G101), .B(n757), .ZN(n759) );
  XNOR2_X1 U812 ( .A(n759), .B(n758), .ZN(n761) );
  NOR2_X1 U813 ( .A1(G898), .A2(n772), .ZN(n760) );
  NOR2_X1 U814 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U815 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U816 ( .A(KEYINPUT125), .B(n764), .ZN(G69) );
  XOR2_X1 U817 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n768) );
  XNOR2_X1 U818 ( .A(n766), .B(n765), .ZN(n767) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(n769) );
  XNOR2_X1 U820 ( .A(n770), .B(n769), .ZN(n774) );
  XNOR2_X1 U821 ( .A(n771), .B(n774), .ZN(n773) );
  NAND2_X1 U822 ( .A1(n773), .A2(n772), .ZN(n778) );
  XOR2_X1 U823 ( .A(G227), .B(n774), .Z(n775) );
  NAND2_X1 U824 ( .A1(n775), .A2(G900), .ZN(n776) );
  NAND2_X1 U825 ( .A1(n776), .A2(G953), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n778), .A2(n777), .ZN(G72) );
  XOR2_X1 U827 ( .A(G137), .B(n779), .Z(G39) );
endmodule

