

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769;

  XNOR2_X1 U369 ( .A(n390), .B(n357), .ZN(n597) );
  OR2_X1 U370 ( .A1(n650), .A2(G902), .ZN(n472) );
  XNOR2_X1 U371 ( .A(n411), .B(G113), .ZN(n486) );
  XNOR2_X2 U372 ( .A(n571), .B(n570), .ZN(n719) );
  NOR2_X1 U373 ( .A1(G953), .A2(G237), .ZN(n391) );
  NOR2_X1 U374 ( .A1(n542), .A2(n541), .ZN(n543) );
  AND2_X1 U375 ( .A1(n399), .A2(n543), .ZN(n404) );
  XNOR2_X1 U376 ( .A(n490), .B(n489), .ZN(n744) );
  INV_X2 U377 ( .A(G953), .ZN(n759) );
  INV_X1 U378 ( .A(n545), .ZN(n347) );
  XNOR2_X1 U379 ( .A(n554), .B(KEYINPUT42), .ZN(n768) );
  AND2_X1 U380 ( .A1(n556), .A2(n543), .ZN(n402) );
  BUF_X2 U381 ( .A(n663), .Z(n671) );
  XNOR2_X2 U382 ( .A(G104), .B(G122), .ZN(n411) );
  NOR2_X1 U383 ( .A1(n523), .A2(n550), .ZN(n429) );
  INV_X1 U384 ( .A(n696), .ZN(n530) );
  NOR2_X2 U385 ( .A1(n769), .A2(n768), .ZN(n555) );
  BUF_X1 U386 ( .A(n597), .Z(n587) );
  XNOR2_X1 U387 ( .A(n347), .B(n546), .ZN(n721) );
  INV_X1 U388 ( .A(n693), .ZN(n560) );
  OR2_X1 U389 ( .A1(n641), .A2(n492), .ZN(n498) );
  XNOR2_X1 U390 ( .A(n514), .B(KEYINPUT113), .ZN(n766) );
  AND2_X1 U391 ( .A1(n533), .A2(n360), .ZN(n540) );
  NOR2_X1 U392 ( .A1(n715), .A2(n583), .ZN(n585) );
  XNOR2_X1 U393 ( .A(n473), .B(KEYINPUT111), .ZN(n559) );
  BUF_X1 U394 ( .A(n523), .Z(n524) );
  OR2_X1 U395 ( .A1(n657), .A2(G902), .ZN(n459) );
  XNOR2_X1 U396 ( .A(n391), .B(KEYINPUT78), .ZN(n466) );
  XNOR2_X1 U397 ( .A(G146), .B(G125), .ZN(n478) );
  XNOR2_X1 U398 ( .A(KEYINPUT100), .B(KEYINPUT23), .ZN(n444) );
  XNOR2_X1 U399 ( .A(KEYINPUT24), .B(KEYINPUT98), .ZN(n445) );
  XNOR2_X1 U400 ( .A(G128), .B(G110), .ZN(n443) );
  XNOR2_X1 U401 ( .A(G119), .B(KEYINPUT99), .ZN(n442) );
  XNOR2_X1 U402 ( .A(n510), .B(n509), .ZN(n674) );
  NOR2_X1 U403 ( .A1(n589), .A2(n709), .ZN(n681) );
  XNOR2_X2 U404 ( .A(n476), .B(n463), .ZN(n757) );
  AND2_X1 U405 ( .A1(n532), .A2(n645), .ZN(n360) );
  XNOR2_X1 U406 ( .A(KEYINPUT46), .B(n555), .ZN(n556) );
  AND2_X1 U407 ( .A1(n351), .A2(n558), .ZN(n400) );
  AND2_X1 U408 ( .A1(n351), .A2(n405), .ZN(n399) );
  NAND2_X1 U409 ( .A1(n363), .A2(n362), .ZN(n361) );
  INV_X1 U410 ( .A(n681), .ZN(n362) );
  NOR2_X1 U411 ( .A1(n624), .A2(KEYINPUT65), .ZN(n618) );
  INV_X1 U412 ( .A(G237), .ZN(n493) );
  OR2_X2 U413 ( .A1(n381), .A2(n378), .ZN(n536) );
  NAND2_X1 U414 ( .A1(n383), .A2(n382), .ZN(n381) );
  XNOR2_X1 U415 ( .A(n364), .B(KEYINPUT39), .ZN(n566) );
  NAND2_X1 U416 ( .A1(n693), .A2(n356), .ZN(n396) );
  NOR2_X1 U417 ( .A1(n375), .A2(n353), .ZN(n373) );
  NAND2_X1 U418 ( .A1(n719), .A2(n376), .ZN(n374) );
  NAND2_X1 U419 ( .A1(n663), .A2(G210), .ZN(n370) );
  INV_X1 U420 ( .A(n358), .ZN(n377) );
  NAND2_X1 U421 ( .A1(n380), .A2(n494), .ZN(n379) );
  NAND2_X1 U422 ( .A1(n674), .A2(n512), .ZN(n383) );
  XNOR2_X1 U423 ( .A(G137), .B(KEYINPUT5), .ZN(n464) );
  XOR2_X1 U424 ( .A(G113), .B(G116), .Z(n465) );
  NAND2_X1 U425 ( .A1(n404), .A2(n350), .ZN(n403) );
  NOR2_X1 U426 ( .A1(n603), .A2(n679), .ZN(n604) );
  XNOR2_X1 U427 ( .A(KEYINPUT3), .B(G119), .ZN(n485) );
  XNOR2_X1 U428 ( .A(KEYINPUT95), .B(KEYINPUT17), .ZN(n480) );
  XNOR2_X1 U429 ( .A(KEYINPUT18), .B(KEYINPUT93), .ZN(n477) );
  NAND2_X1 U430 ( .A1(G234), .A2(G237), .ZN(n430) );
  AND2_X1 U431 ( .A1(n587), .A2(n377), .ZN(n376) );
  NOR2_X1 U432 ( .A1(n587), .A2(n377), .ZN(n375) );
  NOR2_X1 U433 ( .A1(n500), .A2(KEYINPUT19), .ZN(n388) );
  XNOR2_X1 U434 ( .A(G107), .B(G116), .ZN(n488) );
  XNOR2_X1 U435 ( .A(G134), .B(G122), .ZN(n422) );
  XNOR2_X1 U436 ( .A(G107), .B(G104), .ZN(n502) );
  XNOR2_X1 U437 ( .A(n534), .B(n366), .ZN(n365) );
  INV_X1 U438 ( .A(KEYINPUT30), .ZN(n366) );
  AND2_X1 U439 ( .A1(n703), .A2(n536), .ZN(n586) );
  NAND2_X1 U440 ( .A1(n513), .A2(n567), .ZN(n514) );
  NAND2_X1 U441 ( .A1(n393), .A2(n392), .ZN(n513) );
  NAND2_X1 U442 ( .A1(n398), .A2(n501), .ZN(n392) );
  NAND2_X1 U443 ( .A1(n352), .A2(n371), .ZN(n580) );
  INV_X1 U444 ( .A(KEYINPUT56), .ZN(n367) );
  NAND2_X1 U445 ( .A1(n369), .A2(n667), .ZN(n368) );
  XNOR2_X1 U446 ( .A(n370), .B(n642), .ZN(n369) );
  AND2_X1 U447 ( .A1(n347), .A2(n720), .ZN(n348) );
  AND2_X1 U448 ( .A1(n365), .A2(n586), .ZN(n349) );
  AND2_X1 U449 ( .A1(n544), .A2(n556), .ZN(n350) );
  AND2_X1 U450 ( .A1(n646), .A2(n700), .ZN(n351) );
  AND2_X1 U451 ( .A1(n374), .A2(n373), .ZN(n352) );
  OR2_X1 U452 ( .A1(n524), .A2(n578), .ZN(n353) );
  XOR2_X1 U453 ( .A(n521), .B(n520), .Z(n354) );
  AND2_X1 U454 ( .A1(n632), .A2(KEYINPUT2), .ZN(n355) );
  AND2_X1 U455 ( .A1(n348), .A2(KEYINPUT36), .ZN(n356) );
  XOR2_X1 U456 ( .A(n577), .B(KEYINPUT0), .Z(n357) );
  XOR2_X1 U457 ( .A(KEYINPUT81), .B(KEYINPUT34), .Z(n358) );
  NAND2_X1 U458 ( .A1(n359), .A2(n403), .ZN(n632) );
  NAND2_X1 U459 ( .A1(n401), .A2(n400), .ZN(n359) );
  NAND2_X1 U460 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U461 ( .A1(n361), .A2(n590), .ZN(n384) );
  INV_X1 U462 ( .A(n695), .ZN(n363) );
  NAND2_X1 U463 ( .A1(n548), .A2(n349), .ZN(n364) );
  XNOR2_X1 U464 ( .A(n368), .B(n367), .ZN(G51) );
  NAND2_X1 U465 ( .A1(n372), .A2(n358), .ZN(n371) );
  INV_X1 U466 ( .A(n719), .ZN(n372) );
  NOR2_X1 U467 ( .A1(n674), .A2(n379), .ZN(n378) );
  INV_X1 U468 ( .A(n512), .ZN(n380) );
  NAND2_X1 U469 ( .A1(n512), .A2(G902), .ZN(n382) );
  INV_X1 U470 ( .A(n567), .ZN(n705) );
  XNOR2_X2 U471 ( .A(n536), .B(KEYINPUT1), .ZN(n567) );
  NOR2_X2 U472 ( .A1(n581), .A2(n519), .ZN(n521) );
  AND2_X2 U473 ( .A1(n605), .A2(n604), .ZN(n628) );
  NAND2_X1 U474 ( .A1(n649), .A2(n606), .ZN(n619) );
  OR2_X2 U475 ( .A1(n649), .A2(n606), .ZN(n605) );
  NAND2_X1 U476 ( .A1(n384), .A2(n594), .ZN(n603) );
  XNOR2_X1 U477 ( .A(n585), .B(n584), .ZN(n695) );
  AND2_X1 U478 ( .A1(n385), .A2(n389), .ZN(n387) );
  NAND2_X1 U479 ( .A1(n545), .A2(KEYINPUT19), .ZN(n385) );
  NAND2_X1 U480 ( .A1(n387), .A2(n386), .ZN(n576) );
  NAND2_X1 U481 ( .A1(n347), .A2(n388), .ZN(n386) );
  NAND2_X1 U482 ( .A1(n500), .A2(KEYINPUT19), .ZN(n389) );
  NAND2_X1 U483 ( .A1(n576), .A2(n575), .ZN(n390) );
  NAND2_X1 U484 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U485 ( .A1(n559), .A2(KEYINPUT36), .ZN(n394) );
  NAND2_X1 U486 ( .A1(n397), .A2(n396), .ZN(n395) );
  INV_X1 U487 ( .A(n559), .ZN(n397) );
  NAND2_X1 U488 ( .A1(n693), .A2(n348), .ZN(n398) );
  NAND2_X1 U489 ( .A1(n544), .A2(n402), .ZN(n401) );
  INV_X1 U490 ( .A(n558), .ZN(n405) );
  XNOR2_X2 U491 ( .A(n535), .B(KEYINPUT69), .ZN(n703) );
  XNOR2_X1 U492 ( .A(n709), .B(KEYINPUT6), .ZN(n611) );
  XNOR2_X2 U493 ( .A(KEYINPUT68), .B(G101), .ZN(n475) );
  INV_X1 U494 ( .A(KEYINPUT48), .ZN(n557) );
  INV_X1 U495 ( .A(KEYINPUT79), .ZN(n630) );
  XNOR2_X1 U496 ( .A(n557), .B(KEYINPUT72), .ZN(n558) );
  XNOR2_X1 U497 ( .A(n503), .B(n502), .ZN(n506) );
  INV_X1 U498 ( .A(KEYINPUT28), .ZN(n520) );
  XNOR2_X1 U499 ( .A(n486), .B(n412), .ZN(n413) );
  INV_X1 U500 ( .A(KEYINPUT36), .ZN(n501) );
  XNOR2_X1 U501 ( .A(n414), .B(n413), .ZN(n664) );
  XNOR2_X1 U502 ( .A(KEYINPUT105), .B(KEYINPUT31), .ZN(n584) );
  OR2_X2 U503 ( .A1(n553), .A2(n522), .ZN(n528) );
  BUF_X1 U504 ( .A(n545), .Z(n564) );
  XOR2_X1 U505 ( .A(KEYINPUT12), .B(G140), .Z(n407) );
  XNOR2_X1 U506 ( .A(G143), .B(G131), .ZN(n406) );
  XNOR2_X1 U507 ( .A(n407), .B(n406), .ZN(n410) );
  XNOR2_X1 U508 ( .A(n478), .B(KEYINPUT10), .ZN(n452) );
  XNOR2_X1 U509 ( .A(KEYINPUT106), .B(KEYINPUT11), .ZN(n408) );
  XNOR2_X1 U510 ( .A(n452), .B(n408), .ZN(n409) );
  XOR2_X1 U511 ( .A(n410), .B(n409), .Z(n414) );
  NAND2_X1 U512 ( .A1(G214), .A2(n466), .ZN(n412) );
  INV_X1 U513 ( .A(G902), .ZN(n494) );
  NAND2_X1 U514 ( .A1(n664), .A2(n494), .ZN(n418) );
  XNOR2_X1 U515 ( .A(KEYINPUT107), .B(KEYINPUT13), .ZN(n416) );
  INV_X1 U516 ( .A(G475), .ZN(n415) );
  XNOR2_X1 U517 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U518 ( .A(n418), .B(n417), .ZN(n523) );
  XNOR2_X1 U519 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n420) );
  NAND2_X1 U520 ( .A1(n759), .A2(G234), .ZN(n419) );
  XNOR2_X1 U521 ( .A(n420), .B(n419), .ZN(n448) );
  AND2_X1 U522 ( .A1(n448), .A2(G217), .ZN(n427) );
  XNOR2_X1 U523 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n421) );
  XNOR2_X1 U524 ( .A(n421), .B(n488), .ZN(n425) );
  XNOR2_X2 U525 ( .A(G143), .B(G128), .ZN(n461) );
  XNOR2_X1 U526 ( .A(KEYINPUT108), .B(n422), .ZN(n423) );
  XNOR2_X1 U527 ( .A(n461), .B(n423), .ZN(n424) );
  XNOR2_X1 U528 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U529 ( .A(n427), .B(n426), .ZN(n659) );
  NAND2_X1 U530 ( .A1(n659), .A2(n494), .ZN(n428) );
  XNOR2_X1 U531 ( .A(n428), .B(G478), .ZN(n550) );
  XOR2_X2 U532 ( .A(n429), .B(KEYINPUT109), .Z(n693) );
  XNOR2_X1 U533 ( .A(n430), .B(KEYINPUT96), .ZN(n431) );
  XNOR2_X1 U534 ( .A(KEYINPUT14), .B(n431), .ZN(n434) );
  NAND2_X1 U535 ( .A1(n434), .A2(G952), .ZN(n432) );
  XOR2_X1 U536 ( .A(KEYINPUT97), .B(n432), .Z(n733) );
  INV_X1 U537 ( .A(n733), .ZN(n433) );
  NAND2_X1 U538 ( .A1(n433), .A2(n759), .ZN(n574) );
  AND2_X1 U539 ( .A1(n434), .A2(G953), .ZN(n435) );
  NAND2_X1 U540 ( .A1(G902), .A2(n435), .ZN(n572) );
  OR2_X1 U541 ( .A1(G900), .A2(n572), .ZN(n436) );
  NAND2_X1 U542 ( .A1(n574), .A2(n436), .ZN(n547) );
  INV_X1 U543 ( .A(n547), .ZN(n441) );
  XNOR2_X1 U544 ( .A(G902), .B(KEYINPUT15), .ZN(n637) );
  NAND2_X1 U545 ( .A1(n637), .A2(G234), .ZN(n438) );
  XNOR2_X1 U546 ( .A(KEYINPUT20), .B(KEYINPUT102), .ZN(n437) );
  XNOR2_X1 U547 ( .A(n438), .B(n437), .ZN(n454) );
  NAND2_X1 U548 ( .A1(n454), .A2(G221), .ZN(n440) );
  XNOR2_X1 U549 ( .A(KEYINPUT103), .B(KEYINPUT21), .ZN(n439) );
  XNOR2_X1 U550 ( .A(n440), .B(n439), .ZN(n710) );
  INV_X1 U551 ( .A(n710), .ZN(n595) );
  NOR2_X1 U552 ( .A1(n441), .A2(n595), .ZN(n460) );
  XNOR2_X1 U553 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U554 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U555 ( .A(n447), .B(n446), .ZN(n450) );
  NAND2_X1 U556 ( .A1(n448), .A2(G221), .ZN(n449) );
  XNOR2_X1 U557 ( .A(n450), .B(n449), .ZN(n453) );
  INV_X1 U558 ( .A(G140), .ZN(n451) );
  XNOR2_X1 U559 ( .A(n451), .B(G137), .ZN(n504) );
  XNOR2_X1 U560 ( .A(n452), .B(n504), .ZN(n758) );
  XNOR2_X1 U561 ( .A(n453), .B(n758), .ZN(n657) );
  NAND2_X1 U562 ( .A1(n454), .A2(G217), .ZN(n457) );
  XNOR2_X1 U563 ( .A(KEYINPUT80), .B(KEYINPUT101), .ZN(n455) );
  XNOR2_X1 U564 ( .A(n455), .B(KEYINPUT25), .ZN(n456) );
  XNOR2_X1 U565 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X2 U566 ( .A(n459), .B(n458), .ZN(n600) );
  INV_X1 U567 ( .A(n600), .ZN(n612) );
  NAND2_X1 U568 ( .A1(n460), .A2(n612), .ZN(n519) );
  XNOR2_X2 U569 ( .A(n461), .B(KEYINPUT4), .ZN(n476) );
  INV_X1 U570 ( .A(G134), .ZN(n462) );
  XNOR2_X1 U571 ( .A(n462), .B(G131), .ZN(n463) );
  XNOR2_X2 U572 ( .A(n757), .B(G146), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n465), .B(n464), .ZN(n468) );
  NAND2_X1 U574 ( .A1(G210), .A2(n466), .ZN(n467) );
  XNOR2_X1 U575 ( .A(n468), .B(n467), .ZN(n470) );
  XNOR2_X1 U576 ( .A(n485), .B(n475), .ZN(n469) );
  XNOR2_X1 U577 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U578 ( .A(n510), .B(n471), .ZN(n650) );
  XNOR2_X2 U579 ( .A(n472), .B(G472), .ZN(n709) );
  NOR2_X1 U580 ( .A1(n519), .A2(n611), .ZN(n473) );
  XNOR2_X1 U581 ( .A(KEYINPUT74), .B(G110), .ZN(n474) );
  XNOR2_X1 U582 ( .A(n475), .B(n474), .ZN(n507) );
  XNOR2_X1 U583 ( .A(n507), .B(n476), .ZN(n484) );
  XNOR2_X1 U584 ( .A(n478), .B(n477), .ZN(n482) );
  NAND2_X1 U585 ( .A1(n759), .A2(G224), .ZN(n479) );
  XNOR2_X1 U586 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U587 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U588 ( .A(n484), .B(n483), .ZN(n491) );
  XNOR2_X1 U589 ( .A(n486), .B(n485), .ZN(n490) );
  XNOR2_X1 U590 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n487) );
  XNOR2_X1 U591 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U592 ( .A(n491), .B(n744), .ZN(n641) );
  INV_X1 U593 ( .A(n637), .ZN(n492) );
  NAND2_X1 U594 ( .A1(n494), .A2(n493), .ZN(n499) );
  NAND2_X1 U595 ( .A1(n499), .A2(G210), .ZN(n496) );
  INV_X1 U596 ( .A(KEYINPUT83), .ZN(n495) );
  XNOR2_X1 U597 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X2 U598 ( .A(n498), .B(n497), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n499), .A2(G214), .ZN(n720) );
  INV_X1 U600 ( .A(n720), .ZN(n500) );
  NAND2_X1 U601 ( .A1(G227), .A2(n759), .ZN(n503) );
  INV_X1 U602 ( .A(n504), .ZN(n505) );
  XNOR2_X1 U603 ( .A(n506), .B(n505), .ZN(n508) );
  XNOR2_X1 U604 ( .A(n508), .B(n507), .ZN(n509) );
  INV_X1 U605 ( .A(KEYINPUT73), .ZN(n511) );
  XNOR2_X1 U606 ( .A(n511), .B(G469), .ZN(n512) );
  INV_X1 U607 ( .A(n766), .ZN(n516) );
  INV_X1 U608 ( .A(KEYINPUT89), .ZN(n515) );
  NAND2_X1 U609 ( .A1(n516), .A2(n515), .ZN(n518) );
  NAND2_X1 U610 ( .A1(n766), .A2(KEYINPUT89), .ZN(n517) );
  NAND2_X1 U611 ( .A1(n518), .A2(n517), .ZN(n544) );
  INV_X1 U612 ( .A(n709), .ZN(n581) );
  NAND2_X1 U613 ( .A1(n354), .A2(n536), .ZN(n553) );
  INV_X1 U614 ( .A(n576), .ZN(n522) );
  INV_X1 U615 ( .A(n528), .ZN(n690) );
  NAND2_X1 U616 ( .A1(n524), .A2(n550), .ZN(n525) );
  XOR2_X1 U617 ( .A(n525), .B(KEYINPUT110), .Z(n696) );
  NAND2_X1 U618 ( .A1(n530), .A2(n560), .ZN(n590) );
  NAND2_X1 U619 ( .A1(n690), .A2(n590), .ZN(n527) );
  XNOR2_X1 U620 ( .A(KEYINPUT47), .B(KEYINPUT70), .ZN(n526) );
  NOR2_X1 U621 ( .A1(n527), .A2(n526), .ZN(n542) );
  NAND2_X1 U622 ( .A1(n528), .A2(KEYINPUT47), .ZN(n529) );
  XNOR2_X1 U623 ( .A(n529), .B(KEYINPUT86), .ZN(n533) );
  AND2_X1 U624 ( .A1(KEYINPUT47), .A2(n560), .ZN(n531) );
  NAND2_X1 U625 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U626 ( .A1(n709), .A2(n720), .ZN(n534) );
  NAND2_X1 U627 ( .A1(n600), .A2(n710), .ZN(n535) );
  NAND2_X1 U628 ( .A1(n547), .A2(n550), .ZN(n537) );
  OR2_X1 U629 ( .A1(n524), .A2(n537), .ZN(n538) );
  NOR2_X1 U630 ( .A1(n538), .A2(n564), .ZN(n539) );
  NAND2_X1 U631 ( .A1(n349), .A2(n539), .ZN(n645) );
  XNOR2_X1 U632 ( .A(KEYINPUT85), .B(n540), .ZN(n541) );
  INV_X1 U633 ( .A(KEYINPUT38), .ZN(n546) );
  AND2_X1 U634 ( .A1(n721), .A2(n547), .ZN(n548) );
  AND2_X1 U635 ( .A1(n566), .A2(n693), .ZN(n549) );
  XNOR2_X1 U636 ( .A(KEYINPUT40), .B(n549), .ZN(n769) );
  INV_X1 U637 ( .A(n550), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n524), .A2(n578), .ZN(n723) );
  NAND2_X1 U639 ( .A1(n721), .A2(n720), .ZN(n724) );
  NOR2_X1 U640 ( .A1(n723), .A2(n724), .ZN(n552) );
  XNOR2_X1 U641 ( .A(KEYINPUT41), .B(KEYINPUT112), .ZN(n551) );
  XNOR2_X1 U642 ( .A(n552), .B(n551), .ZN(n734) );
  NOR2_X1 U643 ( .A1(n734), .A2(n553), .ZN(n554) );
  NOR2_X1 U644 ( .A1(n560), .A2(n559), .ZN(n561) );
  AND2_X1 U645 ( .A1(n561), .A2(n720), .ZN(n562) );
  NAND2_X1 U646 ( .A1(n562), .A2(n705), .ZN(n563) );
  XNOR2_X1 U647 ( .A(n563), .B(KEYINPUT43), .ZN(n565) );
  NAND2_X1 U648 ( .A1(n565), .A2(n564), .ZN(n646) );
  NAND2_X1 U649 ( .A1(n566), .A2(n696), .ZN(n700) );
  NAND2_X1 U650 ( .A1(n567), .A2(n703), .ZN(n569) );
  INV_X1 U651 ( .A(KEYINPUT77), .ZN(n568) );
  XNOR2_X1 U652 ( .A(n569), .B(n568), .ZN(n582) );
  OR2_X2 U653 ( .A1(n582), .A2(n611), .ZN(n571) );
  XNOR2_X1 U654 ( .A(KEYINPUT92), .B(KEYINPUT33), .ZN(n570) );
  OR2_X1 U655 ( .A1(n572), .A2(G898), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n574), .A2(n573), .ZN(n575) );
  INV_X1 U657 ( .A(KEYINPUT91), .ZN(n577) );
  INV_X1 U658 ( .A(KEYINPUT35), .ZN(n579) );
  XNOR2_X2 U659 ( .A(n580), .B(n579), .ZN(n649) );
  NOR2_X1 U660 ( .A1(KEYINPUT44), .A2(KEYINPUT75), .ZN(n606) );
  OR2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n715) );
  INV_X1 U662 ( .A(n587), .ZN(n583) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n588), .B(KEYINPUT104), .ZN(n589) );
  INV_X1 U665 ( .A(n590), .ZN(n725) );
  INV_X1 U666 ( .A(KEYINPUT44), .ZN(n591) );
  INV_X1 U667 ( .A(KEYINPUT65), .ZN(n620) );
  NAND2_X1 U668 ( .A1(n591), .A2(n620), .ZN(n593) );
  INV_X1 U669 ( .A(KEYINPUT75), .ZN(n621) );
  NAND2_X1 U670 ( .A1(n621), .A2(KEYINPUT44), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U672 ( .A1(n723), .A2(n595), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n599) );
  INV_X1 U674 ( .A(KEYINPUT22), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n599), .B(n598), .ZN(n607) );
  AND2_X1 U676 ( .A1(n600), .A2(n705), .ZN(n601) );
  AND2_X1 U677 ( .A1(n601), .A2(n611), .ZN(n602) );
  AND2_X1 U678 ( .A1(n607), .A2(n602), .ZN(n679) );
  INV_X1 U679 ( .A(n607), .ZN(n616) );
  OR2_X1 U680 ( .A1(n567), .A2(n709), .ZN(n608) );
  NOR2_X1 U681 ( .A1(n616), .A2(n608), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n609), .B(KEYINPUT66), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n610), .A2(n612), .ZN(n648) );
  XNOR2_X1 U684 ( .A(n611), .B(KEYINPUT82), .ZN(n614) );
  AND2_X1 U685 ( .A1(n567), .A2(n612), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n615) );
  OR2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X2 U688 ( .A(n617), .B(KEYINPUT32), .ZN(n647) );
  NAND2_X1 U689 ( .A1(n648), .A2(n647), .ZN(n624) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(n626) );
  NAND2_X1 U691 ( .A1(n620), .A2(KEYINPUT44), .ZN(n622) );
  AND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X2 U695 ( .A(n629), .B(KEYINPUT45), .ZN(n747) );
  NAND2_X1 U696 ( .A1(n355), .A2(n747), .ZN(n631) );
  XNOR2_X1 U697 ( .A(n631), .B(n630), .ZN(n636) );
  XNOR2_X1 U698 ( .A(n632), .B(KEYINPUT88), .ZN(n756) );
  NAND2_X1 U699 ( .A1(n756), .A2(n747), .ZN(n634) );
  INV_X1 U700 ( .A(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n701) );
  NOR2_X2 U703 ( .A1(n701), .A2(n637), .ZN(n638) );
  XNOR2_X2 U704 ( .A(n638), .B(KEYINPUT64), .ZN(n663) );
  XNOR2_X1 U705 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n639) );
  XNOR2_X1 U706 ( .A(n639), .B(KEYINPUT55), .ZN(n640) );
  XNOR2_X1 U707 ( .A(n641), .B(n640), .ZN(n642) );
  INV_X1 U708 ( .A(G952), .ZN(n643) );
  NAND2_X1 U709 ( .A1(n643), .A2(G953), .ZN(n644) );
  XNOR2_X1 U710 ( .A(n644), .B(KEYINPUT94), .ZN(n667) );
  XNOR2_X1 U711 ( .A(n645), .B(G143), .ZN(G45) );
  XNOR2_X1 U712 ( .A(n646), .B(G140), .ZN(G42) );
  XNOR2_X1 U713 ( .A(n647), .B(G119), .ZN(G21) );
  XNOR2_X1 U714 ( .A(n648), .B(G110), .ZN(G12) );
  XNOR2_X1 U715 ( .A(n649), .B(G122), .ZN(G24) );
  NAND2_X1 U716 ( .A1(n663), .A2(G472), .ZN(n652) );
  XOR2_X1 U717 ( .A(KEYINPUT62), .B(n650), .Z(n651) );
  XNOR2_X1 U718 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U719 ( .A1(n653), .A2(n667), .ZN(n655) );
  XNOR2_X1 U720 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n655), .B(n654), .ZN(G57) );
  NAND2_X1 U722 ( .A1(n671), .A2(G217), .ZN(n656) );
  XNOR2_X1 U723 ( .A(n657), .B(n656), .ZN(n658) );
  INV_X1 U724 ( .A(n667), .ZN(n677) );
  NOR2_X1 U725 ( .A1(n658), .A2(n677), .ZN(G66) );
  NAND2_X1 U726 ( .A1(n671), .A2(G478), .ZN(n661) );
  XOR2_X1 U727 ( .A(KEYINPUT124), .B(n659), .Z(n660) );
  XNOR2_X1 U728 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n662), .A2(n677), .ZN(G63) );
  NAND2_X1 U730 ( .A1(n663), .A2(G475), .ZN(n666) );
  XOR2_X1 U731 ( .A(KEYINPUT59), .B(n664), .Z(n665) );
  XNOR2_X1 U732 ( .A(n666), .B(n665), .ZN(n668) );
  NAND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n670) );
  XNOR2_X1 U734 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n670), .B(n669), .ZN(G60) );
  NAND2_X1 U736 ( .A1(n671), .A2(G469), .ZN(n676) );
  XNOR2_X1 U737 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT58), .ZN(n673) );
  XNOR2_X1 U739 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n676), .B(n675), .ZN(n678) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(G54) );
  XOR2_X1 U742 ( .A(G101), .B(n679), .Z(G3) );
  NAND2_X1 U743 ( .A1(n693), .A2(n681), .ZN(n680) );
  XNOR2_X1 U744 ( .A(G104), .B(n680), .ZN(G6) );
  XNOR2_X1 U745 ( .A(G107), .B(KEYINPUT114), .ZN(n685) );
  XOR2_X1 U746 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n683) );
  NAND2_X1 U747 ( .A1(n681), .A2(n696), .ZN(n682) );
  XNOR2_X1 U748 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n685), .B(n684), .ZN(G9) );
  AND2_X1 U750 ( .A1(n690), .A2(n696), .ZN(n689) );
  XOR2_X1 U751 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n687) );
  XNOR2_X1 U752 ( .A(G128), .B(KEYINPUT116), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n689), .B(n688), .ZN(G30) );
  XOR2_X1 U755 ( .A(G146), .B(KEYINPUT117), .Z(n692) );
  NAND2_X1 U756 ( .A1(n690), .A2(n693), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n692), .B(n691), .ZN(G48) );
  NAND2_X1 U758 ( .A1(n695), .A2(n693), .ZN(n694) );
  XNOR2_X1 U759 ( .A(n694), .B(G113), .ZN(G15) );
  NAND2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U761 ( .A(n697), .B(KEYINPUT118), .ZN(n698) );
  XNOR2_X1 U762 ( .A(G116), .B(n698), .ZN(G18) );
  XOR2_X1 U763 ( .A(G134), .B(KEYINPUT119), .Z(n699) );
  XNOR2_X1 U764 ( .A(n700), .B(n699), .ZN(G36) );
  BUF_X1 U765 ( .A(n701), .Z(n702) );
  XOR2_X1 U766 ( .A(KEYINPUT87), .B(n702), .Z(n739) );
  INV_X1 U767 ( .A(n703), .ZN(n704) );
  NAND2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U769 ( .A(n706), .B(KEYINPUT50), .ZN(n707) );
  XNOR2_X1 U770 ( .A(KEYINPUT121), .B(n707), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n709), .A2(n708), .ZN(n714) );
  NOR2_X1 U772 ( .A1(n600), .A2(n710), .ZN(n712) );
  XNOR2_X1 U773 ( .A(KEYINPUT49), .B(KEYINPUT120), .ZN(n711) );
  XNOR2_X1 U774 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U775 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U776 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U777 ( .A(KEYINPUT51), .B(n717), .ZN(n718) );
  NOR2_X1 U778 ( .A1(n734), .A2(n718), .ZN(n730) );
  NOR2_X1 U779 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U780 ( .A1(n723), .A2(n722), .ZN(n727) );
  NOR2_X1 U781 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U782 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U783 ( .A1(n372), .A2(n728), .ZN(n729) );
  NOR2_X1 U784 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U785 ( .A(n731), .B(KEYINPUT52), .ZN(n732) );
  NOR2_X1 U786 ( .A1(n733), .A2(n732), .ZN(n736) );
  NOR2_X1 U787 ( .A1(n734), .A2(n372), .ZN(n735) );
  NOR2_X1 U788 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U789 ( .A(n737), .B(KEYINPUT122), .ZN(n738) );
  NAND2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U791 ( .A1(n740), .A2(G953), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n741), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U793 ( .A(G101), .B(G110), .ZN(n742) );
  XOR2_X1 U794 ( .A(KEYINPUT127), .B(n742), .Z(n743) );
  XNOR2_X1 U795 ( .A(n744), .B(n743), .ZN(n746) );
  NOR2_X1 U796 ( .A1(G898), .A2(n759), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n746), .A2(n745), .ZN(n755) );
  NAND2_X1 U798 ( .A1(n747), .A2(n759), .ZN(n753) );
  XOR2_X1 U799 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n749) );
  NAND2_X1 U800 ( .A1(G224), .A2(G953), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n749), .B(n748), .ZN(n750) );
  NAND2_X1 U802 ( .A1(G898), .A2(n750), .ZN(n751) );
  XNOR2_X1 U803 ( .A(n751), .B(KEYINPUT126), .ZN(n752) );
  NAND2_X1 U804 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U805 ( .A(n755), .B(n754), .ZN(G69) );
  XNOR2_X1 U806 ( .A(n757), .B(n758), .ZN(n761) );
  XNOR2_X1 U807 ( .A(n756), .B(n761), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n760), .A2(n759), .ZN(n765) );
  XOR2_X1 U809 ( .A(G227), .B(n761), .Z(n762) );
  NAND2_X1 U810 ( .A1(n762), .A2(G900), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n763), .A2(G953), .ZN(n764) );
  NAND2_X1 U812 ( .A1(n765), .A2(n764), .ZN(G72) );
  XNOR2_X1 U813 ( .A(n766), .B(G125), .ZN(n767) );
  XNOR2_X1 U814 ( .A(n767), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U815 ( .A(n768), .B(G137), .Z(G39) );
  XOR2_X1 U816 ( .A(G131), .B(n769), .Z(G33) );
endmodule

