

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745;

  NOR2_X2 U369 ( .A1(n644), .A2(n556), .ZN(n593) );
  INV_X1 U370 ( .A(n552), .ZN(n644) );
  XNOR2_X1 U371 ( .A(n416), .B(G110), .ZN(n407) );
  INV_X1 U372 ( .A(G128), .ZN(n404) );
  INV_X2 U373 ( .A(G953), .ZN(n734) );
  NAND2_X2 U374 ( .A1(n368), .A2(n534), .ZN(n535) );
  XNOR2_X2 U375 ( .A(n456), .B(n724), .ZN(n609) );
  XNOR2_X2 U376 ( .A(n455), .B(n454), .ZN(n724) );
  XNOR2_X2 U377 ( .A(n443), .B(n423), .ZN(n732) );
  AND2_X1 U378 ( .A1(n600), .A2(n599), .ZN(n657) );
  NAND2_X2 U379 ( .A1(n367), .A2(n607), .ZN(n608) );
  XNOR2_X2 U380 ( .A(n381), .B(n525), .ZN(n647) );
  AND2_X1 U381 ( .A1(n613), .A2(n618), .ZN(n614) );
  XNOR2_X1 U382 ( .A(n395), .B(n394), .ZN(n393) );
  XNOR2_X1 U383 ( .A(n372), .B(KEYINPUT88), .ZN(n631) );
  NAND2_X1 U384 ( .A1(n521), .A2(n398), .ZN(n372) );
  XNOR2_X1 U385 ( .A(n390), .B(KEYINPUT71), .ZN(n580) );
  NAND2_X1 U386 ( .A1(n391), .A2(n393), .ZN(n390) );
  AND2_X1 U387 ( .A1(n383), .A2(n664), .ZN(n522) );
  XNOR2_X1 U388 ( .A(n392), .B(n571), .ZN(n391) );
  XNOR2_X1 U389 ( .A(n503), .B(n502), .ZN(n526) );
  XNOR2_X1 U390 ( .A(n400), .B(n431), .ZN(n567) );
  XNOR2_X1 U391 ( .A(n667), .B(KEYINPUT102), .ZN(n570) );
  XNOR2_X1 U392 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U393 ( .A(KEYINPUT69), .B(KEYINPUT16), .ZN(n451) );
  XNOR2_X1 U394 ( .A(G107), .B(G104), .ZN(n406) );
  AND2_X1 U395 ( .A1(n744), .A2(n370), .ZN(n361) );
  XNOR2_X2 U396 ( .A(n557), .B(KEYINPUT19), .ZN(n548) );
  XNOR2_X2 U397 ( .A(n450), .B(n415), .ZN(n443) );
  NAND2_X1 U398 ( .A1(n354), .A2(n664), .ZN(n362) );
  XNOR2_X1 U399 ( .A(n490), .B(n489), .ZN(n530) );
  XNOR2_X1 U400 ( .A(n488), .B(n487), .ZN(n489) );
  NOR2_X1 U401 ( .A1(n713), .A2(G902), .ZN(n400) );
  INV_X1 U402 ( .A(KEYINPUT99), .ZN(n371) );
  XNOR2_X1 U403 ( .A(n596), .B(n579), .ZN(n678) );
  XNOR2_X1 U404 ( .A(G116), .B(G122), .ZN(n491) );
  XOR2_X1 U405 ( .A(KEYINPUT95), .B(KEYINPUT7), .Z(n492) );
  XOR2_X1 U406 ( .A(G140), .B(G122), .Z(n481) );
  XNOR2_X1 U407 ( .A(n364), .B(n363), .ZN(n676) );
  INV_X1 U408 ( .A(KEYINPUT41), .ZN(n363) );
  NOR2_X1 U409 ( .A1(n683), .A2(n680), .ZN(n364) );
  INV_X1 U410 ( .A(KEYINPUT1), .ZN(n382) );
  XNOR2_X1 U411 ( .A(n386), .B(n385), .ZN(n546) );
  INV_X1 U412 ( .A(KEYINPUT22), .ZN(n411) );
  XNOR2_X1 U413 ( .A(n401), .B(n425), .ZN(n713) );
  XNOR2_X1 U414 ( .A(n427), .B(n350), .ZN(n401) );
  XNOR2_X1 U415 ( .A(n413), .B(n423), .ZN(n424) );
  INV_X1 U416 ( .A(G237), .ZN(n457) );
  NAND2_X1 U417 ( .A1(n569), .A2(n568), .ZN(n395) );
  INV_X1 U418 ( .A(KEYINPUT72), .ZN(n394) );
  NAND2_X1 U419 ( .A1(n570), .A2(n677), .ZN(n392) );
  NAND2_X1 U420 ( .A1(n387), .A2(n554), .ZN(n386) );
  AND2_X1 U421 ( .A1(n570), .A2(n565), .ZN(n387) );
  XNOR2_X1 U422 ( .A(n543), .B(KEYINPUT106), .ZN(n385) );
  NOR2_X1 U423 ( .A1(G953), .A2(G237), .ZN(n480) );
  XNOR2_X1 U424 ( .A(G137), .B(G101), .ZN(n437) );
  XOR2_X1 U425 ( .A(KEYINPUT5), .B(G146), .Z(n438) );
  XOR2_X1 U426 ( .A(KEYINPUT68), .B(G119), .Z(n435) );
  BUF_X1 U427 ( .A(n657), .Z(n733) );
  XNOR2_X1 U428 ( .A(n399), .B(G140), .ZN(n423) );
  INV_X1 U429 ( .A(G137), .ZN(n399) );
  XOR2_X1 U430 ( .A(G128), .B(G110), .Z(n413) );
  NAND2_X1 U431 ( .A1(G234), .A2(G237), .ZN(n463) );
  NAND2_X1 U432 ( .A1(n397), .A2(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U433 ( .A1(n580), .A2(n678), .ZN(n581) );
  BUF_X1 U434 ( .A(n572), .Z(n596) );
  XNOR2_X1 U435 ( .A(G134), .B(G107), .ZN(n494) );
  XNOR2_X1 U436 ( .A(G113), .B(G104), .ZN(n484) );
  XNOR2_X1 U437 ( .A(n585), .B(n384), .ZN(n586) );
  INV_X1 U438 ( .A(KEYINPUT42), .ZN(n384) );
  NAND2_X1 U439 ( .A1(n582), .A2(n638), .ZN(n623) );
  INV_X1 U440 ( .A(n558), .ZN(n365) );
  INV_X1 U441 ( .A(KEYINPUT35), .ZN(n505) );
  NOR2_X1 U442 ( .A1(n673), .A2(n524), .ZN(n381) );
  BUF_X1 U443 ( .A(n631), .Z(n634) );
  XNOR2_X1 U444 ( .A(n533), .B(n369), .ZN(n368) );
  INV_X1 U445 ( .A(KEYINPUT78), .ZN(n369) );
  XNOR2_X1 U446 ( .A(n713), .B(n712), .ZN(n714) );
  INV_X1 U447 ( .A(G140), .ZN(n651) );
  XNOR2_X1 U448 ( .A(n586), .B(G137), .ZN(G39) );
  XNOR2_X1 U449 ( .A(n360), .B(G119), .ZN(G21) );
  BUF_X1 U450 ( .A(n379), .Z(n360) );
  NOR2_X1 U451 ( .A1(n567), .A2(n518), .ZN(n349) );
  XOR2_X1 U452 ( .A(n422), .B(n421), .Z(n350) );
  XNOR2_X1 U453 ( .A(G146), .B(G125), .ZN(n445) );
  XOR2_X1 U454 ( .A(KEYINPUT18), .B(KEYINPUT82), .Z(n351) );
  AND2_X1 U455 ( .A1(n511), .A2(n553), .ZN(n352) );
  AND2_X1 U456 ( .A1(n514), .A2(n553), .ZN(n353) );
  AND2_X1 U457 ( .A1(n349), .A2(n396), .ZN(n354) );
  AND2_X1 U458 ( .A1(n515), .A2(n514), .ZN(n355) );
  AND2_X1 U459 ( .A1(n599), .A2(n603), .ZN(n356) );
  XOR2_X1 U460 ( .A(KEYINPUT81), .B(KEYINPUT33), .Z(n357) );
  XOR2_X1 U461 ( .A(n616), .B(n615), .Z(n358) );
  AND2_X1 U462 ( .A1(n402), .A2(n602), .ZN(n359) );
  AND2_X2 U463 ( .A1(n361), .A2(n378), .ZN(n377) );
  NAND2_X1 U464 ( .A1(n376), .A2(n540), .ZN(n375) );
  XNOR2_X2 U465 ( .A(n362), .B(n357), .ZN(n688) );
  AND2_X1 U466 ( .A1(n523), .A2(n688), .ZN(n472) );
  XNOR2_X1 U467 ( .A(n532), .B(n371), .ZN(n370) );
  AND2_X1 U468 ( .A1(n366), .A2(n365), .ZN(n559) );
  XNOR2_X1 U469 ( .A(n593), .B(KEYINPUT108), .ZN(n366) );
  NOR2_X1 U470 ( .A1(n563), .A2(n564), .ZN(n578) );
  NAND2_X1 U471 ( .A1(n606), .A2(n605), .ZN(n367) );
  NAND2_X1 U472 ( .A1(n538), .A2(n537), .ZN(n376) );
  NAND2_X2 U473 ( .A1(n379), .A2(n622), .ZN(n516) );
  XNOR2_X2 U474 ( .A(n581), .B(KEYINPUT39), .ZN(n582) );
  XNOR2_X2 U475 ( .A(n373), .B(G472), .ZN(n667) );
  NAND2_X1 U476 ( .A1(n616), .A2(n501), .ZN(n373) );
  XNOR2_X2 U477 ( .A(n374), .B(KEYINPUT45), .ZN(n718) );
  NAND2_X2 U478 ( .A1(n377), .A2(n375), .ZN(n374) );
  NAND2_X1 U479 ( .A1(n408), .A2(n517), .ZN(n378) );
  XNOR2_X2 U480 ( .A(n512), .B(KEYINPUT32), .ZN(n379) );
  NAND2_X1 U481 ( .A1(n380), .A2(n681), .ZN(n532) );
  NAND2_X1 U482 ( .A1(n631), .A2(n647), .ZN(n380) );
  INV_X1 U483 ( .A(n664), .ZN(n514) );
  XNOR2_X2 U484 ( .A(n544), .B(n382), .ZN(n664) );
  AND2_X1 U485 ( .A1(n349), .A2(n667), .ZN(n383) );
  AND2_X2 U486 ( .A1(n657), .A2(n718), .ZN(n606) );
  NAND2_X1 U487 ( .A1(n718), .A2(n388), .ZN(n389) );
  AND2_X1 U488 ( .A1(n600), .A2(n356), .ZN(n388) );
  NAND2_X1 U489 ( .A1(n389), .A2(n359), .ZN(n607) );
  XNOR2_X2 U490 ( .A(n535), .B(KEYINPUT100), .ZN(n744) );
  INV_X1 U491 ( .A(n553), .ZN(n396) );
  INV_X1 U492 ( .A(n606), .ZN(n397) );
  INV_X1 U493 ( .A(n667), .ZN(n398) );
  NAND2_X1 U494 ( .A1(n603), .A2(KEYINPUT2), .ZN(n402) );
  XNOR2_X2 U495 ( .A(n403), .B(n420), .ZN(n544) );
  OR2_X2 U496 ( .A1(n704), .A2(G902), .ZN(n403) );
  INV_X1 U497 ( .A(n414), .ZN(n497) );
  XNOR2_X2 U498 ( .A(n405), .B(n404), .ZN(n414) );
  XNOR2_X2 U499 ( .A(KEYINPUT64), .B(G143), .ZN(n405) );
  XNOR2_X2 U500 ( .A(n407), .B(n406), .ZN(n453) );
  INV_X1 U501 ( .A(n536), .ZN(n408) );
  XNOR2_X2 U502 ( .A(n516), .B(n409), .ZN(n536) );
  INV_X1 U503 ( .A(KEYINPUT79), .ZN(n409) );
  NAND2_X1 U504 ( .A1(n410), .A2(n352), .ZN(n512) );
  NAND2_X1 U505 ( .A1(n410), .A2(n353), .ZN(n533) );
  NAND2_X1 U506 ( .A1(n410), .A2(n355), .ZN(n622) );
  XNOR2_X2 U507 ( .A(n509), .B(n411), .ZN(n410) );
  XNOR2_X1 U508 ( .A(n617), .B(n358), .ZN(n619) );
  NOR2_X2 U509 ( .A1(n518), .A2(n544), .ZN(n569) );
  NAND2_X2 U510 ( .A1(n572), .A2(n677), .ZN(n557) );
  XOR2_X1 U511 ( .A(n609), .B(n611), .Z(n412) );
  NOR2_X1 U512 ( .A1(n734), .A2(G952), .ZN(n717) );
  INV_X1 U513 ( .A(KEYINPUT46), .ZN(n587) );
  INV_X1 U514 ( .A(KEYINPUT11), .ZN(n475) );
  INV_X1 U515 ( .A(n565), .ZN(n566) );
  XNOR2_X1 U516 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U517 ( .A(n478), .B(n477), .ZN(n479) );
  INV_X1 U518 ( .A(KEYINPUT28), .ZN(n543) );
  INV_X1 U519 ( .A(n717), .ZN(n618) );
  XNOR2_X1 U520 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X2 U521 ( .A(n414), .B(KEYINPUT4), .ZN(n450) );
  XNOR2_X1 U522 ( .A(G134), .B(G131), .ZN(n415) );
  XNOR2_X2 U523 ( .A(G101), .B(KEYINPUT83), .ZN(n416) );
  NAND2_X1 U524 ( .A1(n734), .A2(G227), .ZN(n417) );
  XNOR2_X1 U525 ( .A(n417), .B(G146), .ZN(n418) );
  XNOR2_X1 U526 ( .A(n453), .B(n418), .ZN(n419) );
  XNOR2_X1 U527 ( .A(n732), .B(n419), .ZN(n704) );
  XNOR2_X1 U528 ( .A(KEYINPUT67), .B(G469), .ZN(n420) );
  XOR2_X1 U529 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n422) );
  XNOR2_X1 U530 ( .A(G119), .B(KEYINPUT86), .ZN(n421) );
  XNOR2_X1 U531 ( .A(KEYINPUT10), .B(n445), .ZN(n731) );
  XNOR2_X1 U532 ( .A(n731), .B(n424), .ZN(n425) );
  NAND2_X1 U533 ( .A1(G234), .A2(n734), .ZN(n426) );
  XOR2_X1 U534 ( .A(KEYINPUT8), .B(n426), .Z(n496) );
  NAND2_X1 U535 ( .A1(G221), .A2(n496), .ZN(n427) );
  XOR2_X1 U536 ( .A(KEYINPUT25), .B(KEYINPUT73), .Z(n430) );
  XNOR2_X1 U537 ( .A(KEYINPUT15), .B(G902), .ZN(n601) );
  NAND2_X1 U538 ( .A1(n601), .A2(G234), .ZN(n428) );
  XNOR2_X1 U539 ( .A(n428), .B(KEYINPUT20), .ZN(n432) );
  AND2_X1 U540 ( .A1(G217), .A2(n432), .ZN(n429) );
  XNOR2_X1 U541 ( .A(n430), .B(n429), .ZN(n431) );
  AND2_X1 U542 ( .A1(n432), .A2(G221), .ZN(n433) );
  XNOR2_X1 U543 ( .A(n433), .B(KEYINPUT21), .ZN(n668) );
  INV_X1 U544 ( .A(n668), .ZN(n518) );
  XNOR2_X1 U545 ( .A(G116), .B(G113), .ZN(n434) );
  XNOR2_X1 U546 ( .A(n434), .B(KEYINPUT3), .ZN(n436) );
  XNOR2_X1 U547 ( .A(n436), .B(n435), .ZN(n454) );
  XNOR2_X1 U548 ( .A(n438), .B(n437), .ZN(n440) );
  NAND2_X1 U549 ( .A1(n480), .A2(G210), .ZN(n439) );
  XNOR2_X1 U550 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U551 ( .A(n454), .B(n441), .ZN(n442) );
  XNOR2_X1 U552 ( .A(n443), .B(n442), .ZN(n616) );
  INV_X1 U553 ( .A(G902), .ZN(n501) );
  XNOR2_X1 U554 ( .A(n667), .B(KEYINPUT6), .ZN(n553) );
  XNOR2_X1 U555 ( .A(KEYINPUT74), .B(KEYINPUT17), .ZN(n444) );
  XNOR2_X1 U556 ( .A(n351), .B(n444), .ZN(n446) );
  XNOR2_X1 U557 ( .A(n446), .B(n445), .ZN(n448) );
  NAND2_X1 U558 ( .A1(G224), .A2(n734), .ZN(n447) );
  XNOR2_X1 U559 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U560 ( .A(n450), .B(n449), .ZN(n456) );
  XNOR2_X1 U561 ( .A(n451), .B(G122), .ZN(n452) );
  XNOR2_X2 U562 ( .A(n453), .B(n452), .ZN(n455) );
  NAND2_X1 U563 ( .A1(n609), .A2(n601), .ZN(n461) );
  NAND2_X1 U564 ( .A1(n501), .A2(n457), .ZN(n462) );
  NAND2_X1 U565 ( .A1(n462), .A2(G210), .ZN(n459) );
  XNOR2_X1 U566 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X2 U568 ( .A(n461), .B(n460), .ZN(n572) );
  NAND2_X1 U569 ( .A1(n462), .A2(G214), .ZN(n677) );
  XNOR2_X1 U570 ( .A(n463), .B(KEYINPUT14), .ZN(n663) );
  INV_X1 U571 ( .A(G952), .ZN(n464) );
  NAND2_X1 U572 ( .A1(n734), .A2(n464), .ZN(n466) );
  OR2_X1 U573 ( .A1(n734), .A2(G902), .ZN(n465) );
  AND2_X1 U574 ( .A1(n466), .A2(n465), .ZN(n467) );
  AND2_X1 U575 ( .A1(n663), .A2(n467), .ZN(n542) );
  NAND2_X1 U576 ( .A1(G953), .A2(G898), .ZN(n468) );
  AND2_X1 U577 ( .A1(n542), .A2(n468), .ZN(n469) );
  NAND2_X1 U578 ( .A1(n548), .A2(n469), .ZN(n471) );
  INV_X1 U579 ( .A(KEYINPUT0), .ZN(n470) );
  XNOR2_X2 U580 ( .A(n471), .B(n470), .ZN(n523) );
  XNOR2_X1 U581 ( .A(n472), .B(KEYINPUT34), .ZN(n504) );
  XOR2_X1 U582 ( .A(KEYINPUT92), .B(KEYINPUT12), .Z(n474) );
  XNOR2_X1 U583 ( .A(KEYINPUT91), .B(KEYINPUT93), .ZN(n473) );
  XNOR2_X1 U584 ( .A(n474), .B(n473), .ZN(n478) );
  XNOR2_X1 U585 ( .A(G143), .B(G131), .ZN(n476) );
  XOR2_X1 U586 ( .A(n731), .B(n479), .Z(n486) );
  NAND2_X1 U587 ( .A1(G214), .A2(n480), .ZN(n482) );
  XNOR2_X1 U588 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U589 ( .A(n484), .B(n483), .Z(n485) );
  XNOR2_X1 U590 ( .A(n486), .B(n485), .ZN(n626) );
  NOR2_X1 U591 ( .A1(G902), .A2(n626), .ZN(n490) );
  XNOR2_X1 U592 ( .A(KEYINPUT13), .B(KEYINPUT94), .ZN(n488) );
  INV_X1 U593 ( .A(G475), .ZN(n487) );
  XNOR2_X1 U594 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U595 ( .A(n493), .B(KEYINPUT9), .Z(n495) );
  XNOR2_X1 U596 ( .A(n495), .B(n494), .ZN(n500) );
  NAND2_X1 U597 ( .A1(G217), .A2(n496), .ZN(n498) );
  XNOR2_X1 U598 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U599 ( .A(n499), .B(n500), .ZN(n709) );
  NAND2_X1 U600 ( .A1(n709), .A2(n501), .ZN(n503) );
  XOR2_X1 U601 ( .A(KEYINPUT96), .B(G478), .Z(n502) );
  NOR2_X1 U602 ( .A1(n530), .A2(n526), .ZN(n573) );
  NAND2_X1 U603 ( .A1(n504), .A2(n573), .ZN(n506) );
  XNOR2_X2 U604 ( .A(n506), .B(n505), .ZN(n743) );
  INV_X1 U605 ( .A(KEYINPUT44), .ZN(n539) );
  NAND2_X1 U606 ( .A1(n743), .A2(n539), .ZN(n507) );
  NAND2_X1 U607 ( .A1(n507), .A2(KEYINPUT66), .ZN(n517) );
  NAND2_X1 U608 ( .A1(n530), .A2(n526), .ZN(n680) );
  NOR2_X1 U609 ( .A1(n680), .A2(n518), .ZN(n508) );
  NAND2_X1 U610 ( .A1(n523), .A2(n508), .ZN(n509) );
  NAND2_X1 U611 ( .A1(n664), .A2(n567), .ZN(n510) );
  XNOR2_X1 U612 ( .A(n510), .B(KEYINPUT101), .ZN(n511) );
  INV_X1 U613 ( .A(n570), .ZN(n513) );
  AND2_X1 U614 ( .A1(n567), .A2(n513), .ZN(n515) );
  INV_X1 U615 ( .A(n567), .ZN(n534) );
  AND2_X1 U616 ( .A1(n534), .A2(n569), .ZN(n519) );
  NAND2_X1 U617 ( .A1(n523), .A2(n519), .ZN(n520) );
  XNOR2_X1 U618 ( .A(n520), .B(KEYINPUT87), .ZN(n521) );
  XNOR2_X1 U619 ( .A(n522), .B(KEYINPUT89), .ZN(n673) );
  INV_X1 U620 ( .A(n523), .ZN(n524) );
  XNOR2_X1 U621 ( .A(KEYINPUT31), .B(KEYINPUT90), .ZN(n525) );
  INV_X1 U622 ( .A(n526), .ZN(n529) );
  NOR2_X1 U623 ( .A1(n530), .A2(n529), .ZN(n528) );
  INV_X1 U624 ( .A(KEYINPUT97), .ZN(n527) );
  XNOR2_X1 U625 ( .A(n528), .B(n527), .ZN(n552) );
  AND2_X1 U626 ( .A1(n530), .A2(n529), .ZN(n638) );
  NOR2_X1 U627 ( .A1(n552), .A2(n638), .ZN(n531) );
  XOR2_X1 U628 ( .A(KEYINPUT98), .B(n531), .Z(n681) );
  NAND2_X1 U629 ( .A1(n536), .A2(KEYINPUT66), .ZN(n538) );
  AND2_X1 U630 ( .A1(n743), .A2(KEYINPUT44), .ZN(n537) );
  NAND2_X1 U631 ( .A1(n539), .A2(KEYINPUT66), .ZN(n540) );
  AND2_X1 U632 ( .A1(n567), .A2(n668), .ZN(n554) );
  NAND2_X1 U633 ( .A1(G953), .A2(G900), .ZN(n541) );
  AND2_X1 U634 ( .A1(n542), .A2(n541), .ZN(n565) );
  XNOR2_X1 U635 ( .A(n544), .B(KEYINPUT105), .ZN(n545) );
  NAND2_X1 U636 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U637 ( .A(n547), .B(KEYINPUT107), .ZN(n584) );
  AND2_X1 U638 ( .A1(n548), .A2(n584), .ZN(n642) );
  NAND2_X1 U639 ( .A1(n681), .A2(n642), .ZN(n551) );
  INV_X1 U640 ( .A(KEYINPUT47), .ZN(n549) );
  NAND2_X1 U641 ( .A1(n549), .A2(KEYINPUT70), .ZN(n550) );
  XNOR2_X1 U642 ( .A(n551), .B(n550), .ZN(n564) );
  AND2_X1 U643 ( .A1(n554), .A2(n565), .ZN(n555) );
  NAND2_X1 U644 ( .A1(n396), .A2(n555), .ZN(n556) );
  BUF_X1 U645 ( .A(n557), .Z(n558) );
  XNOR2_X1 U646 ( .A(n559), .B(KEYINPUT36), .ZN(n560) );
  NAND2_X1 U647 ( .A1(n560), .A2(n664), .ZN(n650) );
  INV_X1 U648 ( .A(KEYINPUT70), .ZN(n561) );
  NAND2_X1 U649 ( .A1(n561), .A2(KEYINPUT47), .ZN(n562) );
  NAND2_X1 U650 ( .A1(n650), .A2(n562), .ZN(n563) );
  NOR2_X1 U651 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U652 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n571) );
  AND2_X1 U653 ( .A1(n596), .A2(n573), .ZN(n574) );
  NAND2_X1 U654 ( .A1(n580), .A2(n574), .ZN(n576) );
  INV_X1 U655 ( .A(KEYINPUT104), .ZN(n575) );
  XNOR2_X1 U656 ( .A(n576), .B(n575), .ZN(n745) );
  XNOR2_X1 U657 ( .A(n745), .B(KEYINPUT75), .ZN(n577) );
  AND2_X1 U658 ( .A1(n578), .A2(n577), .ZN(n590) );
  INV_X1 U659 ( .A(KEYINPUT38), .ZN(n579) );
  NAND2_X2 U660 ( .A1(n582), .A2(n552), .ZN(n583) );
  XNOR2_X2 U661 ( .A(n583), .B(KEYINPUT40), .ZN(n624) );
  NAND2_X1 U662 ( .A1(n678), .A2(n677), .ZN(n683) );
  AND2_X1 U663 ( .A1(n676), .A2(n584), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n624), .A2(n586), .ZN(n588) );
  XNOR2_X1 U665 ( .A(n588), .B(n587), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n592) );
  INV_X1 U667 ( .A(KEYINPUT48), .ZN(n591) );
  XNOR2_X1 U668 ( .A(n592), .B(n591), .ZN(n600) );
  INV_X1 U669 ( .A(n638), .ZN(n646) );
  AND2_X1 U670 ( .A1(n593), .A2(n677), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n594), .A2(n514), .ZN(n595) );
  XNOR2_X1 U672 ( .A(n595), .B(KEYINPUT43), .ZN(n598) );
  INV_X1 U673 ( .A(n596), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n652) );
  AND2_X1 U675 ( .A1(n623), .A2(n652), .ZN(n599) );
  INV_X1 U676 ( .A(KEYINPUT2), .ZN(n654) );
  INV_X1 U677 ( .A(n601), .ZN(n603) );
  INV_X1 U678 ( .A(KEYINPUT77), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(KEYINPUT77), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n604), .A2(n654), .ZN(n605) );
  XNOR2_X2 U681 ( .A(n608), .B(KEYINPUT65), .ZN(n711) );
  NAND2_X1 U682 ( .A1(n711), .A2(G210), .ZN(n612) );
  XOR2_X1 U683 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n610) );
  XOR2_X1 U684 ( .A(n610), .B(KEYINPUT80), .Z(n611) );
  XNOR2_X1 U685 ( .A(n612), .B(n412), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U687 ( .A1(n711), .A2(G472), .ZN(n617) );
  XNOR2_X1 U688 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n620), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U691 ( .A(G110), .B(KEYINPUT111), .Z(n621) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(G12) );
  XNOR2_X1 U693 ( .A(n623), .B(G134), .ZN(G36) );
  XNOR2_X1 U694 ( .A(n624), .B(G131), .ZN(G33) );
  NAND2_X1 U695 ( .A1(n711), .A2(G475), .ZN(n628) );
  XNOR2_X1 U696 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X2 U698 ( .A1(n629), .A2(n717), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n630), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X1 U700 ( .A1(n634), .A2(n644), .ZN(n632) );
  XOR2_X1 U701 ( .A(KEYINPUT110), .B(n632), .Z(n633) );
  XNOR2_X1 U702 ( .A(G104), .B(n633), .ZN(G6) );
  NOR2_X1 U703 ( .A1(n634), .A2(n646), .ZN(n636) );
  XNOR2_X1 U704 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(G107), .B(n637), .ZN(G9) );
  XOR2_X1 U707 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n640) );
  NAND2_X1 U708 ( .A1(n642), .A2(n638), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U710 ( .A(G128), .B(n641), .ZN(G30) );
  NAND2_X1 U711 ( .A1(n642), .A2(n552), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(G146), .ZN(G48) );
  NOR2_X1 U713 ( .A1(n647), .A2(n644), .ZN(n645) );
  XOR2_X1 U714 ( .A(G113), .B(n645), .Z(G15) );
  NOR2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U716 ( .A(G116), .B(n648), .Z(G18) );
  XOR2_X1 U717 ( .A(G125), .B(KEYINPUT37), .Z(n649) );
  XNOR2_X1 U718 ( .A(n650), .B(n649), .ZN(G27) );
  XNOR2_X1 U719 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U720 ( .A(n653), .B(KEYINPUT113), .ZN(G42) );
  NAND2_X1 U721 ( .A1(n718), .A2(n654), .ZN(n655) );
  NAND2_X1 U722 ( .A1(n656), .A2(n655), .ZN(n660) );
  NOR2_X1 U723 ( .A1(n733), .A2(KEYINPUT2), .ZN(n658) );
  XOR2_X1 U724 ( .A(KEYINPUT76), .B(n658), .Z(n659) );
  NAND2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U726 ( .A1(n676), .A2(n688), .ZN(n661) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n698) );
  NAND2_X1 U728 ( .A1(G952), .A2(n663), .ZN(n695) );
  XNOR2_X1 U729 ( .A(KEYINPUT116), .B(KEYINPUT52), .ZN(n693) );
  NOR2_X1 U730 ( .A1(n349), .A2(n664), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n665), .B(KEYINPUT50), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n534), .A2(n668), .ZN(n669) );
  XNOR2_X1 U734 ( .A(n669), .B(KEYINPUT49), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U737 ( .A(KEYINPUT51), .B(n674), .Z(n675) );
  NAND2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n690) );
  NOR2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n686) );
  INV_X1 U741 ( .A(n681), .ZN(n682) );
  NOR2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U743 ( .A(KEYINPUT114), .B(n684), .ZN(n685) );
  OR2_X1 U744 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U745 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U746 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U747 ( .A(n691), .B(KEYINPUT115), .ZN(n692) );
  XNOR2_X1 U748 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U749 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U750 ( .A(KEYINPUT117), .B(n696), .Z(n697) );
  NOR2_X1 U751 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U752 ( .A1(n734), .A2(n699), .ZN(n700) );
  XOR2_X1 U753 ( .A(KEYINPUT53), .B(n700), .Z(G75) );
  BUF_X1 U754 ( .A(n711), .Z(n701) );
  NAND2_X1 U755 ( .A1(n701), .A2(G469), .ZN(n706) );
  XNOR2_X1 U756 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n702) );
  XOR2_X1 U757 ( .A(n702), .B(KEYINPUT57), .Z(n703) );
  XNOR2_X1 U758 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n717), .A2(n707), .ZN(G54) );
  NAND2_X1 U761 ( .A1(n711), .A2(G478), .ZN(n708) );
  XOR2_X1 U762 ( .A(n709), .B(n708), .Z(n710) );
  NOR2_X1 U763 ( .A1(n717), .A2(n710), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n701), .A2(G217), .ZN(n715) );
  XOR2_X1 U765 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n712) );
  NOR2_X1 U766 ( .A1(n717), .A2(n716), .ZN(G66) );
  NAND2_X1 U767 ( .A1(n718), .A2(n734), .ZN(n723) );
  NAND2_X1 U768 ( .A1(G224), .A2(G953), .ZN(n719) );
  XNOR2_X1 U769 ( .A(n719), .B(KEYINPUT61), .ZN(n720) );
  XNOR2_X1 U770 ( .A(KEYINPUT122), .B(n720), .ZN(n721) );
  NAND2_X1 U771 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n729) );
  XOR2_X1 U773 ( .A(KEYINPUT124), .B(n724), .Z(n726) );
  NOR2_X1 U774 ( .A1(G898), .A2(n734), .ZN(n725) );
  NOR2_X1 U775 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U776 ( .A(KEYINPUT123), .B(n727), .Z(n728) );
  XNOR2_X1 U777 ( .A(n729), .B(n728), .ZN(n730) );
  XOR2_X1 U778 ( .A(KEYINPUT125), .B(n730), .Z(G69) );
  XNOR2_X1 U779 ( .A(n732), .B(n731), .ZN(n736) );
  XNOR2_X1 U780 ( .A(n733), .B(n736), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n735), .A2(n734), .ZN(n741) );
  XOR2_X1 U782 ( .A(G227), .B(n736), .Z(n737) );
  NAND2_X1 U783 ( .A1(n737), .A2(G900), .ZN(n738) );
  XNOR2_X1 U784 ( .A(KEYINPUT126), .B(n738), .ZN(n739) );
  NAND2_X1 U785 ( .A1(G953), .A2(n739), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n741), .A2(n740), .ZN(G72) );
  XOR2_X1 U787 ( .A(G122), .B(KEYINPUT127), .Z(n742) );
  XNOR2_X1 U788 ( .A(n743), .B(n742), .ZN(G24) );
  XNOR2_X1 U789 ( .A(G101), .B(n744), .ZN(G3) );
  XOR2_X1 U790 ( .A(G143), .B(n745), .Z(G45) );
endmodule

