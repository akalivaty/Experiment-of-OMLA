//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT5), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n204));
  XOR2_X1   g003(.A(G141gat), .B(G148gat), .Z(new_n205));
  XNOR2_X1  g004(.A(G155gat), .B(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT2), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n206), .B1(new_n205), .B2(new_n209), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n204), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n212), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT76), .A3(new_n210), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT3), .ZN(new_n216));
  INV_X1    g015(.A(G134gat), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT1), .B1(new_n217), .B2(G127gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n219));
  INV_X1    g018(.A(G120gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G113gat), .ZN(new_n221));
  OAI221_X1 g020(.A(new_n218), .B1(G127gat), .B2(new_n217), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G113gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G120gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n221), .A2(new_n224), .A3(new_n219), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT70), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n225), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n221), .A2(new_n219), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n217), .A2(G127gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT70), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .A4(new_n218), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT68), .B(G134gat), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n234), .A2(G127gat), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n221), .A2(new_n224), .ZN(new_n236));
  OAI22_X1  g035(.A1(new_n235), .A2(new_n229), .B1(KEYINPUT1), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n211), .A2(new_n212), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n216), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT77), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n216), .A2(new_n238), .A3(new_n244), .A4(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n233), .A2(new_n239), .A3(new_n237), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n248), .A2(KEYINPUT4), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(KEYINPUT4), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n213), .A2(new_n215), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n238), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n247), .B1(new_n254), .B2(new_n248), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n203), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n243), .A2(new_n245), .B1(new_n249), .B2(new_n250), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT5), .B1(new_n258), .B2(new_n247), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT6), .ZN(new_n260));
  XOR2_X1   g059(.A(G1gat), .B(G29gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(G85gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT0), .B(G57gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NOR4_X1   g064(.A1(new_n257), .A2(new_n259), .A3(new_n260), .A4(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n203), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n255), .B1(new_n258), .B2(new_n247), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(new_n203), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT6), .B1(new_n270), .B2(new_n265), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT78), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n268), .B(new_n264), .C1(new_n269), .C2(new_n203), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n271), .A2(new_n272), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n267), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G183gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT64), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G183gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n281), .A3(KEYINPUT27), .ZN(new_n282));
  OR2_X1    g081(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n283));
  AOI21_X1  g082(.A(G190gat), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT65), .B1(new_n284), .B2(KEYINPUT28), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n287));
  NOR2_X1   g086(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT64), .B(G183gat), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(KEYINPUT27), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n286), .B(new_n287), .C1(new_n290), .C2(G190gat), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n283), .A2(KEYINPUT66), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT66), .B1(new_n283), .B2(new_n293), .ZN(new_n295));
  OAI211_X1 g094(.A(KEYINPUT28), .B(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT26), .ZN(new_n299));
  NAND2_X1  g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT26), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n299), .B(new_n300), .C1(new_n303), .C2(new_n298), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n298), .A2(KEYINPUT23), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n298), .A2(KEYINPUT23), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n289), .A2(G190gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n300), .B(KEYINPUT24), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n310), .B(KEYINPUT25), .C1(new_n311), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n278), .A2(new_n292), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(new_n309), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n314), .B1(new_n317), .B2(KEYINPUT25), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n306), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n297), .A2(KEYINPUT67), .A3(new_n305), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT67), .B1(new_n297), .B2(new_n305), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n318), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n328));
  XNOR2_X1  g127(.A(G197gat), .B(G204gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330));
  INV_X1    g129(.A(G211gat), .ZN(new_n331));
  INV_X1    g130(.A(G218gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n328), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT75), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(new_n329), .A3(new_n333), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n328), .A2(new_n334), .A3(new_n341), .A4(new_n337), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n319), .A2(new_n325), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(new_n324), .B2(new_n320), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n343), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT30), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(new_n352), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT30), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n349), .B2(new_n352), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n277), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n324), .A2(new_n238), .ZN(new_n361));
  INV_X1    g160(.A(new_n238), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n362), .B(new_n318), .C1(new_n322), .C2(new_n323), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT34), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n364), .B2(new_n366), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT67), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n306), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n297), .A2(KEYINPUT67), .A3(new_n305), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n362), .B1(new_n376), .B2(new_n318), .ZN(new_n377));
  INV_X1    g176(.A(new_n363), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n366), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT32), .ZN(new_n380));
  XNOR2_X1  g179(.A(G15gat), .B(G43gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT33), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n379), .A2(new_n385), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n388), .B2(KEYINPUT71), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT33), .B1(new_n364), .B2(new_n366), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT71), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n390), .A2(new_n391), .B1(KEYINPUT32), .B2(new_n379), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n387), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n372), .B1(new_n393), .B2(KEYINPUT73), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n391), .A3(new_n385), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n365), .B1(new_n361), .B2(new_n363), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT71), .B1(new_n396), .B2(KEYINPUT33), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n395), .A2(new_n397), .A3(new_n380), .A4(new_n383), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n380), .A2(new_n386), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT73), .ZN(new_n401));
  INV_X1    g200(.A(new_n372), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n394), .A2(KEYINPUT36), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT36), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n398), .A2(new_n399), .A3(new_n372), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n372), .B1(new_n398), .B2(new_n399), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n334), .A2(new_n327), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n340), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT3), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n239), .B2(new_n240), .ZN(new_n416));
  OAI221_X1 g215(.A(new_n411), .B1(new_n415), .B2(new_n239), .C1(new_n416), .C2(new_n343), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n343), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n343), .A2(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n240), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n420), .B2(new_n253), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n417), .B1(new_n421), .B2(new_n411), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G22gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n424));
  INV_X1    g223(.A(G22gat), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n425), .B(new_n417), .C1(new_n421), .C2(new_n411), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(G78gat), .B(G106gat), .Z(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n428), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n423), .A2(new_n424), .A3(new_n426), .A4(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n429), .B2(new_n432), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n410), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n429), .A2(new_n432), .ZN(new_n438));
  INV_X1    g237(.A(new_n430), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n433), .ZN(new_n441));
  AND4_X1   g240(.A1(KEYINPUT35), .A2(new_n441), .A3(new_n394), .A4(new_n403), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n360), .B1(new_n437), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT82), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n407), .B2(new_n408), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n400), .A2(new_n402), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(KEYINPUT82), .A3(new_n406), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n358), .B1(new_n440), .B2(new_n433), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n266), .B1(new_n271), .B2(new_n274), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n446), .A2(new_n448), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT35), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT38), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n344), .B(new_n346), .C1(new_n324), .C2(new_n320), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(KEYINPUT37), .A3(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n324), .A2(new_n325), .ZN(new_n460));
  OAI211_X1 g259(.A(KEYINPUT80), .B(new_n343), .C1(new_n460), .C2(new_n321), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT80), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n326), .B2(new_n344), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT37), .B1(new_n345), .B2(new_n348), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n455), .B(new_n352), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n345), .A2(new_n348), .A3(KEYINPUT37), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n352), .B1(new_n468), .B2(new_n466), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n353), .B1(new_n469), .B2(KEYINPUT38), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(new_n470), .A3(new_n450), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n258), .A2(KEYINPUT39), .A3(new_n247), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(new_n264), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n254), .A2(new_n247), .A3(new_n248), .ZN(new_n474));
  OAI211_X1 g273(.A(KEYINPUT39), .B(new_n474), .C1(new_n258), .C2(new_n247), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n473), .A2(KEYINPUT40), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT40), .B1(new_n473), .B2(new_n475), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(new_n358), .A3(new_n274), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n436), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n410), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n454), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n202), .B1(new_n444), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n441), .B1(new_n404), .B2(new_n409), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n277), .B(new_n359), .C1(new_n484), .C2(new_n442), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n453), .A2(new_n452), .B1(new_n410), .B2(new_n480), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT83), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT16), .ZN(new_n490));
  INV_X1    g289(.A(G1gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT87), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G1gat), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G1gat), .B2(new_n498), .ZN(new_n500));
  INV_X1    g299(.A(G8gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR3_X1   g304(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  XOR2_X1   g307(.A(G43gat), .B(G50gat), .Z(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT84), .B1(new_n509), .B2(new_n508), .ZN(new_n511));
  OR3_X1    g310(.A1(new_n509), .A2(KEYINPUT84), .A3(new_n508), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n509), .A2(new_n508), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT86), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT17), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(KEYINPUT17), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n518), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n502), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n502), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n518), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT18), .A3(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n502), .B(new_n518), .Z(new_n530));
  XOR2_X1   g329(.A(new_n528), .B(KEYINPUT13), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537));
  INV_X1    g336(.A(G197gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT11), .B(G169gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n541), .B(KEYINPUT12), .Z(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n542), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n529), .A2(new_n532), .A3(new_n535), .A4(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G57gat), .B(G64gat), .Z(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(KEYINPUT89), .B2(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT89), .Z(new_n551));
  NOR2_X1   g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT90), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n552), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g356(.A(new_n550), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n548), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G211gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n562), .B(new_n564), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n502), .B1(new_n561), .B2(new_n560), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G183gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT92), .Z(new_n572));
  NOR2_X1   g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n569), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n568), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n572), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n566), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n570), .A2(new_n572), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n565), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G134gat), .B(G162gat), .Z(new_n583));
  AOI21_X1  g382(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT7), .ZN(new_n588));
  INV_X1    g387(.A(G99gat), .ZN(new_n589));
  INV_X1    g388(.A(G106gat), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT8), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT93), .B(G85gat), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n588), .B(new_n591), .C1(G92gat), .C2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G99gat), .B(G106gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n522), .B2(new_n523), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT94), .ZN(new_n597));
  AND3_X1   g396(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n595), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n518), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n601), .B(new_n595), .C1(new_n522), .C2(new_n523), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n586), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT95), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n606), .B(new_n607), .C1(new_n605), .C2(new_n603), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n605), .A3(new_n586), .ZN(new_n609));
  INV_X1    g408(.A(new_n603), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n610), .B(new_n604), .C1(KEYINPUT95), .C2(new_n586), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n560), .A2(new_n595), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n599), .A2(new_n556), .A3(new_n559), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n623), .A2(new_n622), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n620), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n619), .B1(new_n621), .B2(new_n623), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n617), .B(new_n618), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n626), .A2(new_n627), .A3(new_n615), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n629), .A2(KEYINPUT96), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(KEYINPUT96), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n582), .A2(new_n612), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n489), .A2(new_n547), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT98), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n489), .A2(new_n636), .A3(new_n547), .A4(new_n633), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n277), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g440(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G8gat), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n638), .A2(new_n358), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT100), .B1(new_n644), .B2(KEYINPUT42), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n501), .B1(new_n638), .B2(new_n358), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(new_n644), .B2(KEYINPUT42), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n638), .A2(new_n358), .A3(new_n643), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n647), .A3(new_n651), .ZN(G1325gat));
  NAND2_X1  g451(.A1(new_n446), .A2(new_n448), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(G15gat), .B1(new_n638), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n410), .B1(new_n635), .B2(new_n637), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(G15gat), .B2(new_n656), .ZN(G1326gat));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n638), .B2(new_n436), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AOI211_X1 g459(.A(KEYINPUT101), .B(new_n441), .C1(new_n635), .C2(new_n637), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT43), .B(G22gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n659), .B2(new_n661), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(G1327gat));
  NAND2_X1  g466(.A1(new_n578), .A2(new_n581), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(new_n546), .A3(new_n632), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n489), .A2(new_n612), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n670), .A2(G29gat), .A3(new_n277), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT45), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n483), .A2(new_n487), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n612), .B1(new_n444), .B2(new_n482), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n674), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n669), .B(KEYINPUT102), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G29gat), .B1(new_n681), .B2(new_n277), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n672), .A2(new_n682), .ZN(G1328gat));
  NOR3_X1   g482(.A1(new_n670), .A2(G36gat), .A3(new_n359), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT46), .ZN(new_n685));
  OAI21_X1  g484(.A(G36gat), .B1(new_n681), .B2(new_n359), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(G1329gat));
  INV_X1    g486(.A(G43gat), .ZN(new_n688));
  INV_X1    g487(.A(new_n410), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n679), .A2(new_n689), .A3(new_n680), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n690), .B2(KEYINPUT104), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(KEYINPUT104), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n670), .A2(new_n653), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT103), .B1(new_n693), .B2(new_n688), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n693), .A2(KEYINPUT103), .A3(new_n688), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n692), .B(KEYINPUT47), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n690), .A2(G43gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(new_n695), .B2(new_n694), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT47), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n696), .A2(new_n700), .ZN(G1330gat));
  NAND3_X1  g500(.A1(new_n679), .A2(G50gat), .A3(new_n680), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n670), .A2(new_n441), .ZN(new_n703));
  OAI22_X1  g502(.A1(new_n441), .A2(new_n702), .B1(new_n703), .B2(G50gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g504(.A1(new_n485), .A2(new_n486), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n668), .A3(new_n673), .ZN(new_n707));
  INV_X1    g506(.A(new_n632), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n707), .A2(new_n547), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n639), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT105), .B(G57gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1332gat));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n358), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT49), .B(G64gat), .Z(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(G1333gat));
  XNOR2_X1  g515(.A(new_n653), .B(KEYINPUT106), .ZN(new_n717));
  AOI21_X1  g516(.A(G71gat), .B1(new_n709), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n689), .A2(G71gat), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n709), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g520(.A1(new_n709), .A2(new_n436), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g522(.A1(new_n668), .A2(new_n547), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n706), .A2(new_n612), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n706), .A2(KEYINPUT51), .A3(new_n612), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT108), .Z(new_n730));
  INV_X1    g529(.A(new_n592), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n731), .A3(new_n632), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n668), .A2(new_n547), .A3(new_n708), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n676), .A2(new_n678), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT107), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n676), .A2(new_n678), .A3(new_n736), .A4(new_n733), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n277), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n732), .A2(new_n277), .B1(new_n731), .B2(new_n738), .ZN(G1336gat));
  INV_X1    g538(.A(G92gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n737), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n358), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n729), .A2(new_n740), .A3(new_n632), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n359), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT52), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n676), .A2(new_n678), .A3(new_n358), .A4(new_n733), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G92gat), .B1(new_n749), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n743), .B2(new_n359), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n748), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  AOI211_X1 g555(.A(G92gat), .B(new_n708), .C1(new_n727), .C2(new_n728), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(new_n757), .B2(new_n358), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n758), .B(KEYINPUT111), .C1(new_n751), .C2(new_n752), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(KEYINPUT109), .B(KEYINPUT52), .C1(new_n742), .C2(new_n744), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n747), .A2(new_n760), .A3(new_n761), .ZN(G1337gat));
  NAND3_X1  g561(.A1(new_n654), .A2(new_n589), .A3(new_n632), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n730), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n410), .B1(new_n735), .B2(new_n737), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n589), .B2(new_n766), .ZN(G1338gat));
  AOI21_X1  g566(.A(new_n590), .B1(new_n741), .B2(new_n436), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n729), .A2(new_n590), .A3(new_n632), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n441), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT53), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n679), .A2(KEYINPUT113), .A3(new_n436), .A4(new_n733), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n734), .B2(new_n441), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n772), .A2(G106gat), .A3(new_n774), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n770), .A2(KEYINPUT53), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n771), .B1(new_n775), .B2(new_n776), .ZN(G1339gat));
  NOR2_X1   g576(.A1(new_n527), .A2(new_n528), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n530), .A2(new_n531), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n541), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n545), .A2(new_n780), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n624), .A2(new_n625), .A3(new_n620), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  OR3_X1    g582(.A1(new_n782), .A2(new_n626), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n616), .B1(new_n626), .B2(new_n783), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n784), .A2(KEYINPUT55), .A3(new_n785), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n788), .B(new_n789), .C1(new_n630), .C2(new_n631), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n612), .B1(new_n781), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n632), .A2(new_n545), .A3(new_n780), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n673), .B(new_n792), .C1(new_n546), .C2(new_n790), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n582), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n668), .A2(new_n546), .A3(new_n673), .A4(new_n708), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT114), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n653), .A2(new_n436), .A3(new_n358), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n639), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n800), .A2(new_n804), .A3(new_n639), .A4(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G113gat), .B1(new_n806), .B2(new_n546), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n441), .A2(new_n394), .A3(new_n403), .ZN(new_n808));
  AND4_X1   g607(.A1(new_n639), .A2(new_n800), .A3(new_n808), .A4(new_n359), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n223), .A3(new_n547), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(G1340gat));
  OAI21_X1  g610(.A(G120gat), .B1(new_n806), .B2(new_n708), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n220), .A3(new_n632), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n812), .A2(KEYINPUT116), .A3(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1341gat));
  INV_X1    g617(.A(G127gat), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n806), .A2(new_n819), .A3(new_n582), .ZN(new_n820));
  AOI21_X1  g619(.A(G127gat), .B1(new_n809), .B2(new_n668), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(G1342gat));
  NAND3_X1  g621(.A1(new_n809), .A2(new_n234), .A3(new_n612), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n824));
  OAI21_X1  g623(.A(G134gat), .B1(new_n806), .B2(new_n673), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(G1343gat));
  NAND2_X1  g626(.A1(new_n800), .A2(new_n436), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(G141gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n639), .A2(new_n359), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n689), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n829), .A2(new_n830), .A3(new_n547), .A4(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n797), .A2(new_n834), .A3(new_n436), .A4(new_n799), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n832), .B(KEYINPUT117), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n796), .A2(new_n436), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT57), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n835), .A2(new_n836), .A3(new_n547), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n839), .B2(G141gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT119), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT118), .A4(new_n838), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n830), .B1(new_n847), .B2(new_n547), .ZN(new_n848));
  INV_X1    g647(.A(new_n833), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT58), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n842), .A2(new_n850), .ZN(G1344gat));
  NOR3_X1   g650(.A1(new_n828), .A2(new_n689), .A3(new_n831), .ZN(new_n852));
  INV_X1    g651(.A(G148gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n632), .ZN(new_n854));
  AOI211_X1 g653(.A(KEYINPUT59), .B(new_n853), .C1(new_n847), .C2(new_n632), .ZN(new_n855));
  XNOR2_X1  g654(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n837), .A2(new_n834), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n828), .B2(new_n834), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n632), .A3(new_n836), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n859), .B2(G148gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n854), .B1(new_n855), .B2(new_n860), .ZN(G1345gat));
  NAND3_X1  g660(.A1(new_n852), .A2(new_n207), .A3(new_n668), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n582), .B1(new_n845), .B2(new_n846), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n207), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(G1346gat));
  AOI21_X1  g665(.A(G162gat), .B1(new_n852), .B2(new_n612), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n673), .B1(new_n845), .B2(new_n846), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n639), .A2(new_n359), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n800), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n808), .ZN(new_n872));
  OR3_X1    g671(.A1(new_n872), .A2(G169gat), .A3(new_n546), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n441), .A3(new_n717), .ZN(new_n874));
  OAI21_X1  g673(.A(G169gat), .B1(new_n874), .B2(new_n546), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1348gat));
  INV_X1    g675(.A(G176gat), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n874), .A2(new_n877), .A3(new_n708), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n872), .B2(new_n708), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT122), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(KEYINPUT122), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(G1349gat));
  INV_X1    g681(.A(new_n872), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n294), .A2(new_n295), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n884), .A3(new_n668), .ZN(new_n885));
  INV_X1    g684(.A(new_n289), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n874), .A2(new_n582), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT60), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n885), .B(new_n890), .C1(new_n886), .C2(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n874), .B2(new_n673), .ZN(new_n893));
  XOR2_X1   g692(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n883), .A2(new_n292), .A3(new_n612), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1351gat));
  NAND2_X1  g696(.A1(new_n870), .A2(new_n410), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n858), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G197gat), .B1(new_n900), .B2(new_n546), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n800), .A2(new_n484), .A3(new_n870), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n538), .A3(new_n547), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1352gat));
  XOR2_X1   g703(.A(KEYINPUT124), .B(G204gat), .Z(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n632), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n902), .A2(new_n909), .A3(new_n632), .A4(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT126), .B1(new_n911), .B2(KEYINPUT62), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT62), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n858), .A2(new_n632), .A3(new_n899), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n905), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n908), .A2(new_n916), .A3(new_n910), .A4(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n912), .A2(new_n913), .A3(new_n915), .A4(new_n918), .ZN(G1353gat));
  NAND3_X1  g718(.A1(new_n858), .A2(new_n668), .A3(new_n899), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G211gat), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT63), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n902), .A2(new_n331), .A3(new_n668), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(KEYINPUT63), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n922), .A2(KEYINPUT63), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n920), .A2(G211gat), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n924), .A3(new_n927), .ZN(G1354gat));
  OAI21_X1  g727(.A(G218gat), .B1(new_n900), .B2(new_n673), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n902), .A2(new_n332), .A3(new_n612), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1355gat));
endmodule


