//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n226), .A2(new_n227), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n211), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n214), .B(new_n220), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  AOI21_X1  g0052(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  AOI21_X1  g0057(.A(G1), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n253), .A2(new_n258), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(KEYINPUT73), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n223), .B1(new_n261), .B2(KEYINPUT73), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  OAI211_X1 g0066(.A(G232), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(G232), .A4(G1698), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G97), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n269), .A2(G226), .A3(new_n273), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n268), .A2(new_n271), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n275), .A2(KEYINPUT72), .A3(new_n253), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT72), .B1(new_n275), .B2(new_n253), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n264), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT13), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n280), .B(new_n264), .C1(new_n276), .C2(new_n277), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G190), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n222), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT12), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n209), .A2(G33), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n288), .B1(new_n224), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n218), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(KEYINPUT11), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n292), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n283), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n208), .A2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G68), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n286), .B(new_n293), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT11), .B1(new_n290), .B2(new_n292), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n282), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n279), .B2(new_n281), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n275), .A2(new_n253), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n275), .A2(KEYINPUT72), .A3(new_n253), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n280), .B1(new_n310), .B2(new_n264), .ZN(new_n311));
  INV_X1    g0111(.A(new_n281), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n305), .B(G169), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n279), .A2(G179), .A3(new_n281), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(G169), .B1(new_n311), .B2(new_n312), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT74), .B1(new_n316), .B2(KEYINPUT14), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n279), .B2(new_n281), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT74), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n319), .A2(new_n320), .A3(new_n305), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n315), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n300), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n304), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT8), .B(G58), .ZN(new_n326));
  INV_X1    g0126(.A(G150), .ZN(new_n327));
  INV_X1    g0127(.A(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n209), .A2(new_n328), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n326), .A2(new_n289), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(G20), .B2(new_n203), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n294), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n296), .A2(G50), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n295), .A2(new_n333), .B1(G50), .B2(new_n283), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT9), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n335), .B(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(G1), .B(G13), .C1(new_n328), .C2(new_n256), .ZN(new_n338));
  OR2_X1    g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NAND2_X1  g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  AOI21_X1  g0140(.A(G1698), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G222), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT68), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n269), .A2(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n265), .A2(new_n266), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n345), .A2(G223), .B1(G77), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n338), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  XOR2_X1   g0148(.A(KEYINPUT67), .B(G226), .Z(new_n349));
  AND2_X1   g0149(.A1(new_n261), .A2(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n260), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G190), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n337), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT10), .ZN(new_n355));
  INV_X1    g0155(.A(new_n352), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(KEYINPUT70), .A3(G200), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n352), .B2(new_n302), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n354), .A2(new_n355), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n357), .A2(new_n359), .A3(new_n353), .A4(new_n337), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT10), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n326), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n296), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n365), .A2(new_n295), .B1(new_n283), .B2(new_n364), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT78), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n339), .A2(new_n209), .A3(new_n340), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n346), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G68), .ZN(new_n373));
  INV_X1    g0173(.A(G58), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(new_n222), .ZN(new_n375));
  OAI21_X1  g0175(.A(G20), .B1(new_n375), .B2(new_n201), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n287), .A2(KEYINPUT75), .A3(G159), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT75), .B1(new_n287), .B2(G159), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n373), .A2(KEYINPUT16), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n380), .B1(new_n372), .B2(G68), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT16), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n294), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT77), .B1(new_n370), .B2(new_n371), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT77), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n368), .B2(new_n369), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT16), .B1(new_n391), .B2(new_n381), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n367), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n341), .A2(G223), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT79), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n341), .A2(KEYINPUT79), .A3(G223), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G226), .ZN(new_n400));
  INV_X1    g0200(.A(G87), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n344), .A2(new_n400), .B1(new_n328), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n338), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n261), .ZN(new_n405));
  INV_X1    g0205(.A(G232), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n259), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(G169), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n407), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n402), .B1(new_n397), .B2(new_n398), .ZN(new_n410));
  OAI211_X1 g0210(.A(G179), .B(new_n409), .C1(new_n410), .C2(new_n338), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT18), .B1(new_n394), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n367), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n385), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n222), .B1(new_n370), .B2(new_n371), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT16), .ZN(new_n418));
  NOR4_X1   g0218(.A1(new_n417), .A2(new_n380), .A3(KEYINPUT76), .A4(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n292), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n415), .B1(new_n420), .B2(new_n392), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n412), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  OAI21_X1  g0225(.A(G200), .B1(new_n404), .B2(new_n407), .ZN(new_n426));
  OAI211_X1 g0226(.A(G190), .B(new_n409), .C1(new_n410), .C2(new_n338), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n425), .B1(new_n421), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n428), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n394), .A2(KEYINPUT17), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n424), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n352), .A2(G169), .ZN(new_n434));
  INV_X1    g0234(.A(G179), .ZN(new_n435));
  AOI211_X1 g0235(.A(new_n335), .B(new_n434), .C1(new_n435), .C2(new_n352), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n326), .A2(new_n329), .B1(new_n209), .B2(new_n224), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT15), .B(G87), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(new_n289), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n292), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n296), .A2(G77), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n441), .B1(G77), .B2(new_n283), .C1(new_n295), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n345), .A2(G238), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n341), .A2(G232), .B1(new_n346), .B2(G107), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n338), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n259), .B1(new_n405), .B2(new_n225), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n443), .B1(new_n449), .B2(G200), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n448), .A2(KEYINPUT69), .A3(G190), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT69), .B1(new_n448), .B2(G190), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n448), .A2(new_n435), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n443), .C1(G169), .C2(new_n448), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n363), .A2(new_n433), .A3(new_n437), .A4(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n325), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G190), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n208), .A2(G45), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT5), .B(G41), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n253), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n464), .A2(new_n463), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n465), .A2(G264), .B1(new_n466), .B2(new_n255), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n269), .A2(G257), .A3(G1698), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n269), .A2(G250), .A3(new_n273), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G294), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT86), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(new_n253), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n472), .B1(new_n471), .B2(new_n253), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n461), .B(new_n467), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n477));
  INV_X1    g0277(.A(new_n467), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n471), .A2(new_n253), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT86), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n480), .B2(new_n473), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT87), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(new_n461), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n467), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n302), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n477), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n401), .A2(KEYINPUT85), .A3(G20), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n269), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n269), .A2(KEYINPUT22), .A3(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G116), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(G20), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT23), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n209), .B2(G107), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(KEYINPUT23), .A3(G20), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n490), .A2(new_n491), .A3(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n499), .A2(KEYINPUT24), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(KEYINPUT24), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n292), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT25), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n283), .B2(G107), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n283), .A2(new_n503), .A3(G107), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n208), .A2(G33), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n283), .A2(new_n507), .A3(new_n218), .A4(new_n291), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n505), .A2(new_n506), .B1(new_n496), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n486), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n479), .A2(new_n467), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G179), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n481), .B2(new_n318), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n511), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G264), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT84), .B1(new_n344), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT84), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n269), .A2(new_n521), .A3(G264), .A4(G1698), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n269), .A2(G257), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n273), .B1(G303), .B2(new_n346), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n253), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n464), .A2(new_n463), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(G270), .A3(new_n338), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT83), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT83), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n465), .A2(new_n531), .A3(G270), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n466), .A2(new_n255), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G283), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT81), .ZN(new_n539));
  INV_X1    g0339(.A(G97), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n209), .B1(new_n540), .B2(G33), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G116), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G20), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n292), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(KEYINPUT20), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT20), .ZN(new_n549));
  OR2_X1    g0349(.A1(new_n538), .A2(KEYINPUT81), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n538), .A2(KEYINPUT81), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n541), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n552), .B2(new_n546), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n283), .A2(G116), .ZN(new_n555));
  INV_X1    g0355(.A(new_n508), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(G116), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n537), .B(new_n559), .C1(new_n536), .C2(new_n461), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n338), .B1(new_n523), .B2(new_n525), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n558), .B(G169), .C1(new_n561), .C2(new_n534), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT21), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT21), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n318), .B1(new_n554), .B2(new_n557), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n536), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n561), .A2(new_n435), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n535), .A3(new_n558), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n560), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G107), .B1(new_n388), .B2(new_n390), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n496), .A2(KEYINPUT6), .A3(G97), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n540), .A2(new_n496), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(new_n205), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n574), .B2(KEYINPUT6), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(G20), .B1(G77), .B2(new_n287), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n292), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n283), .A2(new_n540), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n556), .B2(new_n540), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n580), .B(KEYINPUT80), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(G250), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n583));
  OAI211_X1 g0383(.A(G244), .B(new_n273), .C1(new_n265), .C2(new_n266), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT4), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n539), .B(new_n583), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT4), .B1(new_n341), .B2(G244), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n253), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n465), .A2(G257), .B1(new_n466), .B2(new_n255), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G200), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(G190), .A3(new_n589), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n578), .A2(new_n582), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n318), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n588), .A2(new_n435), .A3(new_n589), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n294), .B1(new_n571), .B2(new_n576), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n594), .B(new_n595), .C1(new_n596), .C2(new_n581), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n269), .A2(G244), .A3(G1698), .ZN(new_n599));
  OAI211_X1 g0399(.A(G238), .B(new_n273), .C1(new_n265), .C2(new_n266), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n492), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n253), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n338), .A2(G250), .A3(new_n462), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n338), .A2(G274), .A3(new_n463), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(new_n435), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n209), .B1(new_n272), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G87), .B2(new_n206), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n608), .B1(new_n289), .B2(new_n540), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n209), .B(G68), .C1(new_n265), .C2(new_n266), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n292), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n439), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n439), .A2(new_n615), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n556), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n439), .A2(new_n284), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n605), .B1(new_n601), .B2(new_n253), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n607), .B(new_n620), .C1(G169), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n602), .A2(new_n606), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(G190), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n556), .A2(G87), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n614), .A2(new_n619), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n598), .A2(new_n622), .A3(new_n628), .ZN(new_n629));
  NOR4_X1   g0429(.A1(new_n460), .A2(new_n518), .A3(new_n570), .A4(new_n629), .ZN(G372));
  INV_X1    g0430(.A(KEYINPUT90), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n394), .A2(new_n413), .A3(KEYINPUT18), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n422), .B1(new_n421), .B2(new_n412), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n414), .A2(KEYINPUT90), .A3(new_n423), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n313), .A2(new_n314), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n320), .B1(new_n319), .B2(new_n305), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n316), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n641), .A2(new_n300), .B1(new_n304), .B2(new_n455), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT91), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n432), .B1(new_n642), .B2(new_n643), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n637), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n363), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n628), .A2(new_n622), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT88), .ZN(new_n650));
  INV_X1    g0450(.A(new_n597), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT88), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n628), .A2(new_n653), .A3(new_n622), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n650), .A2(new_n651), .A3(new_n652), .A4(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT26), .B1(new_n649), .B2(new_n597), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n622), .A3(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT89), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n567), .A2(new_n517), .A3(new_n569), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n628), .A2(new_n653), .A3(new_n622), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n653), .B1(new_n628), .B2(new_n622), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n659), .A2(new_n662), .A3(new_n513), .A4(new_n598), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(KEYINPUT89), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n658), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n459), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n648), .A2(new_n437), .A3(new_n666), .ZN(G369));
  AND2_X1   g0467(.A1(new_n516), .A2(new_n511), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n512), .B2(new_n486), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n511), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT92), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n668), .A2(new_n675), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n567), .A2(new_n569), .ZN(new_n682));
  INV_X1    g0482(.A(new_n675), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n559), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n570), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n675), .B1(new_n567), .B2(new_n569), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n669), .A2(new_n677), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n668), .A2(new_n683), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n212), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n216), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n530), .A2(new_n532), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n484), .A2(new_n623), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n590), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n568), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n590), .A2(new_n435), .A3(new_n484), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n621), .A2(KEYINPUT93), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n621), .A2(KEYINPUT93), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n708), .A2(new_n536), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n703), .A2(KEYINPUT30), .A3(new_n568), .A4(new_n704), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n675), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR4_X1   g0516(.A1(new_n518), .A2(new_n629), .A3(new_n570), .A4(new_n675), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G330), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n652), .B1(new_n649), .B2(new_n597), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT26), .A4(new_n654), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT94), .B(new_n652), .C1(new_n649), .C2(new_n597), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n663), .A3(new_n622), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(new_n683), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n728), .B1(new_n727), .B2(new_n683), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT29), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n665), .A2(new_n683), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n720), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n701), .B1(new_n736), .B2(G1), .ZN(G364));
  AND2_X1   g0537(.A1(new_n209), .A2(G13), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n208), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n696), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n686), .B2(G330), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G330), .B2(new_n686), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n695), .A2(new_n346), .ZN(new_n744));
  NAND2_X1  g0544(.A1(G355), .A2(KEYINPUT96), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G355), .A2(KEYINPUT96), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(G116), .B2(new_n212), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n248), .A2(new_n257), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n695), .A2(new_n269), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n257), .B2(new_n217), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n218), .B1(G20), .B2(new_n318), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n741), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n209), .A2(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(new_n461), .A3(new_n302), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT99), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT99), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT32), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT98), .ZN(new_n769));
  NAND2_X1  g0569(.A1(G20), .A2(G179), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(new_n302), .ZN(new_n771));
  NAND4_X1  g0571(.A1(KEYINPUT98), .A2(G20), .A3(G179), .A4(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n461), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(new_n461), .A3(new_n772), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G50), .A2(new_n774), .B1(new_n776), .B2(G68), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n761), .A2(new_n461), .A3(G200), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT100), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT100), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n496), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n770), .A2(KEYINPUT97), .ZN(new_n783));
  AOI21_X1  g0583(.A(G200), .B1(new_n770), .B2(KEYINPUT97), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(new_n461), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n782), .B1(G77), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G87), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n461), .A2(G179), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n209), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n790), .B(new_n269), .C1(new_n540), .C2(new_n792), .ZN(new_n793));
  AND3_X1   g0593(.A1(new_n783), .A2(G190), .A3(new_n784), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(G58), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n768), .A2(new_n777), .A3(new_n787), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n781), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n797), .A2(G283), .B1(new_n776), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n346), .B1(new_n788), .B2(new_n800), .C1(new_n792), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n765), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(G329), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n794), .A2(G322), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G311), .A2(new_n786), .B1(new_n774), .B2(G326), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n799), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n796), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n760), .B1(new_n808), .B2(new_n757), .ZN(new_n809));
  INV_X1    g0609(.A(new_n756), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n686), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n743), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  INV_X1    g0613(.A(new_n741), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n443), .A2(new_n675), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n453), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n816), .A2(new_n455), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n455), .A2(new_n675), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n733), .B(new_n819), .Z(new_n820));
  INV_X1    g0620(.A(new_n720), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n814), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n822), .A2(KEYINPUT103), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(KEYINPUT103), .B2(new_n822), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G159), .A2(new_n786), .B1(new_n794), .B2(G143), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G137), .A2(new_n774), .B1(new_n776), .B2(G150), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT34), .Z(new_n828));
  NOR2_X1   g0628(.A1(new_n781), .A2(new_n222), .ZN(new_n829));
  INV_X1    g0629(.A(new_n792), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n346), .B1(new_n830), .B2(G58), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n202), .B2(new_n788), .C1(new_n765), .C2(new_n832), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n828), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n797), .A2(G87), .ZN(new_n835));
  INV_X1    g0635(.A(new_n774), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n800), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G294), .A2(new_n794), .B1(new_n776), .B2(G283), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n544), .B2(new_n785), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n269), .B1(new_n830), .B2(G97), .ZN(new_n840));
  INV_X1    g0640(.A(G311), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n496), .B2(new_n788), .C1(new_n765), .C2(new_n841), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n837), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n757), .B1(new_n834), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n757), .A2(new_n754), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT101), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n844), .B(new_n741), .C1(G77), .C2(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT102), .Z(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n755), .B2(new_n819), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n824), .A2(new_n849), .ZN(G384));
  OR2_X1    g0650(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n851), .A2(G116), .A3(new_n219), .A4(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT36), .Z(new_n854));
  OR3_X1    g0654(.A1(new_n216), .A2(new_n224), .A3(new_n375), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n202), .A2(G68), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n208), .B(G13), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n738), .A2(new_n208), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n819), .B1(new_n716), .B2(new_n717), .ZN(new_n860));
  INV_X1    g0660(.A(new_n304), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n300), .A2(new_n683), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(new_n641), .C2(new_n300), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT104), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n322), .A2(new_n323), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n867), .A2(KEYINPUT104), .A3(new_n861), .A4(new_n863), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n641), .B2(new_n861), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n860), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n394), .A2(new_n430), .ZN(new_n873));
  INV_X1    g0673(.A(new_n366), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n384), .A2(KEYINPUT16), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n420), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n412), .ZN(new_n877));
  INV_X1    g0677(.A(new_n673), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n873), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n673), .B(KEYINPUT105), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n394), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n421), .A2(new_n412), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n873), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n879), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n424), .B2(new_n432), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n887), .B2(new_n889), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT40), .B1(new_n872), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  INV_X1    g0695(.A(new_n432), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n883), .B1(new_n636), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n873), .A2(new_n885), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n394), .A2(new_n882), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT37), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n900), .A2(new_n886), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n895), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n890), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n894), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n893), .B1(new_n872), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n460), .A2(new_n718), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n719), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n890), .A2(new_n891), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n902), .A2(new_n903), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n911), .B1(new_n912), .B2(new_n910), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n867), .A2(new_n675), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT104), .B1(new_n324), .B2(new_n863), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n640), .A2(new_n639), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n300), .B1(new_n917), .B2(new_n315), .ZN(new_n918));
  NOR4_X1   g0718(.A1(new_n918), .A2(new_n865), .A3(new_n304), .A4(new_n862), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n871), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n665), .A2(new_n683), .A3(new_n819), .ZN(new_n921));
  INV_X1    g0721(.A(new_n818), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n923), .A3(new_n892), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n637), .A2(new_n882), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n915), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n732), .A2(new_n735), .A3(new_n459), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n437), .B1(new_n646), .B2(new_n647), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n926), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n859), .B1(new_n909), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n932), .A2(new_n933), .B1(new_n931), .B2(new_n909), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n858), .B1(new_n935), .B2(new_n936), .ZN(G367));
  NOR2_X1   g0737(.A1(new_n240), .A2(new_n751), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n758), .B1(new_n212), .B2(new_n439), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n741), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n269), .B1(new_n830), .B2(G107), .ZN(new_n941));
  INV_X1    g0741(.A(G317), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n765), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT112), .B1(new_n788), .B2(new_n544), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n943), .B1(KEYINPUT46), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n794), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n945), .B1(new_n540), .B2(new_n781), .C1(new_n800), .C2(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n786), .A2(G283), .B1(new_n776), .B2(G294), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n948), .B1(KEYINPUT46), .B2(new_n944), .C1(new_n841), .C2(new_n836), .ZN(new_n949));
  AOI22_X1  g0749(.A1(G50), .A2(new_n786), .B1(new_n794), .B2(G150), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n766), .B2(new_n775), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n792), .A2(new_n222), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n269), .B1(new_n788), .B2(new_n374), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(new_n803), .C2(G137), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n781), .A2(new_n224), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G143), .B2(new_n774), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n947), .A2(new_n949), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT113), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT47), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n940), .B1(new_n960), .B2(new_n757), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n627), .A2(new_n683), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n622), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n662), .B2(new_n963), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n961), .B1(new_n810), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n675), .B1(new_n596), .B2(new_n581), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n593), .A2(new_n597), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT108), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n651), .A2(new_n675), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n693), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(KEYINPUT44), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n693), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  AND4_X1   g0776(.A1(KEYINPUT45), .A2(new_n972), .A3(new_n692), .A4(new_n691), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT45), .B1(new_n693), .B2(new_n972), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n974), .A2(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n688), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n689), .B1(new_n977), .B2(new_n978), .C1(new_n974), .C2(new_n976), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  INV_X1    g0783(.A(new_n690), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n681), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n691), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT111), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n986), .B1(new_n687), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT110), .B1(new_n680), .B2(new_n690), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n687), .A2(new_n987), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n736), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n736), .B1(new_n982), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n696), .B(KEYINPUT41), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n740), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n986), .A2(new_n972), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT42), .Z(new_n999));
  NOR2_X1   g0799(.A1(new_n970), .A2(new_n517), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n651), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n675), .B1(new_n1001), .B2(KEYINPUT109), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT109), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n965), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n688), .A2(new_n972), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1004), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT43), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1006), .B1(new_n1012), .B2(new_n965), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1008), .B(new_n1010), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1009), .B1(new_n1015), .B2(new_n1007), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n967), .B1(new_n997), .B2(new_n1017), .ZN(G387));
  OR3_X1    g0818(.A1(new_n992), .A2(KEYINPUT116), .A3(new_n736), .ZN(new_n1019));
  OAI21_X1  g0819(.A(KEYINPUT116), .B1(new_n992), .B2(new_n736), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1019), .A2(new_n696), .A3(new_n993), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n698), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n744), .A2(new_n1022), .B1(new_n496), .B2(new_n695), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n244), .A2(new_n257), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n364), .A2(new_n202), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n698), .B(new_n257), .C1(new_n222), .C2(new_n224), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n750), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1023), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n814), .B1(new_n1029), .B2(new_n758), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n680), .B2(new_n810), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n836), .A2(new_n766), .B1(new_n326), .B2(new_n775), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G50), .B2(new_n794), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n616), .A2(new_n830), .A3(new_n617), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n269), .B1(new_n788), .B2(new_n224), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n803), .B2(G150), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n797), .A2(G97), .B1(G68), .B2(new_n786), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n830), .A2(G283), .B1(new_n789), .B2(G294), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n774), .A2(G322), .B1(new_n794), .B2(G317), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n800), .B2(new_n785), .C1(new_n841), .C2(new_n775), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT114), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1039), .B1(new_n1044), .B2(KEYINPUT48), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(KEYINPUT48), .B2(new_n1044), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(KEYINPUT115), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n781), .A2(new_n544), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n269), .B(new_n1049), .C1(G326), .C2(new_n803), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1047), .A2(KEYINPUT115), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1038), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1031), .B1(new_n1053), .B2(new_n757), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n740), .B2(new_n992), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1021), .A2(new_n1055), .ZN(G393));
  OAI221_X1 g0856(.A(new_n758), .B1(new_n540), .B2(new_n212), .C1(new_n751), .C2(new_n251), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n741), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n774), .A2(G317), .B1(new_n794), .B2(G311), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT52), .Z(new_n1060));
  INV_X1    g0860(.A(G283), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n346), .B1(new_n788), .B2(new_n1061), .C1(new_n792), .C2(new_n544), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n803), .B2(G322), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n786), .A2(G294), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n782), .B1(G303), .B2(new_n776), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n774), .A2(G150), .B1(new_n794), .B2(G159), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  NAND2_X1  g0868(.A1(new_n803), .A2(G143), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n346), .B1(new_n789), .B2(G68), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1068), .A2(new_n835), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n830), .A2(G77), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n202), .B2(new_n775), .C1(new_n326), .C2(new_n785), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT117), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1066), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT118), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1058), .B1(new_n1076), .B2(new_n757), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n970), .A2(new_n756), .A3(new_n971), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n982), .B2(new_n739), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n982), .A2(new_n993), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1081), .A2(new_n697), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n982), .A2(new_n993), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(G390));
  AOI21_X1  g0885(.A(new_n914), .B1(new_n902), .B2(new_n903), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n727), .A2(new_n683), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT95), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n729), .A3(new_n922), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n817), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n870), .B1(new_n866), .B2(new_n868), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1086), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n914), .B1(new_n920), .B2(new_n923), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n913), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n819), .B(G330), .C1(new_n716), .C2(new_n717), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n860), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n920), .A2(G330), .A3(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1093), .B(new_n1100), .C1(new_n1094), .C2(new_n913), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1102), .A2(new_n739), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n913), .A2(new_n755), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n803), .A2(G294), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1105), .A2(new_n346), .A3(new_n790), .A4(new_n1072), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n829), .B(new_n1106), .C1(G97), .C2(new_n786), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n836), .A2(new_n1061), .B1(new_n496), .B2(new_n775), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G116), .B2(new_n794), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n346), .B1(new_n830), .B2(G159), .ZN(new_n1110));
  INV_X1    g0910(.A(G125), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1110), .B1(new_n781), .B2(new_n202), .C1(new_n1111), .C2(new_n765), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n789), .A2(G150), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT53), .ZN(new_n1114));
  INV_X1    g0914(.A(G128), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n836), .A2(new_n1115), .B1(new_n946), .B2(new_n832), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  AOI22_X1  g0918(.A1(new_n786), .A2(new_n1118), .B1(new_n776), .B2(G137), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT120), .Z(new_n1120));
  AOI22_X1  g0920(.A1(new_n1107), .A2(new_n1109), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n757), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n741), .B1(new_n364), .B2(new_n846), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1104), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1103), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n869), .A2(new_n871), .A3(new_n1096), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT119), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT119), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1092), .A2(new_n1128), .A3(new_n1096), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1127), .A2(new_n1100), .A3(new_n1091), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1126), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n923), .B1(new_n1131), .B2(new_n1097), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n720), .A2(new_n459), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n928), .A2(new_n929), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1102), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1098), .A2(new_n1133), .A3(new_n1101), .A4(new_n1136), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n696), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1125), .A2(new_n1140), .ZN(G378));
  AND3_X1   g0941(.A1(new_n915), .A2(new_n924), .A3(new_n925), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n920), .A2(new_n892), .A3(new_n1099), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n894), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n719), .B1(new_n872), .B2(new_n904), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n335), .A2(new_n673), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n647), .A2(new_n436), .A3(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n335), .B(new_n673), .C1(new_n363), .C2(new_n437), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OR3_X1    g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1144), .A2(new_n1145), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1142), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT122), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n872), .A2(new_n904), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(G330), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1160), .B2(new_n893), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1144), .A2(new_n1145), .A3(new_n1153), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n926), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1156), .A2(new_n1157), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1139), .A2(new_n1136), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1142), .B(KEYINPUT122), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1139), .B2(new_n1136), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1156), .A2(new_n1163), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n697), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1164), .A2(new_n740), .A3(new_n1166), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n846), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n814), .B1(new_n1175), .B2(new_n202), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G137), .A2(new_n786), .B1(new_n794), .B2(G128), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n1111), .B2(new_n836), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n830), .A2(G150), .B1(new_n789), .B2(new_n1118), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n832), .B2(new_n775), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n797), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n803), .C2(G124), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n346), .A2(new_n256), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1188), .B(new_n952), .C1(G77), .C2(new_n789), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n1061), .B2(new_n765), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n797), .A2(G58), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n544), .B2(new_n836), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n786), .A2(new_n616), .A3(new_n617), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n540), .B2(new_n775), .C1(new_n496), .C2(new_n946), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1190), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1195), .A2(KEYINPUT58), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(KEYINPUT58), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1188), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1198));
  AND4_X1   g0998(.A1(new_n1187), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1176), .B1(new_n1122), .B2(new_n1199), .C1(new_n1158), .C2(new_n755), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT121), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1174), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1173), .A2(new_n1204), .ZN(G375));
  XNOR2_X1  g1005(.A(new_n739), .B(KEYINPUT123), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1133), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n814), .B1(new_n1175), .B2(new_n222), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n946), .A2(new_n1061), .B1(new_n496), .B2(new_n785), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G116), .B2(new_n776), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n269), .B1(new_n789), .B2(G97), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1034), .B(new_n1212), .C1(new_n765), .C2(new_n800), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n955), .B(new_n1213), .C1(G294), .C2(new_n774), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n346), .B1(new_n789), .B2(G159), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1191), .B(new_n1215), .C1(new_n1115), .C2(new_n765), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G137), .A2(new_n794), .B1(new_n776), .B2(new_n1118), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n832), .B2(new_n836), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n785), .A2(new_n327), .B1(new_n792), .B2(new_n202), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT124), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1211), .A2(new_n1214), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1209), .B1(new_n1122), .B2(new_n1222), .C1(new_n920), .C2(new_n755), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1208), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n648), .A2(new_n437), .A3(new_n927), .A4(new_n1134), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1132), .A3(new_n1130), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1137), .A2(new_n996), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(G381));
  AOI21_X1  g1029(.A(new_n1203), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1230));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(G390), .A2(G387), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1021), .A2(new_n812), .A3(new_n1055), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(G381), .A2(G384), .A3(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1234), .ZN(G407));
  INV_X1    g1035(.A(G213), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(G343), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1230), .A2(new_n1231), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238), .ZN(G409));
  INV_X1    g1039(.A(KEYINPUT126), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1233), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n812), .B1(new_n1021), .B2(new_n1055), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G390), .A2(G387), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1240), .B(new_n1243), .C1(new_n1245), .C2(new_n1232), .ZN(new_n1246));
  OR2_X1    g1046(.A1(G390), .A2(G387), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1242), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1240), .A3(new_n1233), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT126), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1247), .A2(new_n1249), .A3(new_n1244), .A4(new_n1250), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1246), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1173), .A2(G378), .A3(new_n1204), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1164), .A2(new_n1165), .A3(new_n996), .A4(new_n1166), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1201), .B1(new_n1171), .B2(new_n1207), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1231), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1237), .B1(new_n1254), .B2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1226), .A2(new_n1130), .A3(KEYINPUT60), .A4(new_n1132), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n696), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1137), .A2(KEYINPUT60), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n1227), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n824), .B(new_n849), .C1(new_n1263), .C2(new_n1224), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1262), .A2(new_n1227), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G384), .B(new_n1225), .C1(new_n1265), .C2(new_n1261), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1237), .A2(G2897), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1264), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1252), .B(new_n1253), .C1(new_n1259), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1237), .B(new_n1267), .C1(new_n1254), .C2(new_n1258), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(KEYINPUT63), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1237), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1267), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(KEYINPUT125), .A3(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1274), .A2(new_n1277), .A3(new_n1278), .A4(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1252), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1264), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1268), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G378), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1230), .B2(G378), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1289), .B1(new_n1291), .B2(new_n1237), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1279), .A2(new_n1293), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(new_n1294), .A3(new_n1253), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1276), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1286), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1285), .A2(new_n1298), .ZN(G405));
  XNOR2_X1  g1099(.A(new_n1230), .B(new_n1231), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1267), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1300), .A2(new_n1267), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1286), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1303), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n1252), .A3(new_n1301), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(G402));
endmodule


