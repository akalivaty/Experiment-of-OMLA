//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n192), .B1(new_n189), .B2(new_n191), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n187), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT67), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(new_n191), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(new_n187), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(new_n187), .C1(new_n193), .C2(new_n194), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT30), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n204), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n204), .B(KEYINPUT1), .C1(new_n208), .C2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G128), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT64), .A2(G143), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT64), .A2(G143), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n211), .A2(new_n212), .A3(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n205), .A2(G143), .ZN(new_n214));
  OAI22_X1  g028(.A1(new_n207), .A2(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(G146), .B1(new_n211), .B2(new_n212), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n206), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G134), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G137), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n221), .A2(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT11), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n221), .B2(G137), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT11), .A3(G134), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .A4(new_n222), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT68), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n225), .A2(new_n234), .A3(new_n231), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n220), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n227), .A2(new_n222), .A3(new_n229), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n231), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n208), .A2(G146), .ZN(new_n240));
  OR2_X1    g054(.A1(KEYINPUT64), .A2(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT64), .A2(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n243), .B2(G146), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT0), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(new_n217), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n246), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n248), .B(new_n250), .C1(new_n213), .C2(new_n214), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n239), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n203), .B1(new_n236), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n232), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n209), .A2(G128), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT65), .B1(new_n240), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n241), .A2(new_n205), .A3(new_n242), .ZN(new_n258));
  INV_X1    g072(.A(new_n214), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n255), .A2(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n219), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n254), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n262), .A2(new_n203), .A3(new_n252), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n202), .B1(new_n253), .B2(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n225), .A2(new_n234), .A3(new_n231), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n234), .B1(new_n225), .B2(new_n231), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI211_X1 g081(.A(new_n246), .B(new_n249), .C1(new_n258), .C2(new_n259), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n216), .A2(new_n206), .A3(new_n246), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n267), .A2(new_n220), .B1(new_n270), .B2(new_n239), .ZN(new_n271));
  INV_X1    g085(.A(new_n202), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT26), .B(G101), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT69), .B(G953), .ZN(new_n277));
  INV_X1    g091(.A(G237), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(G210), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n276), .B(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n264), .A2(new_n273), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT31), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n264), .A2(new_n284), .A3(new_n273), .A4(new_n281), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n236), .A2(new_n252), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n202), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n271), .A2(KEYINPUT28), .A3(new_n272), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n262), .A2(new_n252), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n202), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n280), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n283), .A2(new_n285), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n294), .B2(new_n296), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n287), .A2(new_n202), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n288), .A2(new_n289), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n281), .A2(KEYINPUT29), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n288), .A2(new_n289), .A3(new_n281), .A4(new_n291), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n264), .A2(new_n273), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n309), .B2(new_n280), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n305), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G472), .ZN(new_n312));
  OAI22_X1  g126(.A1(new_n298), .A2(new_n299), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n314));
  XNOR2_X1  g128(.A(G119), .B(G128), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(KEYINPUT23), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n318), .A2(new_n320), .A3(G119), .A4(new_n217), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT24), .B(G110), .Z(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n315), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n322), .A2(G110), .B1(KEYINPUT72), .B2(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n324), .A2(KEYINPUT72), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT16), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT74), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT16), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n327), .A3(G125), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT75), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n337), .A2(G146), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(G146), .B1(new_n337), .B2(new_n339), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n325), .B(new_n326), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  OAI22_X1  g156(.A1(new_n322), .A2(G110), .B1(new_n315), .B2(new_n323), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n337), .A2(G146), .A3(new_n339), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n334), .A2(new_n205), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT76), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT77), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n342), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G137), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n354), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n342), .A2(new_n350), .A3(new_n347), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n314), .B1(new_n358), .B2(new_n304), .ZN(new_n359));
  AOI211_X1 g173(.A(KEYINPUT25), .B(G902), .C1(new_n355), .C2(new_n357), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G217), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(G234), .B2(new_n304), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G902), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n361), .A2(new_n363), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n313), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G122), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G116), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(G116), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT14), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT94), .B(KEYINPUT14), .C1(new_n368), .C2(G116), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT95), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n377), .A2(KEYINPUT95), .A3(new_n371), .A4(new_n378), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n381), .B(new_n382), .C1(KEYINPUT14), .C2(new_n370), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G107), .ZN(new_n384));
  OAI21_X1  g198(.A(G128), .B1(new_n211), .B2(new_n212), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT92), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n387), .B(G128), .C1(new_n211), .C2(new_n212), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n208), .A2(G128), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT93), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT93), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n393), .B(new_n390), .C1(new_n386), .C2(new_n388), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n392), .A2(new_n394), .A3(new_n221), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n387), .B1(new_n243), .B2(G128), .ZN(new_n396));
  INV_X1    g210(.A(new_n388), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n391), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n393), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n389), .A2(KEYINPUT93), .A3(new_n391), .ZN(new_n400));
  AOI21_X1  g214(.A(G134), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n374), .B(new_n384), .C1(new_n395), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT13), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n390), .B1(new_n389), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n403), .B2(new_n389), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G134), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n221), .B1(new_n392), .B2(new_n394), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n372), .B(new_n373), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT9), .B(G234), .Z(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n411), .A2(new_n362), .A3(G953), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n402), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n402), .B2(new_n409), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n304), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT96), .ZN(new_n416));
  INV_X1    g230(.A(G478), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT15), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT96), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n419), .B(new_n304), .C1(new_n413), .C2(new_n414), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT97), .B1(new_n415), .B2(new_n418), .ZN(new_n422));
  INV_X1    g236(.A(new_n415), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n424));
  INV_X1    g238(.A(new_n418), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n421), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(KEYINPUT69), .A2(G953), .ZN(new_n428));
  NOR2_X1   g242(.A1(KEYINPUT69), .A2(G953), .ZN(new_n429));
  OAI211_X1 g243(.A(G214), .B(new_n278), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n211), .A2(new_n212), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n277), .A2(new_n208), .A3(G214), .A4(new_n278), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n230), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n433), .A3(G131), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT91), .B1(new_n437), .B2(KEYINPUT17), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n340), .A2(new_n341), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT17), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n435), .A2(new_n442), .A3(new_n440), .A4(new_n436), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n438), .A2(new_n439), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n346), .B1(new_n205), .B2(new_n334), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT18), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n434), .B1(new_n446), .B2(new_n230), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n445), .B(new_n447), .C1(new_n446), .C2(new_n436), .ZN(new_n448));
  XNOR2_X1  g262(.A(G113), .B(G122), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT89), .B(G104), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT90), .Z(new_n452));
  NAND3_X1  g266(.A1(new_n444), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(new_n444), .B2(new_n448), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n304), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G475), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n334), .B(KEYINPUT19), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n205), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n437), .A2(new_n344), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n448), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n451), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(G475), .B1(new_n453), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n465), .A3(new_n304), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n465), .B1(new_n464), .B2(new_n304), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n457), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G952), .ZN(new_n471));
  AOI211_X1 g285(.A(G953), .B(new_n471), .C1(G234), .C2(G237), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI211_X1 g287(.A(new_n304), .B(new_n277), .C1(G234), .C2(G237), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT21), .B(G898), .Z(new_n476));
  OAI21_X1  g290(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n427), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G214), .B1(G237), .B2(G902), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(G110), .B(G122), .Z(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT8), .ZN(new_n482));
  OR2_X1    g296(.A1(KEYINPUT78), .A2(G104), .ZN(new_n483));
  NAND2_X1  g297(.A1(KEYINPUT78), .A2(G104), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n373), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT3), .ZN(new_n486));
  INV_X1    g300(.A(G101), .ZN(new_n487));
  AND2_X1   g301(.A1(KEYINPUT78), .A2(G104), .ZN(new_n488));
  NOR2_X1   g302(.A1(KEYINPUT78), .A2(G104), .ZN(new_n489));
  OAI21_X1  g303(.A(G107), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G104), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n491), .A2(KEYINPUT3), .A3(G107), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n486), .A2(new_n487), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  OR3_X1    g308(.A1(new_n373), .A2(KEYINPUT80), .A3(G104), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT80), .B1(new_n373), .B2(G104), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G101), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n193), .A2(new_n194), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT85), .B(KEYINPUT5), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n189), .ZN(new_n503));
  INV_X1    g317(.A(G113), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n499), .B1(new_n507), .B2(new_n198), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n499), .A2(new_n198), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n505), .B1(new_n510), .B2(new_n197), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n482), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G224), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(G953), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT86), .ZN(new_n516));
  OAI21_X1  g330(.A(G125), .B1(new_n268), .B2(new_n269), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n215), .A2(new_n329), .A3(new_n219), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n329), .B1(new_n247), .B2(new_n251), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT86), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n515), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n215), .A2(new_n329), .A3(new_n219), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT86), .B1(new_n523), .B2(new_n520), .ZN(new_n524));
  INV_X1    g338(.A(new_n515), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n517), .A2(new_n516), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n513), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n488), .A2(new_n489), .A3(G107), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT3), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n490), .B(new_n493), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G101), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT79), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n492), .B1(new_n485), .B2(KEYINPUT3), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n487), .B1(new_n538), .B2(new_n490), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT4), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND4_X1   g355(.A1(new_n537), .A2(new_n534), .A3(new_n540), .A4(G101), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n202), .B(new_n536), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n481), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n509), .A2(new_n506), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n529), .B1(new_n519), .B2(new_n521), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(G902), .B1(new_n531), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n545), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n481), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(KEYINPUT6), .A3(new_n546), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT6), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n553), .A3(new_n481), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n554), .A3(new_n528), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT88), .ZN(new_n557));
  OAI21_X1  g371(.A(G210), .B1(G237), .B2(G902), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT87), .Z(new_n559));
  AND3_X1   g373(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n557), .B1(new_n556), .B2(new_n559), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n549), .A2(new_n555), .A3(new_n558), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n480), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT84), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n257), .A2(G128), .A3(new_n209), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n258), .A2(new_n259), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n567), .A2(new_n568), .B1(new_n244), .B2(new_n218), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n499), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n217), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n219), .B1(new_n571), .B2(new_n244), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n494), .A3(new_n498), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT81), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n239), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n574), .B2(new_n239), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n566), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n270), .B(new_n536), .C1(new_n541), .C2(new_n542), .ZN(new_n580));
  INV_X1    g394(.A(new_n239), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT10), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n494), .A4(new_n498), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n580), .A2(new_n581), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n277), .A2(G227), .ZN(new_n586));
  XNOR2_X1  g400(.A(G110), .B(G140), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n570), .A2(new_n573), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT81), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n239), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT12), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(KEYINPUT84), .A3(new_n576), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n579), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n239), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n585), .ZN(new_n598));
  INV_X1    g412(.A(new_n588), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G469), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n304), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n585), .A2(new_n593), .A3(new_n576), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT82), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n585), .A2(new_n593), .A3(KEYINPUT82), .A4(new_n576), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n599), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n585), .A2(new_n588), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT83), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n585), .A2(KEYINPUT83), .A3(new_n588), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n597), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n608), .A2(G469), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(G469), .A2(G902), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n603), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G221), .B1(new_n411), .B2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n367), .A2(new_n478), .A3(new_n565), .A4(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT98), .B(G101), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT99), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n620), .B(new_n622), .ZN(G3));
  AOI21_X1  g437(.A(new_n558), .B1(new_n549), .B2(new_n555), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n479), .B1(new_n563), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT100), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n627), .B(new_n479), .C1(new_n563), .C2(new_n624), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n477), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n402), .A2(new_n409), .A3(new_n412), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n402), .A2(new_n409), .ZN(new_n635));
  INV_X1    g449(.A(new_n412), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n402), .A2(new_n409), .A3(KEYINPUT102), .A4(new_n412), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n634), .A2(new_n637), .A3(KEYINPUT33), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT101), .B(KEYINPUT33), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n413), .B2(new_n414), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n417), .A2(G902), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n631), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n639), .A2(KEYINPUT103), .A3(new_n643), .A4(new_n641), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n469), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n294), .A2(new_n304), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n651), .A2(G472), .B1(new_n296), .B2(new_n294), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n365), .A2(new_n616), .A3(new_n617), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n630), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n491), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT104), .B(KEYINPUT34), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  AOI22_X1  g471(.A1(new_n468), .A2(KEYINPUT105), .B1(new_n456), .B2(G475), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n453), .A2(new_n463), .ZN(new_n659));
  INV_X1    g473(.A(G475), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n304), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT20), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n466), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n427), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n630), .A2(new_n653), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  INV_X1    g483(.A(new_n359), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n358), .A2(new_n314), .A3(new_n304), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n363), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n356), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n348), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n364), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n652), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n478), .A2(new_n565), .A3(new_n678), .A4(new_n619), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  NAND2_X1  g495(.A1(new_n672), .A2(new_n675), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n626), .A2(new_n628), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n313), .A2(new_n617), .A3(new_n616), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n658), .A2(new_n664), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n421), .A2(new_n422), .A3(new_n426), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n473), .B1(new_n475), .B2(G900), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n683), .A2(new_n685), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  NAND2_X1  g506(.A1(new_n562), .A2(new_n564), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT38), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n562), .A2(KEYINPUT38), .A3(new_n564), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n309), .A2(new_n281), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n273), .A2(new_n300), .A3(new_n280), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n699), .A2(new_n304), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n312), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n294), .A2(new_n296), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT32), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n701), .B1(new_n703), .B2(new_n297), .ZN(new_n704));
  OR4_X1    g518(.A1(new_n427), .A2(new_n704), .A3(new_n470), .A4(new_n480), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n688), .B(KEYINPUT39), .Z(new_n708));
  OAI21_X1  g522(.A(new_n707), .B1(new_n618), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n618), .A2(new_n707), .A3(new_n708), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT40), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n711), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n709), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n706), .A2(new_n712), .A3(new_n715), .A4(new_n676), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n431), .ZN(G45));
  AND3_X1   g531(.A1(new_n648), .A2(new_n469), .A3(new_n688), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n683), .A2(new_n685), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT107), .B(G146), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G48));
  AOI21_X1  g535(.A(new_n602), .B1(new_n601), .B2(new_n304), .ZN(new_n722));
  AOI211_X1 g536(.A(G469), .B(G902), .C1(new_n595), .C2(new_n600), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n313), .A2(new_n724), .A3(new_n365), .A4(new_n617), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n629), .A2(new_n725), .A3(new_n649), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT41), .B(G113), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n666), .A2(new_n477), .A3(new_n628), .A4(new_n626), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT108), .B1(new_n729), .B2(new_n725), .ZN(new_n730));
  INV_X1    g544(.A(new_n725), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n630), .A2(new_n731), .A3(new_n732), .A4(new_n666), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  INV_X1    g549(.A(new_n722), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n617), .A3(new_n603), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n683), .A2(new_n313), .A3(new_n478), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  AND2_X1   g554(.A1(new_n687), .A2(new_n469), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n477), .A3(new_n628), .A4(new_n626), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n358), .A2(new_n364), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n672), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n651), .A2(G472), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n301), .A2(new_n280), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n283), .A2(new_n285), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n296), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n738), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n368), .ZN(G24));
  INV_X1    g567(.A(new_n749), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n683), .A2(new_n718), .A3(new_n738), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  INV_X1    g570(.A(new_n561), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n479), .A3(new_n564), .A4(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n688), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n649), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n614), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n608), .A2(KEYINPUT109), .A3(G469), .A4(new_n613), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n603), .A3(new_n615), .A4(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(new_n617), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n761), .A2(new_n367), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n703), .A2(new_n297), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT110), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n308), .A2(new_n310), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n304), .A3(new_n303), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(G472), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n744), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(KEYINPUT42), .A3(new_n761), .A4(new_n766), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n769), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  INV_X1    g592(.A(new_n759), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n766), .A2(new_n690), .A3(new_n367), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  NOR3_X1   g595(.A1(new_n676), .A2(KEYINPUT111), .A3(new_n652), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n682), .B2(new_n677), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n648), .A2(KEYINPUT43), .A3(new_n470), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT43), .B1(new_n648), .B2(new_n470), .ZN(new_n786));
  OAI22_X1  g600(.A1(new_n782), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n787), .A2(new_n790), .A3(new_n788), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n779), .B(new_n789), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n608), .A2(new_n613), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n608), .A2(KEYINPUT45), .A3(new_n613), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(G469), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n615), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n615), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n603), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n617), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(new_n708), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n793), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n228), .ZN(G39));
  NOR2_X1   g621(.A1(new_n313), .A2(new_n365), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n803), .A2(KEYINPUT47), .A3(new_n617), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT47), .B1(new_n803), .B2(new_n617), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n761), .B(new_n808), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(new_n724), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n744), .B(new_n480), .C1(new_n814), .C2(KEYINPUT49), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n470), .A3(new_n617), .A4(new_n648), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT113), .Z(new_n817));
  OR2_X1    g631(.A1(new_n814), .A2(KEYINPUT49), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n697), .A3(new_n704), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n470), .A2(new_n687), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n649), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n653), .A3(new_n565), .A4(new_n477), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n780), .A2(new_n822), .A3(new_n620), .A4(new_n679), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n765), .A2(new_n617), .A3(new_n754), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n686), .A2(new_n427), .ZN(new_n825));
  OAI22_X1  g639(.A1(new_n824), .A2(new_n649), .B1(new_n684), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n676), .A2(new_n760), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n826), .A2(new_n779), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n683), .B(new_n685), .C1(new_n690), .C2(new_n718), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n626), .A2(new_n628), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n704), .A2(new_n682), .A3(new_n760), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n766), .A3(new_n741), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n755), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n755), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n829), .A2(KEYINPUT114), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n837), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n822), .A2(new_n620), .A3(new_n679), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n826), .A2(new_n779), .A3(new_n827), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n780), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n752), .A2(new_n726), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n734), .A2(new_n844), .A3(new_n739), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n840), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n839), .A2(new_n846), .A3(new_n777), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n734), .A2(new_n739), .A3(new_n844), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n829), .A3(new_n835), .A4(new_n837), .ZN(new_n849));
  INV_X1    g663(.A(new_n777), .ZN(new_n850));
  OAI211_X1 g664(.A(KEYINPUT53), .B(new_n838), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT54), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT47), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n804), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n854), .B(new_n809), .C1(new_n617), .C2(new_n814), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n785), .A2(new_n786), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n473), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n750), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n779), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n779), .A2(new_n682), .A3(new_n738), .A4(new_n754), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n724), .A2(new_n480), .A3(new_n617), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n697), .A3(new_n750), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n861), .B1(new_n865), .B2(KEYINPUT50), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n857), .A2(new_n697), .A3(new_n750), .A4(new_n864), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n866), .A2(new_n857), .B1(KEYINPUT50), .B2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n759), .A2(new_n737), .A3(new_n744), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n472), .A3(new_n704), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n870), .B(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n648), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n470), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n860), .A2(new_n868), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n872), .A2(new_n650), .ZN(new_n878));
  INV_X1    g692(.A(G953), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n771), .A2(new_n774), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n857), .A2(new_n880), .A3(new_n869), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT48), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(KEYINPUT118), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n878), .A2(G952), .A3(new_n879), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT48), .B1(new_n881), .B2(KEYINPUT118), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(KEYINPUT118), .B2(new_n881), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n860), .A2(new_n868), .A3(KEYINPUT51), .A4(new_n874), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n877), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n840), .A2(new_n843), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(KEYINPUT53), .A3(new_n777), .A4(new_n848), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n849), .B2(new_n850), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n857), .A2(new_n831), .A3(new_n738), .A4(new_n750), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT117), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n852), .A2(new_n889), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n819), .B1(new_n898), .B2(new_n899), .ZN(G75));
  NAND2_X1  g714(.A1(new_n552), .A2(new_n554), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT119), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n528), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n847), .A2(new_n851), .A3(G902), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n559), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n847), .A2(new_n851), .A3(G210), .A4(G902), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n909), .B2(new_n905), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n277), .A2(G952), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(G51));
  XOR2_X1   g726(.A(new_n615), .B(KEYINPUT57), .Z(new_n913));
  AND3_X1   g727(.A1(new_n847), .A2(new_n851), .A3(KEYINPUT54), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n852), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n601), .ZN(new_n916));
  INV_X1    g730(.A(new_n798), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n911), .B1(new_n916), .B2(new_n918), .ZN(G54));
  AND2_X1   g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n847), .A2(new_n851), .A3(G902), .A4(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n659), .ZN(new_n922));
  OR3_X1    g736(.A1(new_n921), .A2(KEYINPUT120), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n911), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT120), .B1(new_n921), .B2(new_n922), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G60));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT59), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n852), .B2(new_n895), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n642), .ZN(new_n931));
  INV_X1    g745(.A(new_n911), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n642), .A2(new_n928), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n914), .B2(new_n852), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT60), .Z(new_n937));
  NAND3_X1  g751(.A1(new_n847), .A2(new_n851), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n357), .A3(new_n355), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n847), .A2(new_n851), .A3(new_n674), .A4(new_n937), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n932), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(KEYINPUT61), .A3(new_n932), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(G66));
  AOI21_X1  g759(.A(new_n879), .B1(new_n476), .B2(G224), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n848), .A2(new_n841), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n277), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n902), .B1(G898), .B2(new_n277), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT121), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  NOR2_X1   g765(.A1(new_n710), .A2(new_n711), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(new_n367), .A3(new_n779), .A4(new_n821), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n793), .B2(new_n805), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n830), .A2(new_n755), .ZN(new_n956));
  XNOR2_X1  g770(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n716), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n812), .ZN(new_n959));
  NOR2_X1   g773(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n716), .B2(new_n956), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n963), .B(new_n953), .C1(new_n793), .C2(new_n805), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n955), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n253), .A2(new_n263), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n458), .B(KEYINPUT122), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n277), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n968), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n277), .A2(G227), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n775), .A2(new_n831), .A3(new_n741), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n805), .B1(new_n793), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n812), .A2(new_n780), .A3(new_n956), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n850), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n277), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n970), .B(new_n971), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(G900), .B1(new_n970), .B2(G227), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n976), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n969), .A2(new_n977), .A3(new_n979), .ZN(G72));
  INV_X1    g794(.A(new_n947), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n955), .A2(new_n981), .A3(new_n962), .A4(new_n964), .ZN(new_n982));
  XNOR2_X1  g796(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n312), .A2(new_n304), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n983), .B(new_n984), .Z(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n982), .A2(KEYINPUT126), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(KEYINPUT126), .B1(new_n982), .B2(new_n986), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n987), .A2(new_n988), .A3(new_n698), .ZN(new_n989));
  INV_X1    g803(.A(new_n309), .ZN(new_n990));
  NOR4_X1   g804(.A1(new_n973), .A2(new_n974), .A3(new_n947), .A4(new_n850), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n990), .B(new_n280), .C1(new_n991), .C2(new_n985), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n892), .A2(new_n894), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n282), .A2(KEYINPUT127), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n309), .A2(new_n280), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n993), .A2(new_n986), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n992), .A2(new_n997), .A3(new_n932), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n989), .A2(new_n998), .ZN(G57));
endmodule


