//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(new_n204), .B2(new_n205), .ZN(new_n207));
  NOR2_X1   g006(.A1(G127gat), .A2(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G134gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT68), .B(G127gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n207), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G113gat), .B2(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G127gat), .A2(G134gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT69), .B(G113gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G120gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G141gat), .B(G148gat), .Z(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n222), .A2(new_n226), .B1(new_n223), .B2(KEYINPUT77), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n222), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(new_n225), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n221), .B(new_n223), .C1(new_n230), .C2(KEYINPUT77), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n220), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n233), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n203), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n212), .A2(KEYINPUT70), .A3(new_n219), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT70), .B1(new_n212), .B2(new_n219), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n238), .B1(new_n241), .B2(new_n232), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT68), .B(G127gat), .Z(new_n243));
  AOI21_X1  g042(.A(new_n208), .B1(new_n243), .B2(G134gat), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n244), .A2(new_n207), .B1(new_n218), .B2(new_n216), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(new_n232), .A3(new_n238), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT78), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n245), .A2(new_n232), .A3(new_n248), .A4(new_n238), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n237), .B1(new_n242), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n252));
  INV_X1    g051(.A(new_n232), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n220), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(new_n232), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n252), .B1(new_n256), .B2(new_n203), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(KEYINPUT4), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT80), .ZN(new_n259));
  INV_X1    g058(.A(new_n240), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT70), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n238), .A4(new_n232), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT80), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n255), .A2(new_n263), .A3(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n236), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n202), .B(new_n252), .C1(new_n266), .C2(new_n234), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n251), .A2(new_n257), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G1gat), .B(G29gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT0), .ZN(new_n271));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  AOI21_X1  g072(.A(KEYINPUT6), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT81), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n273), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n251), .A2(new_n257), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n265), .A2(new_n268), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n274), .B2(new_n275), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT82), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n269), .A2(new_n273), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT81), .B1(new_n284), .B2(KEYINPUT6), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n276), .A4(new_n281), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n269), .A2(new_n273), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT6), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G8gat), .B(G36gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G64gat), .B(G92gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT64), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT24), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT24), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G169gat), .ZN(new_n308));
  INV_X1    g107(.A(G176gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  XOR2_X1   g111(.A(KEYINPUT65), .B(G176gat), .Z(new_n313));
  NOR2_X1   g112(.A1(new_n311), .A2(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n296), .B1(new_n305), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n303), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(G183gat), .B2(G190gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n296), .B1(new_n314), .B2(new_n309), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n319), .A2(KEYINPUT66), .A3(new_n312), .A4(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n312), .B(new_n320), .C1(new_n304), .C2(new_n297), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT27), .B(G183gat), .ZN(new_n326));
  INV_X1    g125(.A(G190gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n310), .B1(KEYINPUT26), .B2(new_n307), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT26), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT67), .B1(new_n306), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n306), .A2(KEYINPUT67), .A3(new_n332), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(new_n300), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n295), .B1(new_n325), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G226gat), .ZN(new_n339));
  INV_X1    g138(.A(G233gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n295), .A3(new_n336), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT74), .ZN(new_n345));
  XNOR2_X1  g144(.A(G197gat), .B(G204gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT22), .ZN(new_n347));
  INV_X1    g146(.A(G211gat), .ZN(new_n348));
  INV_X1    g147(.A(G218gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n344), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n351), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n356), .A3(KEYINPUT75), .ZN(new_n357));
  OR3_X1    g156(.A1(new_n354), .A2(KEYINPUT75), .A3(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n325), .A2(new_n336), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n341), .A2(KEYINPUT29), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n343), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n325), .A2(new_n295), .A3(new_n336), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n364), .B2(new_n337), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n325), .A2(new_n336), .A3(new_n341), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n359), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n294), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n366), .ZN(new_n369));
  INV_X1    g168(.A(new_n359), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n343), .A2(new_n359), .A3(new_n362), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n293), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(new_n373), .A3(KEYINPUT30), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n363), .A2(new_n367), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n293), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n290), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n358), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n232), .B1(new_n381), .B2(new_n233), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G228gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(new_n340), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n236), .A2(new_n380), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n359), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(KEYINPUT83), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n390));
  INV_X1    g189(.A(new_n388), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(new_n382), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n359), .A2(new_n387), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n352), .B2(new_n356), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n253), .B1(new_n395), .B2(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n386), .ZN(new_n398));
  XNOR2_X1  g197(.A(G78gat), .B(G106gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT31), .B(G50gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G22gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(new_n401), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n393), .A2(new_n398), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n393), .B2(new_n398), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n371), .A2(new_n372), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n343), .A2(new_n370), .A3(new_n362), .ZN(new_n413));
  INV_X1    g212(.A(new_n366), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n338), .A2(new_n342), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(new_n361), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n413), .B(KEYINPUT37), .C1(new_n416), .C2(new_n370), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT38), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n412), .A2(new_n417), .A3(new_n418), .A4(new_n294), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n274), .A2(new_n281), .ZN(new_n420));
  AND4_X1   g219(.A1(new_n289), .A2(new_n419), .A3(new_n373), .A4(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n412), .B(new_n294), .C1(new_n375), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT38), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n410), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT39), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n235), .A2(new_n236), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n265), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT85), .B1(new_n428), .B2(new_n203), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT85), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n430), .B(new_n202), .C1(new_n265), .C2(new_n427), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n426), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n203), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n430), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(KEYINPUT85), .A3(new_n203), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT39), .B1(new_n256), .B2(new_n203), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n432), .B(new_n273), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT40), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n378), .A2(new_n288), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT40), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n379), .A2(new_n410), .B1(new_n425), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G15gat), .B(G43gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n260), .A2(new_n261), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n360), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n241), .A2(new_n336), .A3(new_n325), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G227gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(new_n340), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT71), .ZN(new_n460));
  INV_X1    g259(.A(new_n455), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n451), .B2(new_n452), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT32), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n456), .B(KEYINPUT32), .C1(new_n457), .C2(new_n449), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n461), .A3(new_n452), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n468), .B(KEYINPUT34), .Z(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT73), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n465), .B2(new_n466), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT73), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n471), .A2(KEYINPUT36), .A3(new_n473), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n446), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n473), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n410), .A2(new_n482), .A3(new_n475), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n290), .A3(new_n378), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT35), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n420), .A2(new_n289), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n378), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n476), .B2(new_n474), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G197gat), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT11), .B(G169gat), .Z(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n496), .B(KEYINPUT12), .Z(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  AND2_X1   g297(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G29gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n501), .A2(new_n503), .B1(new_n504), .B2(KEYINPUT15), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT15), .ZN(new_n506));
  INV_X1    g305(.A(G43gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n508));
  INV_X1    g307(.A(G50gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G43gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n506), .B(new_n508), .C1(new_n512), .C2(KEYINPUT89), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n505), .A2(new_n513), .A3(KEYINPUT90), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n501), .A2(KEYINPUT15), .A3(new_n504), .A4(new_n503), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT90), .B1(new_n505), .B2(new_n513), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT17), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n505), .A2(new_n513), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT17), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n521), .A2(new_n522), .A3(new_n515), .A4(new_n514), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n402), .A2(G15gat), .ZN(new_n525));
  INV_X1    g324(.A(G15gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT16), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT92), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n529), .ZN(new_n534));
  INV_X1    g333(.A(G8gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n532), .ZN(new_n538));
  NAND2_X1  g337(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n528), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n530), .A2(KEYINPUT91), .A3(G8gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n532), .A2(G1gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT93), .B1(new_n537), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n541), .A2(new_n542), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n536), .A3(new_n546), .A4(new_n540), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n524), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n516), .A2(new_n517), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n536), .A3(new_n540), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n551), .B(new_n552), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n550), .B(KEYINPUT13), .Z(new_n557));
  AOI22_X1  g356(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n549), .A2(KEYINPUT18), .A3(new_n550), .A4(new_n553), .ZN(new_n559));
  AOI211_X1 g358(.A(KEYINPUT88), .B(new_n497), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n497), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(new_n555), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n557), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT88), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n492), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G57gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G64gat), .ZN(new_n575));
  INV_X1    g374(.A(G64gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G57gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT95), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n573), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n569), .A2(KEYINPUT94), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n569), .A2(KEYINPUT94), .ZN(new_n583));
  NOR2_X1   g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT96), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n581), .A2(new_n585), .A3(KEYINPUT96), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n584), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n569), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT97), .B1(new_n581), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n575), .A2(new_n577), .B1(new_n579), .B2(KEYINPUT95), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n573), .A4(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G127gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n552), .B1(new_n599), .B2(new_n600), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  INV_X1    g406(.A(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G183gat), .B(G211gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n606), .B(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G85gat), .A2(G92gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT99), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(KEYINPUT99), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(G85gat), .A3(G92gat), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n619), .A3(KEYINPUT7), .ZN(new_n620));
  NAND2_X1  g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT8), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n623));
  OR2_X1    g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n622), .B2(new_n624), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n616), .B(new_n620), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G99gat), .B(G106gat), .Z(new_n628));
  OAI21_X1  g427(.A(KEYINPUT101), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n622), .A2(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT100), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n622), .A2(new_n624), .A3(new_n623), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n620), .A2(new_n616), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635));
  INV_X1    g434(.A(new_n628), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n629), .A2(new_n637), .B1(new_n628), .B2(new_n627), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n524), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G190gat), .B(G218gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT102), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n643));
  NAND2_X1  g442(.A1(G232gat), .A2(G233gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n551), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(new_n646), .B2(new_n638), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n641), .A2(KEYINPUT102), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(new_n643), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  XOR2_X1   g451(.A(G134gat), .B(G162gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n640), .B(new_n647), .C1(KEYINPUT102), .C2(new_n641), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n650), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n654), .B1(new_n650), .B2(new_n655), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n629), .A2(new_n637), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n588), .A2(new_n589), .B1(new_n594), .B2(new_n597), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n627), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT103), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n628), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n667), .B(new_n668), .C1(new_n662), .C2(new_n638), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n638), .A2(KEYINPUT10), .A3(new_n662), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n660), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n667), .B1(new_n662), .B2(new_n638), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n660), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  OR2_X1    g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n613), .A2(new_n658), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n568), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n290), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  INV_X1    g484(.A(new_n378), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G8gat), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  NAND3_X1  g489(.A1(new_n682), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n689), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n692), .A2(KEYINPUT104), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(KEYINPUT104), .ZN(new_n694));
  OAI221_X1 g493(.A(new_n688), .B1(new_n689), .B2(new_n691), .C1(new_n693), .C2(new_n694), .ZN(G1325gat));
  NAND2_X1  g494(.A1(new_n474), .A2(new_n476), .ZN(new_n696));
  AOI21_X1  g495(.A(G15gat), .B1(new_n682), .B2(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n478), .A2(KEYINPUT105), .A3(new_n479), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT105), .B1(new_n478), .B2(new_n479), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n526), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT106), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n697), .B1(new_n682), .B2(new_n702), .ZN(G1326gat));
  NAND2_X1  g502(.A1(new_n682), .A2(new_n410), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  NAND2_X1  g505(.A1(new_n612), .A2(new_n680), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n658), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n290), .A2(G29gat), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n492), .A2(new_n567), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n711), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n489), .B1(new_n484), .B2(KEYINPUT35), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n700), .B2(new_n446), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n718), .B2(new_n658), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n658), .A2(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n379), .A2(new_n410), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n425), .A2(new_n445), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n721), .A2(new_n480), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n723), .B2(new_n717), .ZN(new_n724));
  INV_X1    g523(.A(new_n567), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n707), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n719), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n290), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n715), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT109), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n730), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n728), .A4(new_n715), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n492), .A2(new_n567), .A3(new_n708), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n736), .A2(G36gat), .A3(new_n378), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n727), .B2(new_n378), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1329gat));
  OAI21_X1  g539(.A(G43gat), .B1(new_n727), .B2(new_n700), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n696), .A2(new_n507), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1330gat));
  OAI21_X1  g544(.A(G50gat), .B1(new_n727), .B2(new_n409), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n410), .A2(new_n509), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n736), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1331gat));
  NAND3_X1  g549(.A1(new_n613), .A2(new_n658), .A3(new_n679), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n718), .A2(new_n567), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n683), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT110), .B(G57gat), .Z(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1332gat));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n686), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT49), .B(G64gat), .Z(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(G1333gat));
  INV_X1    g558(.A(G71gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n752), .A2(new_n760), .A3(new_n696), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n480), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n478), .A2(KEYINPUT105), .A3(new_n479), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n752), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n761), .B1(new_n766), .B2(new_n760), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n410), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n613), .A2(new_n567), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n679), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n763), .A2(new_n721), .A3(new_n722), .A4(new_n764), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n658), .B1(new_n774), .B2(new_n491), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n724), .B(new_n773), .C1(new_n775), .C2(KEYINPUT44), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n719), .A2(KEYINPUT111), .A3(new_n724), .A4(new_n773), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n683), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G85gat), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n771), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT51), .B1(new_n775), .B2(new_n771), .ZN(new_n784));
  OR3_X1    g583(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT112), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(KEYINPUT112), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n290), .A2(G85gat), .A3(new_n680), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT113), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n782), .B1(new_n787), .B2(new_n789), .ZN(G1336gat));
  NAND3_X1  g589(.A1(new_n778), .A2(new_n686), .A3(new_n779), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(G92gat), .ZN(new_n792));
  INV_X1    g591(.A(G92gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n686), .A2(new_n793), .A3(new_n679), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT114), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n783), .B2(new_n784), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(KEYINPUT115), .B(new_n795), .C1(new_n783), .C2(new_n784), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT52), .B1(new_n792), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n786), .A3(new_n795), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  OAI21_X1  g602(.A(G92gat), .B1(new_n776), .B2(new_n378), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(new_n805), .ZN(G1337gat));
  NAND2_X1  g605(.A1(new_n780), .A2(new_n765), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G99gat), .ZN(new_n808));
  AOI211_X1 g607(.A(G99gat), .B(new_n680), .C1(new_n476), .C2(new_n474), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT116), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n787), .B2(new_n810), .ZN(G1338gat));
  NOR3_X1   g610(.A1(new_n680), .A2(G106gat), .A3(new_n409), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n785), .A2(new_n786), .A3(new_n812), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n776), .A2(new_n409), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT53), .B1(new_n814), .B2(G106gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n778), .A2(new_n410), .A3(new_n779), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n783), .A2(new_n784), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n817), .A2(G106gat), .B1(new_n818), .B2(new_n812), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(G1339gat));
  NAND4_X1  g620(.A1(new_n613), .A2(new_n725), .A3(new_n658), .A4(new_n680), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n564), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n549), .A2(new_n553), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n825), .A2(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n824), .A2(new_n561), .B1(new_n496), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n679), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n829), .B(new_n676), .C1(new_n671), .C2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n669), .A2(new_n660), .A3(new_n670), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n669), .A2(new_n670), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n659), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n669), .A2(KEYINPUT117), .A3(new_n660), .A4(new_n670), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT54), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n831), .A2(new_n838), .A3(KEYINPUT118), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n678), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n676), .B1(new_n671), .B2(new_n830), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n829), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n567), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n828), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n658), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n842), .A2(new_n678), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT118), .B1(new_n831), .B2(new_n838), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT55), .B1(new_n838), .B2(new_n844), .ZN(new_n852));
  NOR4_X1   g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n658), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n827), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n613), .B1(new_n855), .B2(KEYINPUT119), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n848), .A2(new_n658), .B1(new_n853), .B2(new_n827), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n823), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n483), .ZN(new_n861));
  NOR4_X1   g660(.A1(new_n860), .A2(new_n290), .A3(new_n686), .A4(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT120), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n725), .A2(new_n217), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n290), .A2(new_n686), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n696), .A2(new_n409), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n860), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G113gat), .B1(new_n870), .B2(new_n725), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n865), .A2(new_n871), .ZN(G1340gat));
  NAND3_X1  g671(.A1(new_n863), .A2(new_n205), .A3(new_n679), .ZN(new_n873));
  OAI21_X1  g672(.A(G120gat), .B1(new_n870), .B2(new_n680), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1341gat));
  NAND3_X1  g674(.A1(new_n869), .A2(new_n243), .A3(new_n613), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n243), .B1(new_n862), .B2(new_n613), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G1342gat));
  INV_X1    g680(.A(new_n658), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n862), .A2(new_n210), .A3(new_n882), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  OAI21_X1  g683(.A(G134gat), .B1(new_n870), .B2(new_n658), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G1343gat));
  NOR2_X1   g686(.A1(new_n765), .A2(new_n867), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n612), .B1(new_n857), .B2(new_n858), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n849), .A2(new_n858), .A3(new_n854), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n822), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n891), .B2(new_n410), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n855), .A2(new_n612), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n822), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n409), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n567), .B(new_n888), .C1(new_n892), .C2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT122), .B1(new_n898), .B2(G141gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n700), .A2(new_n378), .A3(new_n410), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n725), .A2(G141gat), .ZN(new_n901));
  NOR4_X1   g700(.A1(new_n860), .A2(new_n290), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n898), .B2(G141gat), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n899), .A2(new_n903), .A3(KEYINPUT58), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  AOI221_X4 g704(.A(new_n902), .B1(KEYINPUT122), .B2(new_n905), .C1(new_n898), .C2(G141gat), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n904), .A2(new_n906), .ZN(G1344gat));
  NOR3_X1   g706(.A1(new_n860), .A2(new_n290), .A3(new_n900), .ZN(new_n908));
  INV_X1    g707(.A(G148gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n679), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n700), .A2(new_n866), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n915), .A3(new_n679), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n853), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n846), .A2(new_n882), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT124), .B1(new_n843), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n827), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n613), .B1(new_n921), .B2(new_n849), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n410), .B1(new_n922), .B2(new_n823), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n895), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n891), .A2(new_n896), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n916), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n909), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n911), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n892), .ZN(new_n931));
  INV_X1    g730(.A(new_n897), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n913), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI211_X1 g732(.A(KEYINPUT59), .B(new_n909), .C1(new_n933), .C2(new_n679), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n910), .B1(new_n930), .B2(new_n934), .ZN(G1345gat));
  AND2_X1   g734(.A1(new_n908), .A2(new_n613), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G155gat), .B1(new_n936), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n612), .A2(new_n608), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n938), .A2(new_n939), .B1(new_n933), .B2(new_n940), .ZN(G1346gat));
  INV_X1    g740(.A(G162gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n908), .A2(new_n942), .A3(new_n882), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n933), .A2(new_n882), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n942), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n860), .A2(new_n683), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n861), .A2(new_n378), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n567), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n683), .A2(new_n378), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n860), .A2(new_n868), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n725), .A2(new_n308), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(G1348gat));
  AOI21_X1  g753(.A(G176gat), .B1(new_n948), .B2(new_n679), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n679), .A2(new_n313), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n952), .B2(new_n956), .ZN(G1349gat));
  AND2_X1   g756(.A1(new_n613), .A2(new_n326), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n952), .A2(new_n613), .ZN(new_n959));
  AOI22_X1  g758(.A1(new_n948), .A2(new_n958), .B1(new_n959), .B2(G183gat), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT60), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n960), .B(new_n961), .ZN(G1350gat));
  NAND3_X1  g761(.A1(new_n948), .A2(new_n327), .A3(new_n882), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n952), .A2(new_n882), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G190gat), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1351gat));
  NOR3_X1   g767(.A1(new_n765), .A2(new_n378), .A3(new_n409), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n946), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(G197gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n970), .A2(new_n971), .A3(new_n567), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n924), .A2(new_n925), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n765), .A2(new_n951), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n976), .B2(new_n725), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G197gat), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n976), .A2(new_n973), .A3(new_n725), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n972), .B1(new_n978), .B2(new_n979), .ZN(G1352gat));
  INV_X1    g779(.A(G204gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n970), .A2(new_n981), .A3(new_n679), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  OAI21_X1  g782(.A(G204gat), .B1(new_n976), .B2(new_n680), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(G1353gat));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n348), .A3(new_n613), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n974), .A2(new_n613), .A3(new_n975), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  OAI21_X1  g790(.A(G218gat), .B1(new_n976), .B2(new_n658), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n970), .A2(new_n349), .A3(new_n882), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1355gat));
endmodule


