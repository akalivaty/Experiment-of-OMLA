

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U325 ( .A(n442), .B(n373), .ZN(n374) );
  INV_X1 U326 ( .A(KEYINPUT54), .ZN(n418) );
  XNOR2_X1 U327 ( .A(n418), .B(KEYINPUT122), .ZN(n419) );
  XNOR2_X1 U328 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U329 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U330 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U331 ( .A(n385), .B(n384), .ZN(n477) );
  XNOR2_X1 U332 ( .A(n458), .B(G176GAT), .ZN(n459) );
  XNOR2_X1 U333 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  INV_X1 U334 ( .A(G92GAT), .ZN(n293) );
  NAND2_X1 U335 ( .A1(n293), .A2(G64GAT), .ZN(n296) );
  INV_X1 U336 ( .A(G64GAT), .ZN(n294) );
  NAND2_X1 U337 ( .A1(n294), .A2(G92GAT), .ZN(n295) );
  NAND2_X1 U338 ( .A1(n296), .A2(n295), .ZN(n298) );
  XNOR2_X1 U339 ( .A(G176GAT), .B(G204GAT), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n398) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G71GAT), .Z(n440) );
  XNOR2_X1 U342 ( .A(n398), .B(n440), .ZN(n300) );
  AND2_X1 U343 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U345 ( .A(KEYINPUT32), .B(n301), .Z(n303) );
  XOR2_X1 U346 ( .A(G57GAT), .B(KEYINPUT13), .Z(n353) );
  XNOR2_X1 U347 ( .A(n353), .B(KEYINPUT74), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U349 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n305) );
  XNOR2_X1 U350 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n304) );
  XOR2_X1 U351 ( .A(n305), .B(n304), .Z(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n311) );
  XNOR2_X1 U353 ( .A(G106GAT), .B(G78GAT), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n308), .B(G148GAT), .ZN(n427) );
  XNOR2_X1 U355 ( .A(G99GAT), .B(G85GAT), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n309), .B(KEYINPUT72), .ZN(n378) );
  XNOR2_X1 U357 ( .A(n427), .B(n378), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n392) );
  XNOR2_X1 U359 ( .A(n392), .B(KEYINPUT41), .ZN(n555) );
  XNOR2_X1 U360 ( .A(KEYINPUT106), .B(n555), .ZN(n542) );
  XOR2_X1 U361 ( .A(G57GAT), .B(KEYINPUT4), .Z(n313) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(KEYINPUT88), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n318) );
  XNOR2_X1 U364 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n314), .B(KEYINPUT2), .ZN(n426) );
  XOR2_X1 U366 ( .A(G85GAT), .B(n426), .Z(n316) );
  XOR2_X1 U367 ( .A(G113GAT), .B(KEYINPUT0), .Z(n441) );
  XNOR2_X1 U368 ( .A(n441), .B(G162GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n331) );
  XOR2_X1 U371 ( .A(G120GAT), .B(G127GAT), .Z(n320) );
  XNOR2_X1 U372 ( .A(G29GAT), .B(G134GAT), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U374 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n322) );
  XNOR2_X1 U375 ( .A(G141GAT), .B(G148GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U377 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U378 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n326) );
  NAND2_X1 U379 ( .A1(G225GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U381 ( .A(KEYINPUT90), .B(n327), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n523) );
  XNOR2_X1 U384 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n332), .B(G8GAT), .ZN(n355) );
  XOR2_X1 U386 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U387 ( .A(n355), .B(n431), .Z(n334) );
  XNOR2_X1 U388 ( .A(G50GAT), .B(G36GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n339) );
  XNOR2_X1 U390 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n335), .B(KEYINPUT7), .ZN(n379) );
  XOR2_X1 U392 ( .A(n379), .B(KEYINPUT70), .Z(n337) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U395 ( .A(n339), .B(n338), .Z(n347) );
  XOR2_X1 U396 ( .A(G15GAT), .B(G113GAT), .Z(n341) );
  XNOR2_X1 U397 ( .A(G169GAT), .B(G43GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U399 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n343) );
  XNOR2_X1 U400 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n573) );
  NAND2_X1 U404 ( .A1(n573), .A2(n555), .ZN(n350) );
  XOR2_X1 U405 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n348) );
  XNOR2_X1 U406 ( .A(KEYINPUT115), .B(n348), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n387) );
  XOR2_X1 U408 ( .A(KEYINPUT79), .B(G64GAT), .Z(n352) );
  XNOR2_X1 U409 ( .A(G211GAT), .B(G155GAT), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U411 ( .A(n354), .B(n353), .Z(n357) );
  XOR2_X1 U412 ( .A(G15GAT), .B(G127GAT), .Z(n439) );
  XNOR2_X1 U413 ( .A(n355), .B(n439), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U415 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n359) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U418 ( .A(n361), .B(n360), .Z(n366) );
  XOR2_X1 U419 ( .A(G78GAT), .B(G71GAT), .Z(n363) );
  XNOR2_X1 U420 ( .A(G22GAT), .B(G183GAT), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n364), .B(KEYINPUT12), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n582) );
  XOR2_X1 U424 ( .A(KEYINPUT75), .B(KEYINPUT67), .Z(n368) );
  XNOR2_X1 U425 ( .A(G218GAT), .B(KEYINPUT76), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U427 ( .A(KEYINPUT10), .B(G92GAT), .Z(n370) );
  XNOR2_X1 U428 ( .A(G190GAT), .B(G106GAT), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U430 ( .A(n372), .B(n371), .Z(n377) );
  XOR2_X1 U431 ( .A(G36GAT), .B(KEYINPUT77), .Z(n399) );
  XOR2_X1 U432 ( .A(G50GAT), .B(G162GAT), .Z(n425) );
  XOR2_X1 U433 ( .A(n399), .B(n425), .Z(n375) );
  XOR2_X1 U434 ( .A(G43GAT), .B(G134GAT), .Z(n442) );
  NAND2_X1 U435 ( .A1(G232GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n385) );
  XOR2_X1 U437 ( .A(n379), .B(n378), .Z(n383) );
  XOR2_X1 U438 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n381) );
  XNOR2_X1 U439 ( .A(KEYINPUT65), .B(KEYINPUT11), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n382) );
  INV_X1 U441 ( .A(n477), .ZN(n567) );
  NOR2_X1 U442 ( .A1(n582), .A2(n567), .ZN(n386) );
  AND2_X1 U443 ( .A1(n387), .A2(n386), .ZN(n389) );
  INV_X1 U444 ( .A(KEYINPUT47), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n396) );
  XOR2_X1 U446 ( .A(KEYINPUT36), .B(n477), .Z(n584) );
  NAND2_X1 U447 ( .A1(n582), .A2(n584), .ZN(n391) );
  XOR2_X1 U448 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n393) );
  BUF_X1 U450 ( .A(n392), .Z(n577) );
  NAND2_X1 U451 ( .A1(n393), .A2(n577), .ZN(n394) );
  NOR2_X1 U452 ( .A1(n573), .A2(n394), .ZN(n395) );
  NOR2_X1 U453 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n397), .B(KEYINPUT48), .ZN(n536) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n401) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U458 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n403) );
  XNOR2_X1 U459 ( .A(G8GAT), .B(KEYINPUT91), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U461 ( .A(n405), .B(n404), .Z(n416) );
  XOR2_X1 U462 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n407) );
  XNOR2_X1 U463 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U465 ( .A(n408), .B(KEYINPUT84), .Z(n410) );
  XNOR2_X1 U466 ( .A(G169GAT), .B(G183GAT), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n451) );
  XOR2_X1 U468 ( .A(KEYINPUT21), .B(G218GAT), .Z(n412) );
  XNOR2_X1 U469 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U471 ( .A(G197GAT), .B(n413), .ZN(n436) );
  INV_X1 U472 ( .A(n436), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n451), .B(n414), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n526) );
  XNOR2_X1 U475 ( .A(n526), .B(KEYINPUT121), .ZN(n417) );
  NOR2_X1 U476 ( .A1(n536), .A2(n417), .ZN(n420) );
  NOR2_X1 U477 ( .A1(n523), .A2(n421), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n422), .B(KEYINPUT64), .ZN(n572) );
  XOR2_X1 U479 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT87), .B(G204GAT), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n435) );
  XOR2_X1 U482 ( .A(n426), .B(n425), .Z(n433) );
  XOR2_X1 U483 ( .A(n427), .B(KEYINPUT23), .Z(n429) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n467) );
  NAND2_X1 U490 ( .A1(n572), .A2(n467), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n438), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U492 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n455) );
  XOR2_X1 U495 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n446) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U498 ( .A(n447), .B(KEYINPUT80), .Z(n453) );
  XOR2_X1 U499 ( .A(KEYINPUT81), .B(G176GAT), .Z(n449) );
  XNOR2_X1 U500 ( .A(G99GAT), .B(KEYINPUT20), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X2 U504 ( .A(n455), .B(n454), .Z(n538) );
  NAND2_X1 U505 ( .A1(n456), .A2(n538), .ZN(n457) );
  XNOR2_X1 U506 ( .A(n457), .B(KEYINPUT123), .ZN(n568) );
  NAND2_X1 U507 ( .A1(n542), .A2(n568), .ZN(n460) );
  XOR2_X1 U508 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n458) );
  XOR2_X1 U509 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n482) );
  NAND2_X1 U510 ( .A1(n573), .A2(n577), .ZN(n496) );
  XNOR2_X1 U511 ( .A(KEYINPUT28), .B(n467), .ZN(n489) );
  XNOR2_X1 U512 ( .A(n526), .B(KEYINPUT27), .ZN(n469) );
  NAND2_X1 U513 ( .A1(n523), .A2(n469), .ZN(n535) );
  XOR2_X1 U514 ( .A(n538), .B(KEYINPUT85), .Z(n461) );
  NOR2_X1 U515 ( .A1(n535), .A2(n461), .ZN(n462) );
  NAND2_X1 U516 ( .A1(n489), .A2(n462), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n463), .B(KEYINPUT94), .ZN(n475) );
  NAND2_X1 U518 ( .A1(n526), .A2(n538), .ZN(n464) );
  NAND2_X1 U519 ( .A1(n464), .A2(n467), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n465), .B(KEYINPUT95), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n466), .B(KEYINPUT25), .ZN(n471) );
  NOR2_X1 U522 ( .A1(n467), .A2(n538), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n468), .B(KEYINPUT26), .ZN(n571) );
  NAND2_X1 U524 ( .A1(n469), .A2(n571), .ZN(n470) );
  NAND2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n473) );
  INV_X1 U526 ( .A(n523), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U528 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U529 ( .A(KEYINPUT96), .B(n476), .Z(n493) );
  NAND2_X1 U530 ( .A1(n477), .A2(n582), .ZN(n478) );
  XNOR2_X1 U531 ( .A(KEYINPUT16), .B(n478), .ZN(n479) );
  OR2_X1 U532 ( .A1(n493), .A2(n479), .ZN(n510) );
  NOR2_X1 U533 ( .A1(n496), .A2(n510), .ZN(n480) );
  XOR2_X1 U534 ( .A(KEYINPUT97), .B(n480), .Z(n490) );
  NAND2_X1 U535 ( .A1(n490), .A2(n523), .ZN(n481) );
  XNOR2_X1 U536 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  XOR2_X1 U538 ( .A(G8GAT), .B(KEYINPUT99), .Z(n485) );
  NAND2_X1 U539 ( .A1(n490), .A2(n526), .ZN(n484) );
  XNOR2_X1 U540 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U542 ( .A1(n490), .A2(n538), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U544 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  XOR2_X1 U545 ( .A(G22GAT), .B(KEYINPUT101), .Z(n492) );
  INV_X1 U546 ( .A(n489), .ZN(n540) );
  NAND2_X1 U547 ( .A1(n490), .A2(n540), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n492), .B(n491), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  NOR2_X1 U550 ( .A1(n582), .A2(n493), .ZN(n494) );
  NAND2_X1 U551 ( .A1(n494), .A2(n584), .ZN(n495) );
  XOR2_X1 U552 ( .A(KEYINPUT37), .B(n495), .Z(n520) );
  NOR2_X1 U553 ( .A1(n520), .A2(n496), .ZN(n498) );
  XNOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n498), .B(n497), .ZN(n506) );
  NAND2_X1 U556 ( .A1(n506), .A2(n523), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  XOR2_X1 U558 ( .A(G36GAT), .B(KEYINPUT103), .Z(n502) );
  NAND2_X1 U559 ( .A1(n506), .A2(n526), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(G1329GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n504) );
  NAND2_X1 U562 ( .A1(n506), .A2(n538), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U564 ( .A(G43GAT), .B(n505), .Z(G1330GAT) );
  XOR2_X1 U565 ( .A(G50GAT), .B(KEYINPUT105), .Z(n508) );
  NAND2_X1 U566 ( .A1(n506), .A2(n540), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n508), .B(n507), .ZN(G1331GAT) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n513) );
  INV_X1 U569 ( .A(n573), .ZN(n551) );
  NAND2_X1 U570 ( .A1(n551), .A2(n542), .ZN(n509) );
  XOR2_X1 U571 ( .A(KEYINPUT107), .B(n509), .Z(n521) );
  NOR2_X1 U572 ( .A1(n510), .A2(n521), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(KEYINPUT108), .ZN(n517) );
  NAND2_X1 U574 ( .A1(n523), .A2(n517), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n517), .A2(n526), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U578 ( .A(G71GAT), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U579 ( .A1(n538), .A2(n517), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U582 ( .A1(n517), .A2(n540), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  XOR2_X1 U584 ( .A(G85GAT), .B(KEYINPUT111), .Z(n525) );
  NOR2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(KEYINPUT110), .ZN(n531) );
  NAND2_X1 U587 ( .A1(n523), .A2(n531), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n528) );
  NAND2_X1 U590 ( .A1(n526), .A2(n531), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n531), .A2(n538), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n533) );
  NAND2_X1 U596 ( .A1(n531), .A2(n540), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U598 ( .A(G106GAT), .B(n534), .Z(G1339GAT) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT117), .B(n537), .Z(n550) );
  NAND2_X1 U601 ( .A1(n538), .A2(n550), .ZN(n539) );
  NOR2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n573), .A2(n547), .ZN(n541) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U606 ( .A1(n547), .A2(n542), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n547), .A2(n582), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U612 ( .A1(n547), .A2(n567), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n550), .A2(n571), .ZN(n554) );
  NOR2_X1 U615 ( .A1(n551), .A2(n554), .ZN(n552) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n552), .Z(n553) );
  XNOR2_X1 U617 ( .A(KEYINPUT118), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  INV_X1 U619 ( .A(n554), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n562), .A2(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n560) );
  NAND2_X1 U624 ( .A1(n562), .A2(n582), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n567), .A2(n562), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n568), .A2(n573), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT124), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n568), .A2(n582), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  AND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n585) );
  NAND2_X1 U638 ( .A1(n585), .A2(n573), .ZN(n576) );
  XOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT60), .Z(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT59), .B(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  INV_X1 U643 ( .A(n577), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(G218GAT), .B(n588), .Z(G1355GAT) );
endmodule

