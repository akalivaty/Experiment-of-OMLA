//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT64), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216));
  INV_X1    g015(.A(G169gat), .ZN(new_n217));
  INV_X1    g016(.A(G176gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(G169gat), .A3(G176gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n215), .A2(new_n219), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n227), .A2(new_n210), .A3(new_n228), .A4(new_n211), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n224), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(KEYINPUT66), .A3(new_n231), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n227), .A2(KEYINPUT67), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n213), .A2(new_n237), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n236), .A2(new_n238), .A3(new_n212), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n215), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n223), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT25), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n234), .A2(new_n235), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n209), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT68), .A3(KEYINPUT28), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  OR3_X1    g048(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(new_n209), .A3(new_n246), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n248), .A2(new_n225), .A3(new_n251), .A4(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT29), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n207), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT75), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G211gat), .A2(G218gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT74), .ZN(new_n264));
  INV_X1    g063(.A(G197gat), .ZN(new_n265));
  INV_X1    g064(.A(G204gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G197gat), .A2(G204gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(new_n262), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n261), .A2(new_n271), .A3(new_n262), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n264), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n270), .B1(new_n264), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n258), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n270), .ZN(new_n276));
  INV_X1    g075(.A(new_n272), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n271), .B1(new_n261), .B2(new_n262), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n270), .A3(new_n272), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(KEYINPUT75), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n254), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n243), .B1(new_n232), .B2(new_n233), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(new_n235), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n283), .B1(new_n286), .B2(new_n206), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n257), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n206), .B1(new_n286), .B2(KEYINPUT29), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n255), .A2(new_n207), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n205), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n206), .B1(new_n245), .B2(new_n254), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n282), .B1(new_n257), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n289), .A2(new_n283), .A3(new_n290), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n204), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT76), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT76), .B(KEYINPUT30), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n294), .A2(new_n295), .A3(new_n204), .A4(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n302));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  INV_X1    g102(.A(G155gat), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n306), .B2(KEYINPUT2), .ZN(new_n307));
  AND2_X1   g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT78), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n303), .A2(new_n312), .A3(KEYINPUT2), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G141gat), .B(G148gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n312), .B1(new_n303), .B2(KEYINPUT2), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT77), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(new_n304), .A3(new_n305), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n303), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n311), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G134gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G127gat), .ZN(new_n325));
  INV_X1    g124(.A(G127gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G134gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G113gat), .B(G120gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT1), .ZN(new_n333));
  INV_X1    g132(.A(G113gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(G120gat), .ZN(new_n335));
  INV_X1    g134(.A(G120gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(G113gat), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT70), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n339), .A2(new_n325), .A3(new_n327), .A4(new_n340), .ZN(new_n341));
  OAI22_X1  g140(.A1(new_n331), .A2(new_n333), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n302), .B1(new_n323), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n330), .ZN(new_n344));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n344), .B1(new_n328), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n340), .B1(new_n335), .B2(new_n337), .ZN(new_n347));
  INV_X1    g146(.A(new_n341), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n346), .A2(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n303), .A2(KEYINPUT2), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT78), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(new_n310), .A3(new_n313), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n319), .A2(new_n320), .B1(G155gat), .B2(G162gat), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n354), .A2(new_n355), .B1(new_n310), .B2(new_n307), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(KEYINPUT4), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n342), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n355), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n360), .A2(new_n358), .A3(new_n311), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n343), .B(new_n357), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT79), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n323), .A2(new_n342), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n347), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n350), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n356), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n364), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n365), .A2(KEYINPUT5), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n356), .B(new_n342), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT5), .B1(new_n373), .B2(new_n363), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n323), .A2(KEYINPUT3), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n358), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n342), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n377), .A2(new_n363), .A3(new_n343), .A4(new_n357), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n378), .A3(KEYINPUT79), .ZN(new_n379));
  XOR2_X1   g178(.A(G1gat), .B(G29gat), .Z(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT0), .ZN(new_n381));
  XNOR2_X1  g180(.A(G57gat), .B(G85gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n372), .A2(KEYINPUT6), .A3(new_n379), .A4(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n379), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n374), .B1(KEYINPUT79), .B2(new_n378), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n379), .A3(new_n384), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n299), .A2(new_n301), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n351), .B(new_n284), .C1(new_n285), .C2(new_n235), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n342), .B1(new_n245), .B2(new_n254), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G227gat), .ZN(new_n396));
  INV_X1    g195(.A(G233gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT34), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n230), .A2(KEYINPUT66), .A3(new_n231), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT66), .B1(new_n230), .B2(new_n231), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n400), .A2(new_n401), .A3(new_n243), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n351), .B1(new_n402), .B2(new_n284), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n245), .A2(new_n342), .A3(new_n254), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT34), .ZN(new_n406));
  INV_X1    g205(.A(new_n398), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT33), .B1(new_n395), .B2(new_n398), .ZN(new_n409));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT73), .ZN(new_n411));
  XOR2_X1   g210(.A(G71gat), .B(G99gat), .Z(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n399), .B(new_n408), .C1(new_n409), .C2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n403), .A2(new_n398), .A3(new_n404), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT33), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n420));
  AOI211_X1 g219(.A(KEYINPUT34), .B(new_n398), .C1(new_n403), .C2(new_n404), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(KEYINPUT32), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n424), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n416), .A2(new_n426), .A3(new_n422), .ZN(new_n427));
  XNOR2_X1  g226(.A(G78gat), .B(G106gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT31), .B(G50gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT80), .ZN(new_n431));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n256), .B1(new_n273), .B2(new_n274), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n358), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n323), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n281), .A2(new_n275), .B1(new_n376), .B2(new_n256), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(KEYINPUT81), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n376), .A2(new_n256), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n282), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n432), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(G22gat), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n438), .A2(KEYINPUT82), .B1(new_n281), .B2(new_n275), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT82), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n376), .A2(new_n445), .A3(new_n256), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n432), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n435), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n442), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n443), .B1(new_n442), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n431), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n356), .B1(new_n433), .B2(new_n358), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n439), .B2(new_n440), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n448), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI211_X1 g256(.A(new_n432), .B(new_n454), .C1(new_n444), .C2(new_n446), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n453), .B(G22gat), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n442), .B(new_n449), .C1(KEYINPUT83), .C2(new_n443), .ZN(new_n460));
  INV_X1    g259(.A(new_n430), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n452), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n392), .A2(new_n425), .A3(new_n427), .A4(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(KEYINPUT35), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT91), .B(KEYINPUT35), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n257), .B2(new_n287), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n205), .B1(new_n472), .B2(new_n291), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n294), .B2(new_n295), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT38), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT90), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n291), .A2(KEYINPUT89), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n295), .B1(new_n291), .B2(KEYINPUT89), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT37), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT38), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(new_n205), .C1(new_n472), .C2(new_n291), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n391), .A2(new_n385), .A3(new_n296), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT90), .B(KEYINPUT38), .C1(new_n473), .C2(new_n474), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n477), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n386), .A2(new_n387), .A3(new_n383), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT40), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n490));
  NAND2_X1  g289(.A1(new_n343), .A2(new_n357), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n359), .A2(new_n361), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n364), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n383), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n366), .A2(new_n369), .A3(new_n363), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT39), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n364), .B2(new_n362), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n489), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(KEYINPUT86), .B(new_n489), .C1(new_n494), .C2(new_n497), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n488), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n362), .A2(new_n364), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n495), .A2(KEYINPUT39), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n505), .A2(KEYINPUT40), .A3(new_n383), .A4(new_n493), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n323), .A2(new_n342), .A3(new_n302), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT4), .B1(new_n351), .B2(new_n356), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n363), .B1(new_n511), .B2(new_n377), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n384), .B1(new_n512), .B2(new_n490), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n513), .A2(KEYINPUT87), .A3(KEYINPUT40), .A4(new_n505), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n502), .A2(new_n299), .A3(new_n301), .A4(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(KEYINPUT88), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT88), .ZN(new_n518));
  INV_X1    g317(.A(new_n501), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n383), .B(new_n493), .C1(new_n512), .C2(new_n496), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT86), .B1(new_n520), .B2(new_n489), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n390), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n508), .A2(new_n514), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND4_X1   g323(.A1(new_n294), .A2(new_n295), .A3(new_n204), .A4(new_n300), .ZN(new_n525));
  INV_X1    g324(.A(new_n298), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n256), .B1(new_n402), .B2(new_n284), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n293), .B1(new_n527), .B2(new_n206), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n295), .B1(new_n528), .B2(new_n283), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(new_n529), .B2(new_n205), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n525), .B1(new_n530), .B2(new_n296), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n518), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n463), .B(new_n487), .C1(new_n517), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n299), .A2(new_n301), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n391), .A2(new_n385), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n463), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n416), .A2(new_n426), .A3(new_n422), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n426), .B1(new_n416), .B2(new_n422), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n425), .A2(KEYINPUT36), .A3(new_n427), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n533), .B1(new_n534), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n543), .A2(new_n534), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n470), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n470), .B(KEYINPUT92), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G50gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G43gat), .ZN(new_n552));
  INV_X1    g351(.A(G43gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(G50gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n554), .A3(KEYINPUT15), .ZN(new_n555));
  NAND2_X1  g354(.A1(G29gat), .A2(G36gat), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR3_X1   g358(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n552), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n561), .A2(KEYINPUT96), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n554), .B1(new_n561), .B2(KEYINPUT96), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI221_X1 g363(.A(new_n557), .B1(new_n559), .B2(new_n560), .C1(new_n564), .C2(KEYINPUT15), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n560), .B1(new_n566), .B2(new_n558), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n566), .B2(new_n558), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n556), .ZN(new_n569));
  INV_X1    g368(.A(new_n555), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n569), .A2(KEYINPUT95), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT95), .B1(new_n569), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n565), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G15gat), .B(G22gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT16), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(G1gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(G1gat), .B2(new_n576), .ZN(new_n579));
  INV_X1    g378(.A(G8gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n573), .B2(new_n574), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n575), .A2(new_n583), .B1(new_n573), .B2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(KEYINPUT18), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n588), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n573), .B(new_n582), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n585), .B(KEYINPUT13), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G197gat), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT11), .B(G169gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT93), .B(KEYINPUT12), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n594), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G57gat), .B(G64gat), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT9), .ZN(new_n606));
  INV_X1    g405(.A(G71gat), .ZN(new_n607));
  INV_X1    g406(.A(G78gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(KEYINPUT98), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n606), .B(new_n611), .C1(KEYINPUT98), .C2(new_n610), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT99), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT100), .B1(new_n609), .B2(KEYINPUT9), .ZN(new_n614));
  NOR2_X1   g413(.A1(KEYINPUT100), .A2(KEYINPUT9), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n614), .B(new_n605), .C1(new_n609), .C2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT101), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G127gat), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n613), .A2(new_n618), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n582), .B1(new_n625), .B2(KEYINPUT21), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT102), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n624), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n304), .ZN(new_n630));
  XOR2_X1   g429(.A(G183gat), .B(G211gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n628), .A2(new_n632), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G190gat), .B(G218gat), .Z(new_n636));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n637));
  NAND2_X1  g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638));
  OAI22_X1  g437(.A1(new_n636), .A2(KEYINPUT105), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G85gat), .A2(G92gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT7), .ZN(new_n641));
  NAND2_X1  g440(.A1(G99gat), .A2(G106gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT8), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n641), .B(new_n643), .C1(G85gat), .C2(G92gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G99gat), .B(G106gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n645), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n644), .A2(KEYINPUT103), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT104), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n639), .B1(new_n652), .B2(new_n573), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n651), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n573), .A2(new_n574), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n575), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n636), .A2(KEYINPUT105), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(G134gat), .B(G162gat), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n638), .A2(new_n637), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n635), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n625), .A2(new_n646), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT106), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n668), .B(KEYINPUT106), .C1(new_n625), .C2(new_n651), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT10), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n652), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n672));
  INV_X1    g471(.A(G230gat), .ZN(new_n673));
  OAI22_X1  g472(.A1(new_n671), .A2(new_n672), .B1(new_n673), .B2(new_n397), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n397), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n674), .A2(new_n677), .A3(new_n681), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n667), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n550), .A2(new_n604), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n536), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT107), .B(G1gat), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1324gat));
  INV_X1    g489(.A(new_n687), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n580), .B1(new_n691), .B2(new_n531), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT16), .B(G8gat), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n687), .A2(new_n535), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT42), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(KEYINPUT42), .B2(new_n694), .ZN(G1325gat));
  INV_X1    g495(.A(G15gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n541), .A2(new_n542), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n687), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n425), .A2(new_n427), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n697), .B1(new_n687), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n699), .B1(new_n703), .B2(new_n704), .ZN(G1326gat));
  NOR2_X1   g504(.A1(new_n687), .A2(new_n463), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT43), .B(G22gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n666), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n548), .A2(new_n549), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n470), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n516), .B(new_n518), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n487), .A2(new_n463), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n543), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n533), .A2(new_n717), .A3(new_n543), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n712), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n709), .B1(new_n719), .B2(new_n666), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n711), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n635), .ZN(new_n722));
  INV_X1    g521(.A(new_n685), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n604), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n536), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n724), .A2(new_n666), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n550), .A2(new_n604), .A3(new_n730), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n536), .A2(G29gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n731), .A2(new_n729), .A3(new_n732), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n728), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n728), .A2(new_n734), .A3(KEYINPUT110), .A4(new_n733), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1328gat));
  NOR3_X1   g538(.A1(new_n731), .A2(G36gat), .A3(new_n535), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT46), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n727), .B2(new_n535), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1329gat));
  OAI21_X1  g542(.A(new_n553), .B1(new_n731), .B2(new_n700), .ZN(new_n744));
  INV_X1    g543(.A(new_n698), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n721), .A2(G43gat), .A3(new_n745), .A4(new_n726), .ZN(new_n746));
  NAND2_X1  g545(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n748), .B(new_n749), .Z(G1330gat));
  NOR3_X1   g549(.A1(new_n731), .A2(G50gat), .A3(new_n463), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(KEYINPUT48), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(KEYINPUT48), .ZN(new_n755));
  OAI21_X1  g554(.A(G50gat), .B1(new_n727), .B2(new_n463), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n755), .B1(new_n754), .B2(new_n756), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(G1331gat));
  NAND4_X1  g558(.A1(new_n635), .A2(new_n725), .A3(new_n666), .A4(new_n685), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n719), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n536), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g563(.A1(new_n719), .A2(new_n535), .A3(new_n760), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  AND2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n765), .B2(new_n766), .ZN(G1333gat));
  AOI21_X1  g568(.A(new_n607), .B1(new_n761), .B2(new_n745), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n700), .A2(G71gat), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n761), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1334gat));
  INV_X1    g573(.A(new_n463), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n761), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n533), .A2(new_n717), .A3(new_n543), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n717), .B1(new_n533), .B2(new_n543), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n470), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  INV_X1    g581(.A(new_n666), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n635), .A2(new_n604), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n778), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT114), .B1(new_n719), .B2(new_n666), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n790), .A2(new_n784), .A3(KEYINPUT51), .A4(new_n785), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(KEYINPUT115), .B(new_n778), .C1(new_n786), .C2(new_n787), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n536), .A2(G85gat), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n792), .A2(new_n685), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n785), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n723), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n721), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G85gat), .B1(new_n798), .B2(new_n536), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(G1336gat));
  NOR3_X1   g599(.A1(new_n723), .A2(G92gat), .A3(new_n535), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n792), .A2(new_n793), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n792), .A2(KEYINPUT116), .A3(new_n793), .A4(new_n801), .ZN(new_n805));
  XOR2_X1   g604(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n806));
  NAND3_X1  g605(.A1(new_n721), .A2(new_n531), .A3(new_n797), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(G92gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n807), .A2(G92gat), .ZN(new_n810));
  INV_X1    g609(.A(new_n801), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n788), .B2(new_n791), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT52), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n813), .ZN(G1337gat));
  XOR2_X1   g613(.A(KEYINPUT118), .B(G99gat), .Z(new_n815));
  NOR2_X1   g614(.A1(new_n700), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n792), .A2(new_n685), .A3(new_n793), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n798), .B2(new_n698), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1338gat));
  NOR3_X1   g618(.A1(new_n723), .A2(G106gat), .A3(new_n463), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n792), .A2(new_n793), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n711), .A2(new_n720), .A3(new_n775), .A4(new_n797), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n716), .A2(new_n718), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n666), .B1(new_n827), .B2(new_n470), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n796), .B1(new_n828), .B2(new_n782), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT51), .B1(new_n829), .B2(new_n790), .ZN(new_n830));
  INV_X1    g629(.A(new_n791), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n820), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n824), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n826), .B1(new_n833), .B2(KEYINPUT53), .ZN(new_n834));
  INV_X1    g633(.A(new_n820), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n788), .B2(new_n791), .ZN(new_n836));
  INV_X1    g635(.A(new_n824), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n826), .B(KEYINPUT53), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n825), .B1(new_n834), .B2(new_n839), .ZN(G1339gat));
  OAI21_X1  g639(.A(new_n682), .B1(new_n674), .B2(KEYINPUT54), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n652), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n676), .B(new_n843), .C1(new_n675), .C2(KEYINPUT10), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n674), .A3(KEYINPUT54), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n844), .A2(new_n674), .A3(KEYINPUT54), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n841), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n604), .A2(new_n846), .A3(new_n849), .A4(new_n684), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n584), .A2(new_n585), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n591), .A2(new_n592), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n598), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n685), .A2(new_n602), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n783), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n846), .A2(new_n849), .A3(new_n684), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n602), .A2(new_n853), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n856), .A2(new_n666), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n722), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n686), .A2(new_n725), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n775), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n531), .A2(new_n536), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n861), .A2(new_n427), .A3(new_n425), .A4(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n334), .A3(new_n725), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n536), .B1(new_n859), .B2(new_n860), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n700), .A2(new_n775), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(new_n535), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n604), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n864), .B1(new_n869), .B2(new_n334), .ZN(G1340gat));
  NAND2_X1  g669(.A1(new_n685), .A2(new_n336), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT120), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G120gat), .B1(new_n863), .B2(new_n723), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1341gat));
  NAND3_X1  g674(.A1(new_n868), .A2(new_n326), .A3(new_n635), .ZN(new_n876));
  OAI21_X1  g675(.A(G127gat), .B1(new_n863), .B2(new_n722), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1342gat));
  NOR2_X1   g677(.A1(new_n666), .A2(new_n531), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT121), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n867), .A2(new_n324), .A3(new_n881), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n863), .B2(new_n666), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G1343gat));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n463), .B1(new_n859), .B2(new_n860), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n698), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI211_X1 g690(.A(KEYINPUT57), .B(new_n463), .C1(new_n859), .C2(new_n860), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n891), .A2(new_n604), .A3(new_n862), .A4(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n745), .A2(new_n463), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n865), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n725), .A2(G141gat), .A3(new_n531), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n894), .A2(G141gat), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n894), .A2(G141gat), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n725), .A2(G141gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n865), .A2(KEYINPUT122), .A3(new_n895), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n902), .A2(new_n535), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n887), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n887), .A2(new_n899), .B1(new_n900), .B2(new_n906), .ZN(G1344gat));
  NOR2_X1   g706(.A1(new_n723), .A2(G148gat), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n902), .A2(new_n535), .A3(new_n904), .A4(new_n908), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n685), .A3(new_n862), .A4(new_n893), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n910), .A2(new_n911), .A3(G148gat), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n910), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(G1345gat));
  NOR2_X1   g713(.A1(new_n722), .A2(G155gat), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n902), .A2(new_n535), .A3(new_n904), .A4(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n862), .ZN(new_n917));
  NOR4_X1   g716(.A1(new_n890), .A2(new_n892), .A3(new_n722), .A4(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n918), .B2(new_n304), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT123), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(new_n916), .C1(new_n918), .C2(new_n304), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1346gat));
  NAND2_X1  g722(.A1(new_n891), .A2(new_n893), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n666), .A3(new_n917), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n902), .A2(new_n904), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n881), .A2(new_n305), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n925), .A2(new_n305), .B1(new_n926), .B2(new_n927), .ZN(G1347gat));
  AOI21_X1  g727(.A(new_n762), .B1(new_n859), .B2(new_n860), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n866), .A2(new_n531), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT124), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n604), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n762), .A2(new_n535), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n700), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n861), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n217), .A3(new_n725), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n933), .A2(new_n938), .ZN(G1348gat));
  NAND3_X1  g738(.A1(new_n932), .A2(new_n218), .A3(new_n685), .ZN(new_n940));
  OAI21_X1  g739(.A(G176gat), .B1(new_n937), .B2(new_n723), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT125), .ZN(G1349gat));
  NAND4_X1  g742(.A1(new_n929), .A2(new_n246), .A3(new_n635), .A4(new_n931), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(G183gat), .B1(new_n937), .B2(new_n722), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT60), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1350gat));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n209), .A3(new_n783), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n861), .A2(new_n783), .A3(new_n936), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n954), .A2(new_n955), .A3(G190gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n954), .B2(G190gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G1351gat));
  AND3_X1   g757(.A1(new_n929), .A2(new_n531), .A3(new_n895), .ZN(new_n959));
  AOI21_X1  g758(.A(G197gat), .B1(new_n959), .B2(new_n604), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n924), .A2(new_n935), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n725), .A2(new_n265), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G1352gat));
  NAND3_X1  g762(.A1(new_n959), .A2(new_n266), .A3(new_n685), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n924), .A2(new_n723), .A3(new_n935), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n965), .B(new_n966), .C1(new_n967), .C2(new_n266), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n959), .A2(new_n259), .A3(new_n635), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n891), .A2(new_n635), .A3(new_n893), .A4(new_n934), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  NAND3_X1  g772(.A1(new_n959), .A2(new_n260), .A3(new_n783), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n924), .A2(new_n666), .A3(new_n935), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(new_n260), .ZN(G1355gat));
endmodule


