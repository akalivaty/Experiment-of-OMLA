//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999;
  INV_X1    g000(.A(KEYINPUT24), .ZN(new_n202));
  NAND3_X1  g001(.A1(new_n202), .A2(G183gat), .A3(G190gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G183gat), .B(G190gat), .ZN(new_n204));
  OAI211_X1 g003(.A(KEYINPUT65), .B(new_n203), .C1(new_n204), .C2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT25), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n204), .B2(new_n202), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n213), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n202), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G190gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n215), .B1(new_n220), .B2(KEYINPUT24), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n221), .B(new_n222), .C1(KEYINPUT65), .C2(KEYINPUT25), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G134gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G127gat), .ZN(new_n226));
  INV_X1    g025(.A(G127gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G134gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G113gat), .B2(G120gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G120gat), .ZN(new_n236));
  INV_X1    g035(.A(G113gat), .ZN(new_n237));
  INV_X1    g036(.A(G120gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT1), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(new_n237), .B2(new_n238), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n232), .A2(new_n236), .B1(new_n240), .B2(new_n229), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT27), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G183gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n244), .A3(new_n218), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n216), .B2(new_n218), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n212), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n241), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n224), .A2(new_n252), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n231), .B1(G113gat), .B2(G120gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G127gat), .B(G134gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n239), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n238), .B1(new_n233), .B2(new_n234), .ZN(new_n260));
  OAI22_X1  g059(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n263), .B(KEYINPUT64), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n214), .A2(new_n223), .B1(new_n247), .B2(new_n251), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT67), .A3(new_n241), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n255), .A2(new_n262), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT34), .B1(new_n268), .B2(KEYINPUT71), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT32), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n267), .A3(new_n262), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n274), .B2(new_n264), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT68), .B(KEYINPUT33), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n277), .B1(new_n274), .B2(new_n264), .ZN(new_n278));
  XOR2_X1   g077(.A(G15gat), .B(G43gat), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT69), .ZN(new_n280));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n275), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n276), .B1(new_n283), .B2(KEYINPUT70), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(KEYINPUT70), .B2(new_n283), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n275), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n272), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n275), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n264), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n276), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n292), .A3(new_n282), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n268), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(new_n269), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n295), .A3(new_n287), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n289), .A2(KEYINPUT72), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n298), .B(new_n272), .C1(new_n284), .C2(new_n288), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G78gat), .B(G106gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT31), .B(G50gat), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n301), .B(new_n302), .Z(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G228gat), .A2(G233gat), .ZN(new_n305));
  AND2_X1   g104(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n307));
  OAI21_X1  g106(.A(G218gat), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(G197gat), .B(G204gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G218gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G211gat), .ZN(new_n316));
  INV_X1    g115(.A(G211gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G218gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n311), .A2(KEYINPUT75), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT73), .B(G211gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT22), .B1(new_n325), .B2(G218gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n312), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n326), .A2(KEYINPUT74), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n310), .B2(new_n312), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n324), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT74), .B1(new_n326), .B2(new_n327), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n310), .A2(new_n329), .A3(new_n312), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(KEYINPUT76), .A3(new_n324), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n314), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339));
  NAND2_X1  g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT2), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G155gat), .B(G162gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G141gat), .B(G148gat), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n340), .A2(KEYINPUT2), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G141gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G148gat), .ZN(new_n349));
  INV_X1    g148(.A(G148gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n341), .B(new_n352), .C1(new_n355), .C2(new_n342), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n339), .B1(new_n358), .B2(KEYINPUT3), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n305), .B1(new_n338), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT76), .B1(new_n336), .B2(new_n324), .ZN(new_n361));
  AOI211_X1 g160(.A(new_n332), .B(new_n323), .C1(new_n334), .C2(new_n335), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n313), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT3), .B1(new_n363), .B2(new_n339), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n360), .B1(new_n364), .B2(new_n357), .ZN(new_n365));
  INV_X1    g164(.A(G22gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n368));
  OR2_X1    g167(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n315), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n312), .B1(new_n371), .B2(KEYINPUT22), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n313), .A2(new_n368), .B1(new_n372), .B2(new_n319), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n310), .A2(KEYINPUT82), .A3(new_n311), .A4(new_n312), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n367), .B(new_n358), .C1(new_n375), .C2(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n319), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n311), .A2(new_n312), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n368), .B1(new_n326), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n379), .A3(new_n374), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT3), .B1(new_n380), .B2(new_n339), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT83), .B1(new_n381), .B2(new_n357), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n313), .B(new_n359), .C1(new_n361), .C2(new_n362), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n376), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n305), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n366), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n304), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n365), .A2(new_n366), .A3(new_n385), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n366), .B1(new_n365), .B2(new_n385), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT85), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n384), .A2(new_n305), .ZN(new_n394));
  INV_X1    g193(.A(new_n305), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n383), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n396), .B1(new_n398), .B2(new_n358), .ZN(new_n399));
  OAI21_X1  g198(.A(G22gat), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n393), .B1(new_n400), .B2(new_n386), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n389), .B1(new_n392), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT0), .ZN(new_n404));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT81), .B1(new_n241), .B2(new_n357), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n261), .A2(new_n410), .A3(new_n356), .A4(new_n347), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n241), .A2(new_n357), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT79), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n241), .A2(new_n357), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n408), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT5), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n347), .A2(new_n356), .A3(KEYINPUT3), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT78), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n347), .A2(new_n356), .A3(KEYINPUT78), .A4(KEYINPUT3), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n241), .B1(new_n397), .B2(new_n357), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n408), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n414), .A2(new_n427), .A3(new_n416), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n427), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT80), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n241), .A2(new_n357), .A3(new_n415), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n415), .B1(new_n241), .B2(new_n357), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n429), .B1(new_n436), .B2(new_n427), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(KEYINPUT80), .A3(new_n426), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n419), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n413), .A2(new_n427), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(new_n417), .B2(KEYINPUT4), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT5), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n426), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n407), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n409), .A2(new_n411), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n443), .B1(new_n448), .B2(new_n408), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT80), .B1(new_n437), .B2(new_n426), .ZN(new_n450));
  AND4_X1   g249(.A1(KEYINPUT80), .A2(new_n426), .A3(new_n428), .A4(new_n430), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(new_n406), .A3(new_n444), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n446), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(KEYINPUT6), .B(new_n407), .C1(new_n439), .C2(new_n445), .ZN(new_n456));
  AND2_X1   g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n256), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n266), .A2(KEYINPUT29), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n363), .B(new_n458), .C1(new_n459), .C2(new_n457), .ZN(new_n460));
  INV_X1    g259(.A(new_n458), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n457), .B1(new_n256), .B2(new_n339), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n338), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465));
  XNOR2_X1  g264(.A(G8gat), .B(G36gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(G64gat), .B(G92gat), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n466), .B(new_n467), .Z(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n460), .A2(new_n463), .ZN(new_n470));
  INV_X1    g269(.A(new_n468), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n460), .A2(new_n463), .A3(new_n468), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(KEYINPUT30), .A3(new_n473), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n455), .A2(new_n456), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT85), .B1(new_n390), .B2(new_n391), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n400), .A2(new_n393), .A3(new_n386), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n388), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n300), .A2(new_n402), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT90), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n482), .A3(KEYINPUT35), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT35), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n289), .A2(new_n484), .A3(new_n296), .ZN(new_n485));
  AND4_X1   g284(.A1(new_n475), .A2(new_n402), .A3(new_n478), .A4(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n481), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n476), .A2(new_n388), .A3(new_n477), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n388), .B1(new_n476), .B2(new_n477), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT86), .B1(new_n402), .B2(new_n478), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n455), .A2(new_n456), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n469), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OAI22_X1  g296(.A1(new_n492), .A2(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT36), .B1(new_n289), .B2(new_n296), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n300), .B2(KEYINPUT36), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n424), .A2(new_n425), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n440), .C1(new_n436), .C2(new_n427), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT39), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n408), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n502), .A2(new_n408), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT39), .B1(new_n448), .B2(new_n408), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n406), .B(new_n504), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n502), .A2(new_n408), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n510), .B(KEYINPUT39), .C1(new_n408), .C2(new_n448), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(KEYINPUT40), .A3(new_n406), .A4(new_n504), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n446), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(new_n496), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n489), .A2(new_n490), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n464), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT88), .B1(new_n470), .B2(KEYINPUT37), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n468), .B1(new_n470), .B2(KEYINPUT37), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT89), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n521), .A2(KEYINPUT89), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT38), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n463), .A2(KEYINPUT87), .A3(new_n363), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(new_n517), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n464), .A2(KEYINPUT87), .ZN(new_n528));
  AOI211_X1 g327(.A(KEYINPUT38), .B(new_n468), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n520), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n495), .A2(new_n525), .A3(new_n530), .A4(new_n473), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n500), .B1(new_n515), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n498), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n488), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT93), .B(G43gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n537));
  INV_X1    g336(.A(G50gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT94), .B1(new_n535), .B2(G50gat), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n538), .A2(G43gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT15), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(KEYINPUT95), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(KEYINPUT95), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n538), .A2(G43gat), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n541), .A2(KEYINPUT15), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G29gat), .ZN(new_n551));
  INV_X1    g350(.A(G36gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT14), .ZN(new_n554));
  NAND2_X1  g353(.A1(G29gat), .A2(G36gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT96), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n550), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n549), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT92), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n559), .A2(KEYINPUT17), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n557), .B1(new_n545), .B2(new_n546), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(new_n562), .ZN(new_n567));
  XNOR2_X1  g366(.A(G15gat), .B(G22gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT16), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(G1gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(G1gat), .B2(new_n568), .ZN(new_n571));
  INV_X1    g370(.A(G8gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n564), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n563), .ZN(new_n576));
  INV_X1    g375(.A(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT18), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n574), .A2(KEYINPUT18), .A3(new_n575), .A4(new_n578), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n559), .A2(new_n563), .A3(new_n573), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n575), .B(KEYINPUT13), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G169gat), .B(G197gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT12), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n581), .A2(new_n582), .A3(new_n586), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n534), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT97), .Z(new_n602));
  NAND2_X1  g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT9), .ZN(new_n604));
  XNOR2_X1  g403(.A(G57gat), .B(G64gat), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n603), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n605), .B1(new_n604), .B2(new_n603), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n609), .A2(KEYINPUT99), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT99), .B1(new_n609), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n573), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT101), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n614), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT100), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n623), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n617), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n617), .A2(new_n624), .A3(new_n625), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  INV_X1    g432(.A(new_n631), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n626), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(KEYINPUT41), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G134gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G162gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(G85gat), .A2(G92gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT7), .ZN(new_n643));
  NAND2_X1  g442(.A1(G99gat), .A2(G106gat), .ZN(new_n644));
  INV_X1    g443(.A(G85gat), .ZN(new_n645));
  INV_X1    g444(.A(G92gat), .ZN(new_n646));
  AOI22_X1  g445(.A1(KEYINPUT8), .A2(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G99gat), .B(G106gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT102), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n643), .A2(new_n652), .A3(new_n649), .A4(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n576), .A2(new_n654), .B1(KEYINPUT41), .B2(new_n638), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n564), .A2(new_n567), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G190gat), .B(G218gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT103), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n641), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n658), .A2(new_n661), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n660), .B1(new_n655), .B2(new_n657), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(KEYINPUT104), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n669), .A2(new_n641), .B1(new_n665), .B2(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G120gat), .B(G148gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(G176gat), .B(G204gat), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(G230gat), .A2(G233gat), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n654), .A2(new_n613), .ZN(new_n678));
  INV_X1    g477(.A(new_n650), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n679), .B(new_n606), .C1(new_n611), .C2(new_n612), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT10), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR3_X1    g482(.A1(new_n656), .A2(new_n682), .A3(new_n613), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n677), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n678), .A2(new_n677), .A3(new_n680), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n675), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT10), .B1(new_n678), .B2(new_n680), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n656), .A2(new_n682), .A3(new_n613), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n676), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(new_n686), .A3(new_n674), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n637), .A2(new_n671), .A3(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n598), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n494), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT105), .B(G1gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1324gat));
  INV_X1    g498(.A(new_n696), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n572), .B1(new_n700), .B2(new_n497), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT16), .B(G8gat), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n696), .A2(new_n496), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT42), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(KEYINPUT42), .B2(new_n703), .ZN(G1325gat));
  INV_X1    g504(.A(G15gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n289), .A2(new_n296), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n696), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT106), .ZN(new_n709));
  INV_X1    g508(.A(new_n500), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n696), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n709), .A2(new_n711), .ZN(G1326gat));
  NOR2_X1   g511(.A1(new_n492), .A2(new_n493), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n696), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  AND2_X1   g515(.A1(new_n668), .A2(new_n670), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n693), .B1(new_n632), .B2(new_n635), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT107), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n534), .A2(new_n597), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n551), .A3(new_n495), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT45), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n486), .B1(new_n480), .B2(KEYINPUT90), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n725), .A2(new_n483), .B1(new_n498), .B2(new_n532), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n726), .B2(new_n671), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n479), .A2(new_n482), .A3(KEYINPUT35), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n482), .B1(new_n479), .B2(KEYINPUT35), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n728), .A2(new_n729), .A3(new_n486), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n498), .A2(new_n532), .ZN(new_n731));
  OAI211_X1 g530(.A(KEYINPUT44), .B(new_n717), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n718), .A2(new_n597), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G29gat), .B1(new_n735), .B2(new_n494), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n723), .A2(new_n736), .ZN(G1328gat));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n552), .A3(new_n497), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT46), .Z(new_n739));
  OAI21_X1  g538(.A(G36gat), .B1(new_n735), .B2(new_n496), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(G1329gat));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(KEYINPUT109), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n707), .A2(new_n536), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n534), .A2(new_n597), .A3(new_n720), .A4(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n727), .A2(new_n500), .A3(new_n732), .A4(new_n734), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n536), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n743), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n742), .A2(KEYINPUT109), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1330gat));
  NOR2_X1   g551(.A1(new_n713), .A2(G50gat), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n534), .A2(new_n597), .A3(new_n720), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT48), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n489), .A2(new_n490), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n727), .A2(new_n757), .A3(new_n732), .A4(new_n734), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(G50gat), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  INV_X1    g561(.A(new_n713), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n733), .A2(new_n763), .A3(new_n734), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n764), .A2(G50gat), .B1(new_n721), .B2(new_n753), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n761), .A2(new_n762), .B1(new_n765), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g565(.A1(new_n717), .A2(new_n636), .A3(new_n597), .A4(new_n694), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n534), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n495), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g570(.A1(new_n768), .A2(new_n496), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  AND2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n772), .B2(new_n773), .ZN(G1333gat));
  AOI21_X1  g575(.A(new_n599), .B1(new_n769), .B2(new_n500), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n768), .A2(G71gat), .A3(new_n707), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n768), .A2(new_n713), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(new_n600), .ZN(G1335gat));
  INV_X1    g581(.A(new_n596), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n579), .A2(new_n580), .B1(new_n584), .B2(new_n585), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n595), .B1(new_n784), .B2(new_n582), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n636), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT111), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n694), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n733), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n494), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  NOR4_X1   g591(.A1(new_n726), .A2(new_n792), .A3(new_n788), .A4(new_n671), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n671), .B1(new_n488), .B2(new_n533), .ZN(new_n794));
  INV_X1    g593(.A(new_n788), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT51), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n495), .A2(new_n645), .A3(new_n693), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n791), .B1(new_n797), .B2(new_n798), .ZN(G1336gat));
  NAND4_X1  g598(.A1(new_n727), .A2(new_n497), .A3(new_n732), .A4(new_n789), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G92gat), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n694), .A2(G92gat), .A3(new_n496), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT113), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n801), .A2(KEYINPUT112), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n794), .A2(new_n795), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n792), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n794), .A2(KEYINPUT51), .A3(new_n795), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n802), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(new_n801), .C1(KEYINPUT112), .C2(new_n810), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n805), .A2(new_n812), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n790), .B2(new_n710), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n694), .A2(new_n707), .A3(G99gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n797), .B2(new_n815), .ZN(G1338gat));
  NAND4_X1  g615(.A1(new_n727), .A2(new_n757), .A3(new_n732), .A4(new_n789), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G106gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n756), .A2(G106gat), .A3(new_n694), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n793), .B2(new_n796), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n727), .A2(new_n763), .A3(new_n732), .A4(new_n789), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n821), .B1(new_n824), .B2(new_n820), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT114), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n809), .A2(new_n819), .B1(G106gat), .B2(new_n823), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n821), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n830), .ZN(G1339gat));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n683), .A2(new_n684), .A3(new_n677), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n833), .A2(KEYINPUT54), .A3(new_n691), .ZN(new_n834));
  XOR2_X1   g633(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n675), .B1(new_n691), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n832), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n674), .B1(new_n685), .B2(new_n835), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n691), .A3(KEYINPUT54), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n838), .A2(new_n692), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n584), .A2(new_n585), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n575), .B1(new_n574), .B2(new_n578), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n592), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n596), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n717), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n597), .A2(new_n842), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n596), .A2(new_n693), .A3(new_n845), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n717), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n636), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n695), .A2(new_n597), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n763), .A2(new_n707), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n494), .A2(new_n497), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n786), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n494), .B1(new_n853), .B2(new_n855), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n756), .A2(new_n496), .A3(new_n300), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n597), .A2(new_n233), .A3(new_n234), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(G1340gat));
  INV_X1    g665(.A(new_n864), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n238), .A3(new_n693), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n856), .A2(new_n693), .A3(new_n859), .A4(new_n857), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n869), .A2(new_n870), .A3(G120gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n869), .B2(G120gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT117), .ZN(G1341gat));
  OAI21_X1  g673(.A(G127gat), .B1(new_n860), .B2(new_n636), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n867), .A2(new_n227), .A3(new_n637), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1342gat));
  NAND3_X1  g676(.A1(new_n867), .A2(new_n225), .A3(new_n717), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n860), .B2(new_n671), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n710), .A2(new_n859), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n756), .B1(new_n853), .B2(new_n855), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n841), .A2(new_n692), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n839), .A2(new_n840), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n832), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n887), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n850), .B1(new_n892), .B2(new_n597), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(new_n893), .B2(new_n717), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n841), .A2(new_n692), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n890), .B1(new_n889), .B2(new_n832), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT118), .B(KEYINPUT55), .C1(new_n839), .C2(new_n840), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n851), .B1(new_n898), .B2(new_n786), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n671), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n894), .A2(new_n901), .A3(new_n847), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n636), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n713), .B1(new_n903), .B2(new_n855), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n597), .B(new_n886), .C1(new_n904), .C2(new_n885), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G141gat), .ZN(new_n906));
  AND4_X1   g705(.A1(new_n496), .A2(new_n862), .A3(new_n757), .A4(new_n710), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n348), .A3(new_n597), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g708(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n910), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n906), .A2(new_n912), .A3(new_n908), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n907), .A2(new_n350), .A3(new_n693), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n713), .A2(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n847), .B1(new_n893), .B2(new_n717), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n918), .A2(KEYINPUT121), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n637), .B1(new_n918), .B2(KEYINPUT121), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n921), .B2(new_n854), .ZN(new_n922));
  INV_X1    g721(.A(new_n883), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n856), .A2(new_n757), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT57), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n922), .A2(new_n693), .A3(new_n923), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n916), .B1(new_n926), .B2(G148gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n916), .A2(G148gat), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n904), .A2(new_n885), .ZN(new_n929));
  INV_X1    g728(.A(new_n886), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(new_n693), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n915), .B1(new_n927), .B2(new_n932), .ZN(G1345gat));
  OAI211_X1 g732(.A(new_n637), .B(new_n886), .C1(new_n904), .C2(new_n885), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G155gat), .ZN(new_n935));
  INV_X1    g734(.A(G155gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n907), .A2(new_n936), .A3(new_n637), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT122), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n935), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1346gat));
  AOI21_X1  g741(.A(G162gat), .B1(new_n907), .B2(new_n717), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n717), .A2(G162gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n931), .B2(new_n944), .ZN(G1347gat));
  AOI21_X1  g744(.A(new_n495), .B1(new_n853), .B2(new_n855), .ZN(new_n946));
  AND4_X1   g745(.A1(new_n497), .A2(new_n946), .A3(new_n756), .A4(new_n300), .ZN(new_n947));
  INV_X1    g746(.A(G169gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n947), .A2(new_n948), .A3(new_n597), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n494), .A2(new_n497), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n858), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n597), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT124), .B1(new_n954), .B2(G169gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(G1348gat));
  OAI21_X1  g756(.A(G176gat), .B1(new_n952), .B2(new_n694), .ZN(new_n958));
  INV_X1    g757(.A(G176gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n947), .A2(new_n959), .A3(new_n693), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT125), .ZN(G1349gat));
  NAND4_X1  g761(.A1(new_n947), .A2(new_n242), .A3(new_n244), .A4(new_n637), .ZN(new_n963));
  OAI21_X1  g762(.A(G183gat), .B1(new_n952), .B2(new_n636), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n947), .A2(new_n218), .A3(new_n717), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n717), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(G190gat), .ZN(new_n970));
  AOI211_X1 g769(.A(KEYINPUT61), .B(new_n218), .C1(new_n953), .C2(new_n717), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(G1351gat));
  AND4_X1   g771(.A1(new_n497), .A2(new_n946), .A3(new_n757), .A4(new_n710), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n597), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n951), .A2(new_n710), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n854), .B1(new_n919), .B2(new_n920), .ZN(new_n977));
  INV_X1    g776(.A(new_n917), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n925), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n597), .A2(G197gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n974), .B1(new_n980), .B2(new_n981), .ZN(G1352gat));
  XNOR2_X1  g781(.A(KEYINPUT126), .B(G204gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n694), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n973), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n985), .B(KEYINPUT62), .Z(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n979), .B2(new_n694), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1353gat));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n369), .A3(new_n370), .A4(new_n637), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT63), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n990), .A2(KEYINPUT127), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n317), .B1(KEYINPUT127), .B2(new_n990), .ZN(new_n992));
  OAI211_X1 g791(.A(new_n991), .B(new_n992), .C1(new_n979), .C2(new_n636), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n922), .A2(new_n637), .A3(new_n925), .A4(new_n976), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n991), .B1(new_n995), .B2(new_n992), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n989), .B1(new_n994), .B2(new_n996), .ZN(G1354gat));
  OAI21_X1  g796(.A(G218gat), .B1(new_n979), .B2(new_n671), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n973), .A2(new_n315), .A3(new_n717), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1355gat));
endmodule


