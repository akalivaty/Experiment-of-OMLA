//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT80), .Z(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT70), .B(G953), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XOR2_X1   g008(.A(G110), .B(G140), .Z(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT0), .B(G128), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n211), .A2(KEYINPUT3), .A3(G107), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT81), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT81), .A2(G104), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(G107), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(G107), .B1(new_n215), .B2(new_n216), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n213), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT84), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT84), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n220), .A2(new_n224), .A3(new_n221), .A4(G101), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n210), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n221), .B1(new_n220), .B2(G101), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT83), .ZN(new_n228));
  INV_X1    g042(.A(G107), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT81), .A2(G104), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT81), .A2(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n212), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT82), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n230), .A2(new_n231), .ZN(new_n235));
  AOI21_X1  g049(.A(G101), .B1(new_n235), .B2(G107), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n233), .B2(new_n236), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n227), .B(new_n228), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n213), .B1(new_n218), .B2(new_n219), .ZN(new_n241));
  INV_X1    g055(.A(G101), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n217), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT82), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n228), .B1(new_n246), .B2(new_n227), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n226), .B1(new_n240), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n250), .B(new_n205), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT10), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT85), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n211), .A2(G107), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n242), .B1(new_n232), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n254), .B1(new_n246), .B2(new_n257), .ZN(new_n258));
  AOI211_X1 g072(.A(KEYINPUT85), .B(new_n256), .C1(new_n244), .C2(new_n245), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT11), .A3(G134), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G137), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT11), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n263), .B2(G137), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n265), .A2(KEYINPUT65), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n268), .A2(new_n262), .A3(new_n266), .A4(new_n264), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n264), .A3(new_n262), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n269), .A2(new_n272), .B1(G131), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n256), .B1(new_n244), .B2(new_n245), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n250), .B(new_n199), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n252), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n248), .A2(new_n260), .A3(new_n274), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n257), .B1(new_n237), .B2(new_n238), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT85), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n254), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n251), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n277), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n273), .A2(G131), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n270), .A2(new_n271), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n270), .A2(new_n271), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n280), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(KEYINPUT12), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n274), .B(new_n292), .C1(new_n284), .C2(new_n277), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n197), .B(new_n279), .C1(new_n290), .C2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n227), .B1(new_n237), .B2(new_n238), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT83), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n239), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n297), .A2(new_n226), .B1(new_n252), .B2(new_n277), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n274), .B1(new_n298), .B2(new_n260), .ZN(new_n299));
  AND4_X1   g113(.A1(new_n274), .A2(new_n248), .A3(new_n260), .A4(new_n278), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n196), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n192), .B1(new_n302), .B2(new_n190), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n248), .A2(new_n260), .A3(new_n278), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n289), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n197), .A3(new_n279), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n285), .A2(new_n289), .ZN(new_n307));
  INV_X1    g121(.A(new_n280), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n285), .B(new_n289), .C1(new_n291), .C2(KEYINPUT12), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n300), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(G469), .B(new_n306), .C1(new_n311), .C2(new_n197), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n189), .B1(new_n303), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n314));
  INV_X1    g128(.A(G110), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n249), .A2(G119), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n249), .A2(KEYINPUT23), .A3(G119), .ZN(new_n319));
  INV_X1    g133(.A(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G128), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n315), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n323), .B2(new_n322), .ZN(new_n325));
  XNOR2_X1  g139(.A(G125), .B(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(G146), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G146), .B1(new_n327), .B2(new_n329), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n316), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT24), .B(G110), .ZN(new_n334));
  OAI221_X1 g148(.A(new_n325), .B1(new_n331), .B2(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n326), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n330), .B1(G146), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n333), .A2(new_n334), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n318), .A2(new_n319), .A3(new_n315), .A4(new_n321), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT77), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n340), .A2(KEYINPUT78), .A3(new_n341), .A4(new_n342), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n337), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI211_X1 g163(.A(KEYINPUT79), .B(new_n337), .C1(new_n345), .C2(new_n346), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n335), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G137), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n335), .B(new_n354), .C1(new_n349), .C2(new_n350), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n314), .B1(new_n358), .B2(G902), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n356), .A2(KEYINPUT25), .A3(new_n191), .A4(new_n357), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G217), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(G234), .B2(new_n191), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(G902), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n356), .A2(new_n357), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G472), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT68), .B1(new_n274), .B2(new_n210), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n289), .A2(new_n371), .A3(new_n209), .ZN(new_n372));
  INV_X1    g186(.A(G113), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT2), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT2), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G113), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G116), .B(G119), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT67), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT67), .B1(new_n377), .B2(new_n378), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n261), .A2(G134), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n266), .B1(new_n383), .B2(new_n264), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n269), .B2(new_n272), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n382), .B1(new_n385), .B2(new_n276), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n370), .A2(new_n372), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT69), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT69), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n370), .A2(new_n372), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n385), .A2(new_n276), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n370), .A2(new_n372), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n382), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT74), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(KEYINPUT74), .A3(new_n382), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT28), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n274), .A2(new_n210), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT28), .B1(new_n401), .B2(new_n386), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G237), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n193), .A2(G210), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT72), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(G101), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n406), .B(new_n409), .Z(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT29), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n399), .A2(new_n403), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n191), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n370), .A2(new_n372), .A3(KEYINPUT30), .A4(new_n392), .ZN(new_n417));
  INV_X1    g231(.A(new_n384), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n287), .B2(new_n288), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT66), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n251), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n385), .A2(KEYINPUT66), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n400), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n382), .B(new_n417), .C1(new_n423), .C2(KEYINPUT30), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n410), .B1(new_n424), .B2(new_n391), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT73), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n422), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n401), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n382), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n391), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n402), .B1(new_n430), .B2(KEYINPUT28), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT29), .B1(new_n431), .B2(new_n410), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n415), .A2(new_n416), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n402), .B1(new_n398), .B2(KEYINPUT28), .ZN(new_n434));
  AOI211_X1 g248(.A(new_n416), .B(G902), .C1(new_n434), .C2(new_n413), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n369), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n424), .A2(new_n391), .A3(new_n410), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT31), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT31), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n424), .A2(new_n391), .A3(new_n440), .A4(new_n410), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n439), .B(new_n441), .C1(new_n431), .C2(new_n410), .ZN(new_n442));
  NOR2_X1   g256(.A1(G472), .A2(G902), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT32), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n442), .A2(KEYINPUT32), .A3(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n313), .B(new_n368), .C1(new_n437), .C2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n450));
  MUX2_X1   g264(.A(new_n251), .B(new_n210), .S(G125), .Z(new_n451));
  INV_X1    g265(.A(G224), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n451), .B(new_n453), .Z(new_n454));
  NAND2_X1  g268(.A1(new_n377), .A2(new_n378), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT67), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n223), .A2(new_n225), .B1(new_n379), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n240), .B2(new_n247), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n378), .A2(KEYINPUT5), .ZN(new_n462));
  INV_X1    g276(.A(G116), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n463), .A2(KEYINPUT5), .A3(G119), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(new_n373), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n258), .B2(new_n259), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G122), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n461), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT87), .A2(KEYINPUT6), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n461), .A2(new_n469), .ZN(new_n475));
  INV_X1    g289(.A(new_n470), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n476), .A3(new_n473), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n454), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n470), .B(KEYINPUT8), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n467), .B1(new_n282), .B2(new_n283), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n275), .A2(new_n468), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT7), .B1(new_n452), .B2(G953), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n451), .B(new_n485), .Z(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n471), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n191), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n450), .B1(new_n480), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n487), .A2(new_n191), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n470), .B(new_n472), .C1(new_n461), .C2(new_n469), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n477), .B2(new_n474), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n490), .B(KEYINPUT88), .C1(new_n492), .C2(new_n454), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n478), .A2(new_n479), .ZN(new_n497));
  INV_X1    g311(.A(new_n454), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n488), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT89), .B1(new_n499), .B2(new_n494), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n193), .A2(G214), .A3(new_n404), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n203), .ZN(new_n504));
  NAND2_X1  g318(.A1(KEYINPUT18), .A2(G131), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT90), .B(G143), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n193), .A2(new_n506), .A3(G214), .A4(new_n404), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n505), .B1(new_n504), .B2(new_n507), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n326), .B(G146), .ZN(new_n510));
  OR3_X1    g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G113), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n211), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n504), .A2(new_n507), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G131), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n504), .A2(new_n266), .A3(new_n507), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n332), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n330), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT91), .B1(new_n331), .B2(new_n332), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n521), .B(new_n522), .C1(new_n515), .C2(new_n516), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n511), .B(new_n513), .C1(new_n518), .C2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n513), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n326), .B(KEYINPUT19), .Z(new_n526));
  OAI21_X1  g340(.A(new_n330), .B1(new_n526), .B2(G146), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n515), .B2(new_n517), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(G475), .A2(G902), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT20), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT20), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT92), .ZN(new_n538));
  INV_X1    g352(.A(G122), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G116), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n463), .A2(G122), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n229), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n203), .A2(G128), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n249), .A2(G143), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n544), .A2(new_n545), .ZN(new_n549));
  OAI21_X1  g363(.A(G134), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n544), .A2(new_n547), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n263), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n543), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n551), .B(new_n263), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n542), .A2(new_n229), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n541), .A2(KEYINPUT14), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n541), .A2(KEYINPUT14), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n540), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G107), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n538), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n187), .A2(new_n362), .A3(G953), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n560), .A3(new_n538), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n563), .ZN(new_n566));
  INV_X1    g380(.A(new_n564), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(new_n561), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n568), .A3(new_n191), .ZN(new_n569));
  INV_X1    g383(.A(G478), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT15), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n569), .B(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n511), .B1(new_n518), .B2(new_n523), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n525), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n524), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n191), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G475), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n537), .A2(new_n573), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G952), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G953), .ZN(new_n581));
  INV_X1    g395(.A(G234), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n404), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n193), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(G902), .C1(new_n582), .C2(new_n404), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT93), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT21), .B(G898), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT94), .B1(new_n579), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n535), .B1(new_n531), .B2(new_n532), .ZN(new_n592));
  INV_X1    g406(.A(new_n532), .ZN(new_n593));
  AOI211_X1 g407(.A(KEYINPUT20), .B(new_n593), .C1(new_n524), .C2(new_n530), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n575), .B2(new_n524), .ZN(new_n595));
  INV_X1    g409(.A(G475), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n592), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n599));
  INV_X1    g413(.A(new_n590), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n573), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n591), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G214), .B1(G237), .B2(G902), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n489), .A2(KEYINPUT89), .A3(new_n493), .A4(new_n495), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n501), .A2(new_n602), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n449), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n242), .ZN(G3));
  OAI21_X1  g421(.A(KEYINPUT95), .B1(new_n499), .B2(new_n494), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n490), .B(new_n494), .C1(new_n492), .C2(new_n454), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n610), .B(new_n495), .C1(new_n480), .C2(new_n488), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n567), .A2(new_n566), .A3(new_n561), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n565), .A2(new_n568), .A3(KEYINPUT33), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n570), .A2(G902), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n569), .A2(new_n570), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n597), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n590), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n612), .A2(new_n603), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n444), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n369), .B1(new_n442), .B2(new_n191), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n189), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n279), .A2(new_n197), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n309), .B2(new_n310), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n197), .B1(new_n305), .B2(new_n279), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n190), .B(new_n191), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n633), .B(new_n312), .C1(new_n190), .C2(new_n191), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n628), .A2(new_n368), .A3(new_n629), .A4(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n625), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT34), .B(G104), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  NAND3_X1  g452(.A1(new_n534), .A2(KEYINPUT96), .A3(new_n536), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n592), .B2(new_n594), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n573), .ZN(new_n643));
  AND4_X1   g457(.A1(new_n600), .A2(new_n642), .A3(new_n578), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n612), .A2(new_n603), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n635), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT35), .B(G107), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  INV_X1    g462(.A(new_n363), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n359), .B2(new_n360), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n355), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT97), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(new_n351), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n351), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n655), .A2(G902), .A3(new_n363), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n313), .A2(new_n628), .A3(new_n658), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n605), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n424), .A2(new_n391), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n411), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT73), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT73), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n425), .A2(new_n666), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n390), .A2(new_n388), .B1(new_n428), .B2(new_n382), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT28), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n410), .B(new_n403), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n665), .A2(new_n412), .A3(new_n667), .A4(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(G902), .B1(new_n434), .B2(new_n413), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n671), .B1(new_n672), .B2(KEYINPUT75), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n673), .B2(new_n435), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n442), .A2(KEYINPUT32), .A3(new_n443), .ZN(new_n675));
  AOI21_X1  g489(.A(KEYINPUT32), .B1(new_n442), .B2(new_n443), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n657), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n611), .A2(new_n609), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n490), .B1(new_n492), .B2(new_n454), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n610), .B1(new_n680), .B2(new_n495), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n603), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n642), .A2(new_n578), .ZN(new_n684));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n584), .B1(new_n588), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n684), .A2(new_n643), .A3(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n678), .A2(new_n683), .A3(new_n313), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  NAND2_X1  g504(.A1(new_n501), .A2(new_n604), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT38), .ZN(new_n692));
  INV_X1    g506(.A(new_n603), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n598), .A2(new_n693), .A3(new_n573), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n657), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT98), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n686), .B(KEYINPUT39), .Z(new_n697));
  NAND2_X1  g511(.A1(new_n313), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n663), .A2(new_n410), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n700), .B(new_n191), .C1(new_n410), .C2(new_n398), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G472), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n446), .A2(new_n447), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n696), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n692), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n203), .ZN(G45));
  NOR2_X1   g521(.A1(new_n623), .A2(new_n686), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n603), .B(new_n708), .C1(new_n679), .C2(new_n681), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT99), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n612), .A2(KEYINPUT99), .A3(new_n603), .A4(new_n708), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n313), .A4(new_n678), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  AOI21_X1  g528(.A(new_n367), .B1(new_n674), .B2(new_n677), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n302), .A2(new_n190), .ZN(new_n716));
  AOI211_X1 g530(.A(G469), .B(G902), .C1(new_n294), .C2(new_n301), .ZN(new_n717));
  INV_X1    g531(.A(new_n188), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n625), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT100), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n721), .B(new_n723), .ZN(G15));
  NOR2_X1   g538(.A1(new_n720), .A2(new_n645), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n463), .ZN(G18));
  NAND4_X1  g540(.A1(new_n719), .A2(new_n612), .A3(new_n603), .A4(new_n602), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n658), .B1(new_n437), .B2(new_n448), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT101), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n302), .A2(new_n190), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n188), .A3(new_n633), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n682), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT101), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n602), .A4(new_n678), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n719), .A2(new_n612), .A3(new_n600), .A4(new_n694), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n439), .B1(new_n434), .B2(new_n410), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT102), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(new_n439), .C1(new_n434), .C2(new_n410), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n441), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n627), .B1(new_n743), .B2(new_n443), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n368), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n737), .B1(new_n738), .B2(new_n745), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n627), .B(new_n367), .C1(new_n743), .C2(new_n443), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n731), .A2(new_n590), .ZN(new_n748));
  INV_X1    g562(.A(new_n694), .ZN(new_n749));
  INV_X1    g563(.A(new_n679), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n749), .B1(new_n750), .B2(new_n608), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n747), .A2(new_n748), .A3(new_n751), .A4(KEYINPUT103), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  AOI211_X1 g568(.A(new_n627), .B(new_n657), .C1(new_n743), .C2(new_n443), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n732), .A2(new_n708), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  AOI21_X1  g571(.A(new_n693), .B1(new_n501), .B2(new_n604), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n192), .B(KEYINPUT104), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n302), .B2(new_n190), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n718), .B1(new_n761), .B2(new_n312), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n758), .A2(new_n715), .A3(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n623), .A2(KEYINPUT42), .A3(new_n686), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n758), .A2(new_n708), .A3(new_n762), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n674), .A2(new_n447), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n676), .B(KEYINPUT105), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n368), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT42), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n266), .ZN(G33));
  NAND4_X1  g586(.A1(new_n758), .A2(new_n715), .A3(new_n688), .A4(new_n762), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n598), .A2(new_n622), .A3(new_n775), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n618), .A2(new_n619), .B1(new_n570), .B2(new_n569), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT43), .B1(new_n777), .B2(new_n597), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n776), .B2(new_n778), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n658), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n628), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(KEYINPUT44), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT109), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n783), .A2(new_n787), .A3(KEYINPUT44), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n782), .B2(new_n628), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n758), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n306), .B1(new_n311), .B2(new_n197), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n190), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n796), .B2(new_n795), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT46), .B1(new_n798), .B2(new_n759), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n717), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n759), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n718), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n697), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n697), .ZN(new_n805));
  INV_X1    g619(.A(new_n803), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n794), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(new_n261), .ZN(G39));
  NAND2_X1  g623(.A1(new_n691), .A2(new_n603), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n674), .A2(new_n677), .A3(new_n367), .A4(new_n708), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n802), .A2(KEYINPUT47), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n814), .B(new_n718), .C1(new_n800), .C2(new_n801), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n812), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT110), .B(G140), .Z(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(G42));
  NOR4_X1   g632(.A1(new_n777), .A2(new_n597), .A3(new_n693), .A4(new_n189), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n368), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT111), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n716), .A2(new_n717), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n821), .B1(KEYINPUT49), .B2(new_n823), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT112), .Z(new_n825));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n703), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n692), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT113), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n719), .A2(new_n693), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT117), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n776), .A2(new_n778), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n584), .A2(new_n744), .A3(new_n368), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n692), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT50), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n810), .A2(new_n731), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n703), .A2(new_n583), .A3(new_n367), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n598), .A3(new_n777), .ZN(new_n839));
  INV_X1    g653(.A(new_n755), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n584), .A3(new_n832), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n802), .B(KEYINPUT47), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n823), .A2(new_n629), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n758), .B(new_n833), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT118), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n843), .A2(new_n846), .A3(new_n850), .A4(KEYINPUT51), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n841), .A2(new_n769), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT48), .Z(new_n854));
  NAND2_X1  g668(.A1(new_n833), .A2(new_n732), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n838), .A2(new_n597), .A3(new_n622), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n581), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n847), .B2(new_n848), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n713), .A2(new_n689), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n650), .A2(new_n656), .A3(new_n686), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n762), .A2(new_n703), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n612), .A2(new_n694), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT114), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n633), .A2(new_n312), .A3(new_n759), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n862), .A2(new_n866), .A3(new_n188), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n751), .A2(new_n867), .A3(new_n868), .A4(new_n703), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n861), .A2(KEYINPUT52), .A3(new_n756), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n713), .A2(new_n689), .A3(new_n756), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n865), .A2(new_n869), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n765), .A2(new_n770), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n720), .B1(new_n625), .B2(new_n645), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n777), .A2(new_n597), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n579), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n590), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n501), .A2(new_n603), .A3(new_n881), .A4(new_n604), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n605), .A2(new_n659), .B1(new_n882), .B2(new_n635), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n878), .A2(new_n606), .A3(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n734), .A2(new_n729), .B1(new_n746), .B2(new_n752), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n758), .A2(new_n755), .A3(new_n708), .A4(new_n762), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n684), .A2(new_n573), .A3(new_n687), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n758), .A2(new_n678), .A3(new_n887), .A4(new_n313), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n886), .A2(new_n773), .A3(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n877), .A2(new_n884), .A3(new_n885), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n860), .B1(new_n876), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n770), .A3(new_n765), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n883), .A2(new_n606), .ZN(new_n894));
  INV_X1    g708(.A(new_n625), .ZN(new_n895));
  INV_X1    g709(.A(new_n645), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n715), .B(new_n719), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n894), .A2(new_n735), .A3(new_n753), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n871), .A2(new_n875), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(KEYINPUT53), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n891), .A2(new_n892), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT116), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n891), .A2(new_n904), .A3(new_n892), .A4(new_n901), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n891), .A2(new_n901), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT115), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n903), .A2(new_n908), .A3(KEYINPUT115), .A4(new_n905), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n859), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(G952), .A2(G953), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n829), .B1(new_n912), .B2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n193), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n907), .A2(G210), .A3(G902), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n497), .A2(new_n498), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n480), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT55), .Z(new_n922));
  OAI21_X1  g736(.A(new_n916), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n919), .A2(new_n922), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n919), .A2(KEYINPUT119), .A3(new_n922), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G51));
  AND2_X1   g742(.A1(new_n908), .A2(new_n902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n759), .B(KEYINPUT57), .ZN(new_n930));
  OAI22_X1  g744(.A1(new_n929), .A2(new_n930), .B1(new_n632), .B2(new_n631), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n899), .A2(KEYINPUT53), .A3(new_n900), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT53), .B1(new_n899), .B2(new_n900), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR3_X1    g748(.A1(new_n934), .A2(new_n191), .A3(new_n798), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n915), .B1(new_n931), .B2(new_n935), .ZN(G54));
  NAND4_X1  g750(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n937));
  INV_X1    g751(.A(new_n531), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n915), .ZN(G60));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT59), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n618), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n916), .B1(new_n929), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n910), .A2(new_n911), .A3(new_n944), .ZN(new_n947));
  INV_X1    g761(.A(new_n618), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(G63));
  INV_X1    g763(.A(new_n655), .ZN(new_n950));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  OAI211_X1 g766(.A(new_n950), .B(new_n952), .C1(new_n932), .C2(new_n933), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n952), .B1(new_n932), .B2(new_n933), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n358), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n907), .A2(new_n957), .A3(new_n950), .A4(new_n952), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n954), .A2(new_n956), .A3(new_n958), .A4(new_n916), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT61), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT61), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(G66));
  OAI21_X1  g777(.A(G953), .B1(new_n589), .B2(new_n452), .ZN(new_n964));
  INV_X1    g778(.A(new_n898), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n585), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n492), .B1(G898), .B2(new_n193), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT122), .Z(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(G69));
  OAI21_X1  g783(.A(new_n417), .B1(new_n423), .B2(KEYINPUT30), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(new_n526), .Z(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT123), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n698), .A2(new_n880), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n715), .A3(new_n758), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n816), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n808), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(KEYINPUT62), .B1(new_n706), .B2(new_n873), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n706), .C2(new_n873), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OR3_X1    g795(.A1(new_n706), .A2(KEYINPUT62), .A3(new_n873), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n976), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n972), .B1(new_n983), .B2(new_n585), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n771), .B1(new_n688), .B2(new_n763), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(new_n816), .A3(new_n756), .A4(new_n861), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n769), .A2(new_n864), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AOI22_X1  g802(.A1(new_n794), .A2(new_n988), .B1(new_n807), .B2(new_n804), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT125), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n873), .B1(new_n844), .B2(new_n812), .ZN(new_n991));
  INV_X1    g805(.A(new_n804), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n803), .B1(new_n802), .B2(new_n697), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n792), .B1(new_n786), .B2(new_n788), .ZN(new_n994));
  OAI22_X1  g808(.A1(new_n992), .A2(new_n993), .B1(new_n994), .B2(new_n987), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n991), .A2(new_n995), .A3(new_n996), .A4(new_n985), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n990), .A2(new_n997), .A3(new_n193), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n971), .B1(G900), .B2(new_n585), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n984), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G72));
  NAND3_X1  g817(.A1(new_n990), .A2(new_n997), .A3(new_n965), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n663), .A2(new_n410), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n976), .A2(new_n981), .A3(new_n982), .A4(new_n965), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n1006), .ZN(new_n1011));
  INV_X1    g825(.A(new_n700), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1006), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n426), .A2(KEYINPUT126), .ZN(new_n1015));
  INV_X1    g829(.A(new_n438), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(new_n426), .B2(KEYINPUT126), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1014), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n915), .B1(new_n907), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1009), .A2(new_n1013), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1009), .A2(new_n1013), .A3(KEYINPUT127), .A4(new_n1019), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1022), .A2(new_n1023), .ZN(G57));
endmodule


