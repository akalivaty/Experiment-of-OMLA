//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1207,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  AND2_X1   g0019(.A1(KEYINPUT67), .A2(G68), .ZN(new_n220));
  NOR2_X1   g0020(.A1(KEYINPUT67), .A2(G68), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G20), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT64), .ZN(new_n233));
  INV_X1    g0033(.A(G68), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n217), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g0035(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n236), .A2(G50), .A3(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT66), .Z(new_n239));
  AOI211_X1 g0039(.A(new_n209), .B(new_n229), .C1(new_n233), .C2(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n242), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G238), .B(G244), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G222), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G223), .A2(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n260), .B(new_n261), .C1(G77), .C2(new_n256), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n231), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n264), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n262), .B(new_n267), .C1(new_n212), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G200), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n230), .ZN(new_n276));
  OAI21_X1  g0076(.A(G20), .B1(new_n235), .B2(G50), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  INV_X1    g0078(.A(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n268), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n276), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n285), .A2(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(KEYINPUT68), .ZN(new_n287));
  INV_X1    g0087(.A(G13), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(new_n279), .A3(G1), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n286), .A2(new_n287), .B1(new_n211), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n276), .B1(new_n263), .B2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n273), .B1(new_n274), .B2(new_n272), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n294), .B2(new_n293), .ZN(new_n296));
  XOR2_X1   g0096(.A(new_n296), .B(KEYINPUT10), .Z(new_n297));
  INV_X1    g0097(.A(new_n293), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n272), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(G179), .B2(new_n272), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n282), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G20), .A2(G33), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n304), .A2(new_n305), .B1(G20), .B2(G77), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT15), .B(G87), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n283), .B2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n308), .A2(new_n276), .B1(new_n213), .B2(new_n289), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n291), .A2(G77), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G238), .A2(G1698), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n256), .B(new_n313), .C1(new_n218), .C2(G1698), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n261), .C1(G107), .C2(new_n256), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n267), .C1(new_n214), .C2(new_n271), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n299), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n312), .B(new_n317), .C1(G179), .C2(new_n316), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n297), .A2(new_n303), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n304), .A2(new_n289), .ZN(new_n320));
  INV_X1    g0120(.A(new_n291), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n304), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT69), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n268), .ZN(new_n325));
  NAND2_X1  g0125(.A1(KEYINPUT69), .A2(G33), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(KEYINPUT3), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G33), .ZN(new_n329));
  OR2_X1    g0129(.A1(G223), .A2(G1698), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n212), .A2(G1698), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n327), .A2(new_n329), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G87), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT75), .Z(new_n334));
  AOI21_X1  g0134(.A(new_n270), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n271), .A2(new_n218), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT77), .B(G190), .Z(new_n337));
  NOR4_X1   g0137(.A1(new_n335), .A2(new_n336), .A3(new_n266), .A4(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT78), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n335), .A2(new_n336), .A3(new_n266), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(G200), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n338), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(new_n343), .B2(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n329), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT7), .B1(new_n346), .B2(new_n279), .ZN(new_n347));
  AND2_X1   g0147(.A1(KEYINPUT69), .A2(G33), .ZN(new_n348));
  NOR2_X1   g0148(.A1(KEYINPUT69), .A2(G33), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n328), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(G20), .B1(new_n350), .B2(new_n345), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n347), .B1(new_n351), .B2(KEYINPUT7), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT73), .B1(new_n352), .B2(new_n223), .ZN(new_n353));
  OR2_X1    g0153(.A1(KEYINPUT67), .A2(G68), .ZN(new_n354));
  NAND2_X1  g0154(.A1(KEYINPUT67), .A2(G68), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G58), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n279), .B1(new_n356), .B2(new_n235), .ZN(new_n357));
  INV_X1    g0157(.A(G159), .ZN(new_n358));
  NOR4_X1   g0158(.A1(new_n358), .A2(KEYINPUT71), .A3(G20), .A4(G33), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT71), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n305), .B2(G159), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT3), .B1(new_n325), .B2(new_n326), .ZN(new_n364));
  INV_X1    g0164(.A(new_n345), .ZN(new_n365));
  OAI211_X1 g0165(.A(KEYINPUT7), .B(new_n279), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n256), .B2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(new_n370), .A3(new_n222), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n353), .A2(new_n363), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n276), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n327), .A2(new_n329), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n279), .ZN(new_n377));
  NAND2_X1  g0177(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n234), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n376), .A2(new_n279), .A3(new_n378), .A4(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT72), .B1(new_n357), .B2(new_n362), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT72), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT71), .B1(new_n280), .B2(new_n358), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n305), .A2(new_n360), .A3(G159), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G58), .A2(G68), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n222), .B2(G58), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n384), .B(new_n387), .C1(new_n389), .C2(new_n279), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n380), .A2(new_n382), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n375), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n374), .A2(new_n392), .A3(KEYINPUT74), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT74), .B1(new_n374), .B2(new_n392), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n323), .B(new_n344), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT74), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n370), .B1(new_n369), .B2(new_n222), .ZN(new_n399));
  AOI211_X1 g0199(.A(KEYINPUT73), .B(new_n223), .C1(new_n366), .C2(new_n368), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT16), .B1(new_n401), .B2(new_n363), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n380), .A2(new_n382), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n383), .A2(new_n390), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n276), .B1(new_n405), .B2(new_n373), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n398), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n374), .A2(new_n392), .A3(KEYINPUT74), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n323), .A4(new_n344), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n397), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n322), .B1(new_n407), .B2(new_n408), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n341), .A2(G179), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n299), .B2(new_n341), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT76), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT76), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n414), .B(new_n417), .C1(new_n299), .C2(new_n341), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n412), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n323), .B1(new_n393), .B2(new_n394), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT18), .A3(new_n419), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n411), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n222), .A2(new_n279), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n280), .A2(new_n211), .B1(new_n283), .B2(new_n213), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n276), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XOR2_X1   g0227(.A(new_n427), .B(KEYINPUT11), .Z(new_n428));
  INV_X1    g0228(.A(KEYINPUT12), .ZN(new_n429));
  OAI21_X1  g0229(.A(G68), .B1(new_n291), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n223), .A2(new_n289), .A3(KEYINPUT12), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n430), .B(new_n431), .C1(KEYINPUT12), .C2(new_n289), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G97), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n218), .A2(G1698), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G226), .B2(G1698), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n436), .B2(new_n346), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n266), .B1(new_n437), .B2(new_n261), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n219), .B2(new_n271), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT13), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n433), .B1(new_n440), .B2(new_n274), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(G200), .B2(new_n440), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(G169), .ZN(new_n443));
  XOR2_X1   g0243(.A(new_n443), .B(KEYINPUT14), .Z(new_n444));
  INV_X1    g0244(.A(G179), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n440), .ZN(new_n446));
  INV_X1    g0246(.A(new_n433), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n442), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n316), .A2(G200), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n311), .B(new_n449), .C1(new_n274), .C2(new_n316), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n424), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n319), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(new_n279), .C1(G33), .C2(new_n202), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n276), .C1(new_n279), .C2(G116), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n455), .B(KEYINPUT20), .ZN(new_n456));
  AOI211_X1 g0256(.A(new_n276), .B(new_n289), .C1(new_n263), .C2(G33), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(G116), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n289), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(G116), .B2(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n327), .A2(new_n329), .ZN(new_n461));
  OR2_X1    g0261(.A1(G257), .A2(G1698), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n461), .B(new_n462), .C1(G264), .C2(new_n257), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n346), .A2(G303), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n270), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n261), .B1(KEYINPUT5), .B2(new_n269), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n263), .A2(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT81), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT81), .B1(new_n467), .B2(new_n468), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n466), .A2(G274), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n261), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G270), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OR3_X1    g0278(.A1(new_n465), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n460), .A2(new_n479), .A3(G169), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT21), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR4_X1   g0282(.A1(new_n465), .A2(new_n474), .A3(new_n478), .A4(new_n445), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n460), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(new_n481), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n465), .A2(new_n474), .A3(new_n478), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n337), .ZN(new_n488));
  INV_X1    g0288(.A(G200), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n487), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n486), .B1(new_n460), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n461), .B1(G257), .B2(new_n257), .ZN(new_n492));
  NOR2_X1   g0292(.A1(G250), .A2(G1698), .ZN(new_n493));
  INV_X1    g0293(.A(G294), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n348), .A2(new_n349), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n492), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n261), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n476), .A2(G264), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(G190), .A3(new_n473), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT24), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n327), .A2(new_n279), .A3(G87), .A4(new_n329), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT22), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n504), .A2(KEYINPUT87), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(KEYINPUT87), .ZN(new_n506));
  NOR4_X1   g0306(.A1(new_n346), .A2(KEYINPUT22), .A3(G20), .A4(new_n225), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G116), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n495), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n279), .B2(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n510), .A2(new_n279), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n502), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n504), .B(KEYINPUT87), .ZN(new_n517));
  OAI211_X1 g0317(.A(KEYINPUT24), .B(new_n514), .C1(new_n517), .C2(new_n507), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n276), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n457), .A2(G107), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n289), .A2(new_n203), .ZN(new_n521));
  XOR2_X1   g0321(.A(new_n521), .B(KEYINPUT25), .Z(new_n522));
  NAND4_X1  g0322(.A1(new_n501), .A2(new_n519), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n499), .A2(new_n474), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(new_n489), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n499), .A2(G179), .A3(new_n474), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n500), .A2(new_n473), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n299), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n491), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G238), .A2(G1698), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n214), .B2(G1698), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n461), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n510), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n261), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT82), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n468), .A2(new_n226), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n263), .A2(new_n265), .A3(G45), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n270), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n539), .A2(new_n540), .A3(new_n445), .A4(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n510), .B1(new_n461), .B2(new_n535), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n445), .B(new_n543), .C1(new_n545), .C2(new_n270), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT82), .ZN(new_n547));
  INV_X1    g0347(.A(new_n543), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n538), .B2(new_n261), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n544), .B(new_n547), .C1(G169), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT83), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n461), .A2(new_n279), .A3(G68), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT19), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n283), .B2(new_n202), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n279), .B1(new_n434), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G87), .B2(new_n204), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n276), .B1(new_n289), .B2(new_n307), .ZN(new_n558));
  INV_X1    g0358(.A(new_n457), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n307), .B(KEYINPUT84), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n539), .A2(new_n543), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n299), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT83), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n544), .A4(new_n547), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n551), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n557), .A2(new_n276), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n307), .A2(new_n289), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n457), .A2(G87), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT85), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n562), .B2(new_n274), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n549), .A2(KEYINPUT85), .A3(G190), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n549), .A2(new_n489), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n566), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT86), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT86), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n566), .A2(new_n580), .A3(new_n577), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT4), .B1(new_n346), .B2(new_n226), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n376), .A2(new_n214), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n584), .B(new_n585), .C1(KEYINPUT4), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n261), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n476), .A2(G257), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n473), .A3(new_n589), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n590), .A2(new_n274), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n559), .A2(new_n202), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n459), .A2(G97), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n369), .A2(G107), .B1(G77), .B2(new_n305), .ZN(new_n595));
  XNOR2_X1  g0395(.A(G97), .B(G107), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT79), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(KEYINPUT6), .ZN(new_n598));
  MUX2_X1   g0398(.A(new_n597), .B(new_n203), .S(KEYINPUT6), .Z(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT80), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n595), .B1(new_n602), .B2(new_n279), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n594), .B1(new_n603), .B2(new_n276), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n590), .A2(G200), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n591), .A2(new_n593), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n276), .ZN(new_n607));
  INV_X1    g0407(.A(new_n594), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n593), .A3(new_n608), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n590), .A2(G179), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n590), .A2(new_n299), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n582), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n452), .A2(new_n533), .A3(new_n614), .ZN(G372));
  INV_X1    g0415(.A(new_n612), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n579), .A2(KEYINPUT26), .A3(new_n581), .A4(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n572), .A2(new_n573), .B1(new_n575), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n570), .A2(KEYINPUT89), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT89), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n558), .A2(new_n622), .A3(new_n569), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n576), .A2(KEYINPUT88), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n620), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n561), .A2(new_n563), .A3(new_n546), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n618), .B1(new_n628), .B2(new_n612), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n617), .A2(KEYINPUT91), .A3(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n566), .A2(new_n580), .A3(new_n577), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n580), .B1(new_n566), .B2(new_n577), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT91), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT26), .A4(new_n616), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT90), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n531), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT90), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n486), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n523), .A2(new_n525), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n640), .A2(new_n613), .A3(new_n628), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n630), .A2(new_n635), .A3(new_n627), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n452), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n397), .A2(new_n410), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n446), .A2(new_n447), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n442), .A2(new_n318), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n422), .A2(new_n415), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(new_n412), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n302), .B1(new_n652), .B2(new_n297), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n644), .A2(new_n653), .ZN(G369));
  NAND3_X1  g0454(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n288), .A2(G20), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n263), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n460), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n491), .B2(new_n663), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n530), .A2(new_n662), .ZN(new_n669));
  INV_X1    g0469(.A(new_n662), .ZN(new_n670));
  OAI22_X1  g0470(.A1(new_n532), .A2(new_n669), .B1(new_n531), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n486), .A2(new_n662), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n531), .A3(new_n526), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n637), .A2(new_n638), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n670), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n207), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n238), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT26), .B1(new_n628), .B2(new_n612), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n627), .B(KEYINPUT95), .ZN(new_n688));
  INV_X1    g0488(.A(new_n613), .ZN(new_n689));
  INV_X1    g0489(.A(new_n628), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n526), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n655), .B1(new_n530), .B2(new_n529), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n687), .B(new_n688), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n582), .A2(KEYINPUT26), .A3(new_n612), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n670), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n643), .A2(new_n697), .A3(new_n670), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n524), .A2(new_n549), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n445), .A3(new_n479), .A4(new_n590), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n483), .A2(KEYINPUT92), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n590), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(KEYINPUT93), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n499), .B1(new_n483), .B2(KEYINPUT92), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n704), .A2(new_n549), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(KEYINPUT93), .ZN(new_n709));
  AND4_X1   g0509(.A1(new_n549), .A2(new_n704), .A3(new_n709), .A4(new_n707), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n702), .B(new_n708), .C1(new_n710), .C2(new_n706), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT31), .B1(new_n711), .B2(new_n662), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT94), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n662), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n712), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n533), .A2(new_n614), .A3(new_n670), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n715), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n700), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n686), .B1(new_n725), .B2(G1), .ZN(G364));
  INV_X1    g0526(.A(new_n668), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n656), .A2(G45), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n682), .A2(G1), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n666), .A2(new_n667), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n666), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n461), .A2(new_n680), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G45), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n737), .B1(new_n239), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n738), .B2(new_n251), .ZN(new_n740));
  INV_X1    g0540(.A(G355), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n256), .A2(new_n207), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n740), .B1(G116), .B2(new_n207), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n230), .B1(G20), .B2(new_n299), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n729), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n279), .A2(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(G190), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G87), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n279), .A2(new_n445), .A3(new_n489), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT98), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT98), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(new_n337), .A3(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n279), .A2(new_n445), .A3(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n274), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n751), .B1(new_n755), .B2(new_n211), .C1(new_n760), .C2(new_n213), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT32), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n748), .A2(new_n274), .A3(new_n489), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT99), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT99), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n762), .B1(new_n766), .B2(new_n358), .ZN(new_n767));
  INV_X1    g0567(.A(new_n766), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(KEYINPUT32), .A3(G159), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n761), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n274), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n279), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G97), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n748), .A2(new_n274), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n203), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n337), .A2(new_n756), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT96), .Z(new_n778));
  AOI21_X1  g0578(.A(new_n776), .B1(new_n778), .B2(G58), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n753), .A2(new_n274), .A3(new_n754), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT100), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n346), .B1(new_n781), .B2(G68), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n770), .A2(new_n774), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n786), .B2(new_n775), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G303), .B2(new_n750), .ZN(new_n788));
  INV_X1    g0588(.A(new_n757), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G311), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n256), .B1(new_n768), .B2(G329), .ZN(new_n791));
  INV_X1    g0591(.A(G326), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n755), .A2(new_n792), .B1(new_n494), .B2(new_n772), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT101), .Z(new_n794));
  NAND4_X1  g0594(.A1(new_n788), .A2(new_n790), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n777), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n796), .A2(G322), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n783), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n744), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n735), .A2(new_n746), .A3(new_n747), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n731), .A2(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n643), .A2(new_n670), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n318), .A2(new_n662), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n450), .B1(new_n311), .B2(new_n670), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n318), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n802), .B(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(new_n723), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n729), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n781), .B(KEYINPUT102), .ZN(new_n812));
  INV_X1    g0612(.A(new_n760), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n812), .A2(G283), .B1(G116), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n755), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G303), .B1(G294), .B2(new_n796), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n774), .C1(new_n817), .C2(new_n766), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G107), .B2(new_n750), .ZN(new_n819));
  INV_X1    g0619(.A(new_n775), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G87), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n814), .A2(new_n819), .A3(new_n346), .A4(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n781), .A2(G150), .B1(G159), .B2(new_n813), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  INV_X1    g0624(.A(G143), .ZN(new_n825));
  INV_X1    g0625(.A(new_n778), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n823), .B1(new_n824), .B2(new_n755), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT34), .Z(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G50), .B2(new_n750), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n775), .A2(new_n234), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n768), .A2(G132), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n773), .A2(G58), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n829), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n822), .B1(new_n834), .B2(new_n376), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(new_n744), .B1(new_n732), .B2(new_n807), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n744), .A2(new_n732), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n213), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n747), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT103), .Z(new_n840));
  NAND2_X1  g0640(.A1(new_n811), .A2(new_n840), .ZN(G384));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT37), .B1(new_n422), .B2(new_n419), .ZN(new_n843));
  INV_X1    g0643(.A(new_n660), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n422), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n395), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n415), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n395), .B1(new_n413), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT107), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n650), .A2(KEYINPUT107), .A3(new_n395), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n845), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n847), .B1(new_n853), .B2(KEYINPUT37), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n845), .B1(new_n651), .B2(new_n645), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n842), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n391), .A2(KEYINPUT16), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n323), .B1(new_n406), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n415), .B2(new_n844), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n857), .B1(new_n395), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n846), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n859), .A2(new_n844), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT38), .B(new_n863), .C1(new_n424), .C2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT108), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n413), .A2(new_n412), .A3(new_n420), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT18), .B1(new_n422), .B2(new_n419), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n397), .B(new_n410), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n864), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n871), .A2(new_n872), .B1(new_n846), .B2(new_n862), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(KEYINPUT108), .A3(KEYINPUT38), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n856), .A2(new_n867), .A3(new_n868), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT109), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT108), .B1(new_n873), .B2(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n421), .A2(new_n423), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n864), .B1(new_n645), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n395), .B1(new_n413), .B2(new_n660), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n861), .B1(new_n881), .B2(new_n843), .ZN(new_n882));
  NOR4_X1   g0682(.A1(new_n879), .A2(new_n882), .A3(new_n866), .A4(new_n842), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT109), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n884), .A2(new_n885), .A3(new_n868), .A4(new_n856), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n842), .B1(new_n879), .B2(new_n882), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n865), .A3(KEYINPUT105), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT105), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n889), .B(new_n842), .C1(new_n879), .C2(new_n882), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT106), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n888), .A2(KEYINPUT106), .A3(KEYINPUT39), .A4(new_n890), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n876), .A2(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n646), .A2(new_n662), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n651), .A2(new_n844), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n643), .A2(new_n670), .A3(new_n808), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n804), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n447), .A2(new_n662), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n647), .A2(new_n662), .B1(new_n448), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n888), .A2(new_n890), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n898), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n699), .A2(new_n452), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n653), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n721), .A2(new_n718), .A3(new_n712), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n808), .A3(new_n904), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n856), .B2(new_n884), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(KEYINPUT110), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(KEYINPUT110), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n913), .A2(new_n808), .A3(new_n904), .A4(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n918), .A2(new_n920), .A3(new_n907), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n452), .A2(new_n913), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(new_n667), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n912), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n263), .B2(new_n656), .ZN(new_n927));
  INV_X1    g0727(.A(new_n602), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n509), .B1(new_n928), .B2(KEYINPUT35), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n233), .C1(KEYINPUT35), .C2(new_n928), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT36), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n234), .A2(G50), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT104), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n356), .A2(G77), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n933), .B1(new_n238), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(G1), .A3(new_n288), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n927), .A2(new_n931), .A3(new_n936), .ZN(G367));
  NOR2_X1   g0737(.A1(new_n675), .A2(new_n613), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n609), .A2(new_n662), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n689), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n612), .B1(new_n941), .B2(new_n531), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n670), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n621), .A2(new_n623), .A3(new_n662), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n690), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n627), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n939), .A2(new_n943), .B1(KEYINPUT43), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n941), .B1(new_n612), .B2(new_n670), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n674), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n950), .B(new_n953), .Z(new_n954));
  XNOR2_X1  g0754(.A(new_n681), .B(KEYINPUT41), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT112), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n668), .A2(new_n673), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n676), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n725), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT112), .B1(new_n724), .B2(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n675), .A2(new_n678), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n952), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n952), .ZN(new_n966));
  XOR2_X1   g0766(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n965), .A2(new_n674), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n674), .B1(new_n965), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n961), .A2(new_n962), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT113), .Z(new_n973));
  AOI21_X1  g0773(.A(new_n956), .B1(new_n973), .B2(new_n725), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n728), .A2(G1), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n954), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n775), .A2(new_n202), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G107), .B2(new_n773), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n755), .B2(new_n817), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n813), .A2(G283), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT46), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n749), .B2(new_n509), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n750), .A2(KEYINPUT46), .A3(G116), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n980), .A2(new_n376), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n979), .B(new_n984), .C1(G317), .C2(new_n768), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n812), .A2(G294), .ZN(new_n986));
  INV_X1    g0786(.A(G303), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n985), .B(new_n986), .C1(new_n987), .C2(new_n826), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT114), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n820), .A2(G77), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n256), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n812), .A2(G159), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n813), .A2(G50), .B1(KEYINPUT114), .B2(new_n991), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n773), .A2(G68), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n825), .C2(new_n755), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G58), .B2(new_n750), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n993), .B(new_n997), .C1(new_n824), .C2(new_n766), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n777), .A2(new_n278), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n988), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n744), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n945), .A2(new_n734), .A3(new_n946), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n745), .B1(new_n207), .B2(new_n307), .C1(new_n243), .C2(new_n737), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1003), .A2(new_n747), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n976), .A2(new_n1006), .ZN(G387));
  OR3_X1    g0807(.A1(new_n282), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT50), .B1(new_n282), .B2(G50), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1008), .A2(new_n1009), .A3(new_n738), .A4(new_n683), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n234), .A2(new_n213), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n736), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT116), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n738), .B2(new_n247), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(G107), .B2(new_n207), .C1(new_n683), .C2(new_n742), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n729), .B1(new_n1015), .B2(new_n745), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT117), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n560), .A2(new_n772), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n211), .B2(new_n777), .C1(new_n278), .C2(new_n766), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n977), .B(new_n1019), .C1(G159), .C2(new_n815), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n750), .A2(G77), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n789), .A2(G68), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n376), .B1(new_n781), .B2(new_n304), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n812), .A2(G311), .B1(G322), .B2(new_n815), .ZN(new_n1025));
  INV_X1    g0825(.A(G317), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1025), .B1(new_n987), .B2(new_n760), .C1(new_n1026), .C2(new_n826), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n786), .B2(new_n772), .C1(new_n494), .C2(new_n749), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT49), .Z(new_n1030));
  OAI221_X1 g0830(.A(new_n376), .B1(new_n509), .B2(new_n775), .C1(new_n766), .C2(new_n792), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1024), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT118), .Z(new_n1033));
  AOI21_X1  g0833(.A(new_n1017), .B1(new_n1033), .B2(new_n744), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n671), .A2(G20), .A3(new_n733), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1034), .A2(new_n1035), .B1(new_n975), .B2(new_n960), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n961), .A2(new_n962), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n725), .B2(new_n960), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1036), .B1(new_n1038), .B2(new_n682), .ZN(G393));
  OAI21_X1  g0839(.A(new_n1037), .B1(new_n969), .B2(new_n970), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n973), .A2(new_n681), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n952), .A2(new_n734), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n755), .A2(new_n278), .B1(new_n358), .B2(new_n777), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT51), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n222), .B2(new_n750), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n813), .A2(new_n304), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n812), .A2(G50), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n821), .B1(new_n213), .B2(new_n772), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n376), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G143), .B2(new_n768), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n812), .A2(G303), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n755), .A2(new_n1026), .B1(new_n817), .B2(new_n777), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n773), .A2(G116), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n768), .A2(G322), .B1(G294), .B2(new_n789), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n749), .A2(new_n786), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n1057), .A2(new_n256), .A3(new_n776), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n744), .B1(new_n1051), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n745), .B1(new_n202), .B2(new_n207), .C1(new_n737), .C2(new_n254), .ZN(new_n1061));
  AND4_X1   g0861(.A1(new_n747), .A2(new_n1042), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n971), .B2(new_n975), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1041), .A2(new_n1063), .ZN(G390));
  NAND2_X1  g0864(.A1(new_n886), .A2(new_n876), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n893), .A2(new_n894), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n905), .A2(new_n897), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n670), .B(new_n806), .C1(new_n693), .C2(new_n694), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n804), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n896), .B1(new_n1070), .B2(new_n904), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n884), .A2(new_n856), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n722), .A2(G330), .A3(new_n808), .A4(new_n904), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1068), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n913), .A2(G330), .A3(new_n808), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1077), .A2(new_n903), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n722), .A2(G330), .A3(new_n808), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n903), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n1078), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n901), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1077), .A2(new_n903), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1070), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1074), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n452), .A2(new_n913), .A3(G330), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n910), .A2(new_n653), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n682), .B1(new_n1081), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1091), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1095));
  OAI211_X1 g0895(.A(KEYINPUT119), .B(new_n1095), .C1(new_n1076), .C2(new_n1080), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1068), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1073), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n895), .B2(new_n1067), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1100), .B2(new_n1079), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT119), .B1(new_n1101), .B2(new_n1095), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1094), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n975), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n895), .A2(new_n732), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n812), .A2(G107), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n777), .A2(new_n509), .B1(new_n213), .B2(new_n772), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT121), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n830), .B(new_n1108), .C1(G283), .C2(new_n815), .ZN(new_n1109));
  AND4_X1   g0909(.A1(new_n346), .A2(new_n1106), .A3(new_n1109), .A4(new_n751), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n202), .B2(new_n760), .C1(new_n494), .C2(new_n766), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT122), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n812), .A2(G137), .B1(G50), .B2(new_n820), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n815), .A2(G128), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n749), .A2(new_n278), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n256), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n772), .A2(new_n358), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT54), .B(G143), .Z(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n760), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n796), .A2(G132), .ZN(new_n1122));
  INV_X1    g0922(.A(G125), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n766), .B2(new_n1123), .ZN(new_n1124));
  NOR4_X1   g0924(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n744), .B1(new_n1112), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n729), .B1(new_n282), .B2(new_n837), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT120), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1105), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1103), .A2(new_n1104), .A3(new_n1129), .ZN(G378));
  INV_X1    g0930(.A(KEYINPUT57), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1095), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT119), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1091), .B1(new_n1134), .B2(new_n1096), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n297), .A2(new_n303), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1137));
  XOR2_X1   g0937(.A(new_n1136), .B(new_n1137), .Z(new_n1138));
  NAND2_X1  g0938(.A1(new_n293), .A2(new_n844), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1138), .B(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n922), .B2(new_n667), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1140), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1142), .B(G330), .C1(new_n917), .C2(new_n921), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n909), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n898), .A4(new_n908), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1131), .B1(new_n1135), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1092), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(KEYINPUT57), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n1151), .A3(new_n681), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1142), .A2(new_n732), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n757), .A2(new_n824), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1120), .A2(new_n749), .B1(new_n772), .B2(new_n278), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n781), .C2(G132), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1156), .B1(new_n1123), .B2(new_n755), .C1(new_n1157), .C2(new_n777), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n820), .A2(G159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G41), .B1(new_n768), .B2(G124), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1159), .A2(new_n268), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1163));
  AOI21_X1  g0963(.A(G41), .B1(new_n348), .B2(KEYINPUT3), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n1162), .A2(new_n1163), .B1(G50), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n820), .A2(G58), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n995), .B(new_n1166), .C1(new_n766), .C2(new_n786), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1021), .B1(new_n203), .B2(new_n777), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n269), .B(new_n376), .C1(new_n560), .C2(new_n757), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n509), .B2(new_n755), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G97), .B2(new_n781), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT58), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n744), .B1(new_n1165), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n837), .A2(new_n211), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1153), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n747), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n975), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1177), .B1(new_n1147), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1152), .A2(new_n1180), .ZN(G375));
  NAND2_X1  g0981(.A1(new_n768), .A2(G303), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n256), .B1(new_n796), .B2(G283), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n750), .A2(G97), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1182), .A2(new_n990), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n812), .A2(G116), .B1(G294), .B2(new_n815), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1186), .B(new_n1018), .C1(new_n203), .C2(new_n760), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n757), .A2(new_n278), .B1(new_n772), .B2(new_n211), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1166), .B1(new_n826), .B2(new_n824), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(G132), .C2(new_n815), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n376), .B1(new_n812), .B2(new_n1119), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n358), .C2(new_n749), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n766), .A2(new_n1157), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1185), .A2(new_n1187), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n744), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n747), .B(new_n1195), .C1(new_n904), .C2(new_n733), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n234), .B2(new_n837), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1089), .B2(new_n975), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n955), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n1095), .ZN(G381));
  INV_X1    g1000(.A(G390), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n976), .A3(new_n1006), .ZN(new_n1202));
  OR2_X1    g1002(.A1(G381), .A2(G384), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1202), .A2(G396), .A3(G393), .A4(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(G375), .A2(G378), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(G407));
  OAI21_X1  g1006(.A(new_n1205), .B1(new_n1204), .B2(new_n661), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(G213), .ZN(G409));
  NAND2_X1  g1008(.A1(G375), .A2(G378), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT60), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1085), .A2(KEYINPUT60), .A3(new_n1091), .A4(new_n1088), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1211), .A2(new_n681), .A3(new_n1093), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1198), .ZN(new_n1214));
  INV_X1    g1014(.A(G384), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(G384), .A3(new_n1198), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(G213), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(G343), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1135), .A2(new_n956), .A3(new_n1147), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1223), .A2(G378), .A3(new_n1179), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1209), .A2(new_n1219), .A3(new_n1222), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1221), .A2(G2897), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1219), .B2(KEYINPUT123), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1218), .A2(new_n1229), .A3(G2897), .A4(new_n1221), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1219), .A2(KEYINPUT123), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1221), .B1(G375), .B2(G378), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1232), .B1(new_n1233), .B2(new_n1225), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT63), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1226), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT61), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT124), .B1(new_n1226), .B2(new_n1235), .ZN(new_n1238));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1152), .B2(new_n1180), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1240), .A2(new_n1218), .A3(new_n1224), .A4(new_n1221), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT124), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(KEYINPUT63), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G393), .B(G396), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1202), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1201), .B1(new_n976), .B2(new_n1006), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G387), .A2(G390), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1202), .A3(new_n1245), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT126), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1241), .B2(KEYINPUT62), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1233), .A2(KEYINPUT62), .A3(new_n1219), .A4(new_n1225), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT127), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1240), .A2(new_n1221), .A3(new_n1224), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(KEYINPUT62), .A4(new_n1219), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1226), .A2(KEYINPUT126), .A3(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1254), .A2(new_n1256), .A3(new_n1259), .A4(new_n1261), .ZN(new_n1262));
  XOR2_X1   g1062(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1263));
  NOR3_X1   g1063(.A1(new_n1252), .A2(new_n1234), .A3(new_n1263), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1244), .A2(new_n1252), .B1(new_n1262), .B2(new_n1264), .ZN(G405));
  NAND2_X1  g1065(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1205), .A2(new_n1240), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1249), .B(new_n1251), .C1(new_n1205), .C2(new_n1240), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(new_n1219), .ZN(G402));
endmodule


