//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT64), .Z(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G137), .A4(new_n463), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(G2105), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT65), .B1(new_n473), .B2(G101), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n463), .A2(KEYINPUT65), .A3(G101), .A4(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT66), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n475), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(new_n483), .A3(new_n472), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n467), .B1(new_n478), .B2(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n469), .A2(new_n471), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n486), .A2(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NOR3_X1   g067(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n493));
  OAI221_X1 g068(.A(G2104), .B1(G112), .B2(new_n463), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n488), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  NAND4_X1  g071(.A1(new_n469), .A2(new_n471), .A3(G138), .A4(new_n463), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT68), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n464), .A2(G138), .A3(new_n463), .A4(new_n499), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n464), .A2(G126), .A3(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT69), .A2(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(KEYINPUT69), .A2(KEYINPUT6), .A3(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n518), .A2(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n514), .A2(new_n521), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n524), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n522), .A2(new_n523), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT70), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n511), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n528), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  INV_X1    g112(.A(new_n520), .ZN(new_n538));
  INV_X1    g113(.A(G51), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n535), .A2(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n533), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n524), .A2(G90), .B1(new_n520), .B2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND3_X1  g123(.A1(new_n530), .A2(new_n532), .A3(G56), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT71), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n553), .A3(new_n550), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(G651), .A3(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n524), .A2(G81), .B1(new_n520), .B2(G43), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(KEYINPUT72), .ZN(new_n565));
  INV_X1    g140(.A(new_n519), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT6), .B1(KEYINPUT69), .B2(G651), .ZN(new_n567));
  OAI211_X1 g142(.A(G543), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n520), .A2(new_n570), .A3(new_n565), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n511), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n569), .A2(new_n571), .B1(G651), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n566), .A2(new_n567), .B1(new_n510), .B2(new_n509), .ZN(new_n577));
  INV_X1    g152(.A(G91), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n524), .A2(KEYINPUT73), .A3(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n575), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G168), .ZN(G286));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  NOR3_X1   g159(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT70), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n531), .B1(new_n522), .B2(new_n523), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n524), .A2(G87), .B1(new_n520), .B2(G49), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G288));
  INV_X1    g165(.A(G651), .ZN(new_n591));
  OAI21_X1  g166(.A(G61), .B1(new_n509), .B2(new_n510), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n524), .A2(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n520), .A2(G48), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND3_X1  g173(.A1(new_n530), .A2(new_n532), .A3(G60), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n591), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n524), .A2(G85), .B1(new_n520), .B2(G47), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n524), .A2(G92), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT10), .Z(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT74), .B(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n511), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n606), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n606), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(G286), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(G299), .B(KEYINPUT75), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G297));
  XOR2_X1   g195(.A(G297), .B(KEYINPUT76), .Z(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n614), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n614), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n487), .A2(G2104), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n487), .A2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n489), .A2(G123), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT79), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT80), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n653), .B2(new_n654), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n660), .B2(KEYINPUT81), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(KEYINPUT81), .B2(new_n660), .ZN(new_n665));
  INV_X1    g240(.A(new_n659), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n660), .B(KEYINPUT17), .Z(new_n667));
  INV_X1    g242(.A(new_n661), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n665), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n668), .A3(new_n659), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n663), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT82), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT83), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT85), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT84), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G35), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G162), .B2(new_n695), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT29), .Z(new_n698));
  INV_X1    g273(.A(G2090), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G20), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT23), .ZN(new_n702));
  INV_X1    g277(.A(G299), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n700), .ZN(new_n704));
  INV_X1    g279(.A(G1956), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  OAI22_X1  g282(.A1(new_n698), .A2(new_n699), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT98), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n614), .A2(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G4), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1348), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n698), .A2(new_n699), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT97), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(new_n713), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n487), .A2(G140), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n489), .A2(G128), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g296(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n722));
  OAI221_X1 g297(.A(G2104), .B1(G116), .B2(new_n463), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n718), .A2(new_n719), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n695), .A2(G26), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G2067), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  AND4_X1   g305(.A1(new_n714), .A2(new_n716), .A3(new_n717), .A4(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n708), .A2(new_n709), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n700), .A2(G19), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n557), .B2(new_n700), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1341), .Z(new_n735));
  AND4_X1   g310(.A1(new_n710), .A2(new_n731), .A3(new_n732), .A4(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n695), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n487), .A2(G139), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT91), .Z(new_n742));
  AOI22_X1  g317(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n463), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(G29), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(new_n442), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT92), .ZN(new_n747));
  NOR2_X1   g322(.A1(G27), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT95), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(new_n443), .ZN(new_n751));
  NAND2_X1  g326(.A1(G160), .A2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n753), .B2(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT24), .B2(new_n753), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(G2084), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n700), .A2(G5), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G171), .B2(new_n700), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n745), .A2(new_n442), .B1(G1961), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n747), .A2(new_n751), .A3(new_n756), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G29), .A2(G32), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n489), .A2(G129), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT93), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n473), .A2(G105), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT26), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n764), .B(new_n766), .C1(G141), .C2(new_n487), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n763), .A2(KEYINPUT94), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(KEYINPUT94), .B1(new_n763), .B2(new_n767), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n761), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(G2084), .B1(new_n752), .B2(new_n755), .ZN(new_n775));
  INV_X1    g350(.A(new_n758), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G168), .A2(new_n700), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n700), .B2(G21), .ZN(new_n780));
  INV_X1    g355(.A(G1966), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT30), .B(G28), .ZN(new_n783));
  OR2_X1    g358(.A1(KEYINPUT31), .A2(G11), .ZN(new_n784));
  NAND2_X1  g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n783), .A2(new_n695), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n638), .B2(new_n695), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n780), .B2(new_n781), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n778), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n774), .A2(new_n789), .ZN(new_n790));
  OR3_X1    g365(.A1(new_n760), .A2(KEYINPUT96), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(KEYINPUT96), .B1(new_n760), .B2(new_n790), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n736), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT99), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT99), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n736), .A2(new_n791), .A3(new_n795), .A4(new_n792), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n700), .A2(G23), .ZN(new_n797));
  INV_X1    g372(.A(G288), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n700), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT33), .B(G1976), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G22), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G166), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT88), .B(G1971), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n801), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n700), .A2(G24), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n604), .B2(new_n700), .ZN(new_n813));
  INV_X1    g388(.A(G1986), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n695), .A2(G25), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n487), .A2(G131), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n489), .A2(G119), .ZN(new_n818));
  OR2_X1    g393(.A1(G95), .A2(G2105), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n819), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT86), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT86), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n816), .B1(new_n825), .B2(new_n695), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT35), .B(G1991), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT87), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n810), .A2(new_n811), .A3(new_n815), .A4(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT89), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT36), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n831), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n794), .A2(new_n796), .B1(new_n833), .B2(new_n835), .ZN(G311));
  NAND2_X1  g411(.A1(new_n794), .A2(new_n796), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(G150));
  NAND2_X1  g414(.A1(new_n614), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n530), .A2(new_n532), .A3(G67), .ZN(new_n842));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n591), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n520), .A2(G55), .ZN(new_n845));
  INV_X1    g420(.A(G93), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n577), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n557), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n555), .A2(new_n556), .ZN(new_n850));
  INV_X1    g425(.A(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n841), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n855));
  AOI21_X1  g430(.A(G860), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT100), .Z(G145));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n862));
  XNOR2_X1  g437(.A(G160), .B(G162), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n638), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n489), .A2(G130), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n463), .A2(G118), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G142), .B2(new_n487), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n824), .B(new_n869), .Z(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(new_n630), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n724), .B(new_n506), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n769), .B2(new_n770), .ZN(new_n874));
  INV_X1    g449(.A(new_n770), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(KEYINPUT101), .A3(new_n768), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n744), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n763), .A2(new_n767), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n744), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n872), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n872), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n874), .A2(new_n876), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n882), .B(new_n879), .C1(new_n883), .C2(new_n744), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n871), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n881), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n870), .B(new_n630), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n864), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n864), .B1(new_n886), .B2(new_n888), .ZN(new_n894));
  AOI21_X1  g469(.A(G37), .B1(new_n894), .B2(new_n885), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n893), .B1(new_n892), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n862), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n892), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT103), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n898), .A2(new_n902), .ZN(G395));
  XNOR2_X1  g478(.A(new_n853), .B(new_n624), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n613), .A2(new_n703), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT104), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n613), .A2(new_n907), .A3(new_n703), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n614), .A2(G299), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(KEYINPUT41), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n906), .A2(new_n909), .A3(new_n913), .A4(new_n908), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n911), .B1(new_n904), .B2(new_n915), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n917));
  XOR2_X1   g492(.A(G303), .B(KEYINPUT105), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G305), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n604), .B(G288), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n917), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g501(.A(new_n925), .B1(G868), .B2(new_n848), .ZN(G331));
  AND2_X1   g502(.A1(new_n849), .A2(new_n852), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n545), .A2(new_n929), .A3(new_n546), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n545), .B2(new_n546), .ZN(new_n932));
  OAI21_X1  g507(.A(G286), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n932), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(G168), .A3(new_n930), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n853), .A2(new_n935), .A3(new_n933), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n928), .A2(KEYINPUT107), .A3(new_n936), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n940), .A2(new_n912), .A3(new_n914), .A4(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n937), .A2(new_n910), .A3(new_n938), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n921), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G37), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  INV_X1    g523(.A(new_n921), .ZN(new_n949));
  INV_X1    g524(.A(new_n910), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n940), .B2(new_n941), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n915), .B1(new_n937), .B2(new_n938), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n946), .A2(new_n947), .A3(new_n948), .A4(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n953), .A2(new_n944), .A3(new_n948), .A4(new_n945), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT108), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n944), .A2(new_n945), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n921), .B1(new_n942), .B2(new_n943), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n953), .A2(new_n945), .A3(new_n944), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n963), .B2(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(new_n958), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n946), .A2(new_n948), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT109), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n964), .A2(new_n966), .A3(KEYINPUT109), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n962), .B1(new_n967), .B2(new_n968), .ZN(G397));
  INV_X1    g544(.A(KEYINPUT127), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n506), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n465), .A2(new_n466), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G2105), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n482), .A2(new_n483), .A3(new_n472), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n483), .B1(new_n482), .B2(new_n472), .ZN(new_n978));
  OAI211_X1 g553(.A(G40), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n724), .B(G2067), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(G1996), .B2(new_n878), .ZN(new_n982));
  INV_X1    g557(.A(new_n771), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(G1996), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n824), .B(new_n828), .Z(new_n985));
  OAI21_X1  g560(.A(new_n980), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(G290), .A2(G1986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n604), .A2(new_n814), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n980), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT110), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT122), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  INV_X1    g568(.A(G2084), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n506), .A2(new_n995), .A3(new_n971), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n506), .B2(new_n971), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n996), .A2(new_n979), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G40), .ZN(new_n999));
  AOI211_X1 g574(.A(new_n999), .B(new_n467), .C1(new_n478), .C2(new_n484), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n974), .A3(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n994), .A2(new_n998), .B1(new_n1002), .B2(new_n781), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n993), .B1(new_n1003), .B2(G168), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n992), .B1(new_n1004), .B2(KEYINPUT51), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(KEYINPUT121), .A3(KEYINPUT51), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n506), .B2(new_n971), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(new_n979), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n972), .A2(KEYINPUT50), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n506), .A2(new_n995), .A3(new_n971), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1000), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  OAI22_X1  g587(.A1(G1966), .A2(new_n1009), .B1(new_n1012), .B2(G2084), .ZN(new_n1013));
  OAI21_X1  g588(.A(G8), .B1(new_n1013), .B2(G286), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(KEYINPUT122), .A3(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT51), .B(G8), .C1(new_n1013), .C2(G286), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1005), .A2(new_n1006), .A3(new_n1016), .A4(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1013), .A2(G8), .A3(G286), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1976), .B1(new_n588), .B2(new_n589), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1023), .B(G8), .C1(new_n979), .C2(new_n972), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G8), .B1(new_n979), .B2(new_n972), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1024), .B(new_n1025), .C1(new_n1027), .C2(new_n1030), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(G1981), .B1(new_n594), .B2(KEYINPUT113), .ZN(new_n1035));
  XNOR2_X1  g610(.A(G305), .B(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1027), .B1(new_n1036), .B2(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  OAI211_X1 g613(.A(G305), .B(G1981), .C1(KEYINPUT113), .C2(new_n594), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1035), .A2(new_n596), .A3(new_n597), .A4(new_n595), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT114), .B(KEYINPUT49), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1037), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G303), .A2(G8), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n1046), .B(KEYINPUT55), .Z(new_n1047));
  INV_X1    g622(.A(G1971), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1002), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1000), .A2(new_n699), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n993), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1034), .B(new_n1045), .C1(new_n1047), .C2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1009), .B2(G1971), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(G8), .A3(new_n1047), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT111), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1056), .A3(new_n1047), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1052), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1007), .A2(new_n1008), .A3(G2078), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n979), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(G160), .A2(KEYINPUT123), .A3(G40), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1059), .A2(KEYINPUT53), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1000), .A2(new_n443), .A3(new_n974), .A4(new_n1001), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1012), .A2(new_n777), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1063), .A2(new_n1066), .A3(G301), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT124), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1065), .A2(new_n1064), .B1(new_n1012), .B2(new_n777), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(G301), .A4(new_n1063), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1059), .A2(KEYINPUT53), .A3(new_n1000), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1066), .A2(new_n1073), .A3(new_n1067), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G171), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1070), .A2(new_n1063), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G171), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(KEYINPUT54), .C1(G171), .C2(new_n1074), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1058), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT56), .B(G2072), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1000), .A2(new_n974), .A3(new_n1001), .A4(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n998), .B2(G1956), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n575), .A2(new_n1087), .A3(new_n581), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n575), .B2(new_n581), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1083), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1085), .B(new_n1090), .C1(new_n998), .C2(G1956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT120), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1092), .A2(new_n1096), .A3(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1996), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1000), .A2(new_n1102), .A3(new_n974), .A4(new_n1001), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n979), .B2(new_n972), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1101), .B(new_n850), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1101), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(new_n557), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n979), .A2(new_n972), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n729), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n998), .B2(G1348), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n614), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1113), .B(new_n613), .C1(new_n998), .C2(G1348), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1012), .A2(new_n713), .B1(new_n729), .B2(new_n1112), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(new_n1111), .A3(new_n614), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1110), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n996), .A2(new_n997), .ZN(new_n1122));
  AOI21_X1  g697(.A(G1956), .B1(new_n1122), .B2(new_n1000), .ZN(new_n1123));
  AND4_X1   g698(.A1(new_n1000), .A2(new_n974), .A3(new_n1001), .A4(new_n1084), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT118), .B(new_n1091), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1083), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1093), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT119), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1093), .A2(new_n1129), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1012), .A2(new_n705), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1090), .B1(new_n1133), .B2(new_n1085), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1135), .A2(new_n1126), .A3(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1098), .B(new_n1121), .C1(new_n1131), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1093), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1128), .B1(new_n1139), .B2(new_n1115), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1082), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1034), .A2(new_n1045), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1051), .A2(new_n1047), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1075), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1022), .B1(new_n1142), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1034), .A2(new_n1045), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1144), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1003), .A2(new_n993), .A3(G286), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1147), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1156), .A2(KEYINPUT116), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1156), .B2(KEYINPUT116), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1147), .A2(new_n1143), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1045), .A2(new_n1029), .A3(new_n798), .ZN(new_n1162));
  NOR2_X1   g737(.A1(G305), .A2(G1981), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT115), .Z(new_n1164));
  AOI21_X1  g739(.A(new_n1027), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1145), .A2(new_n1147), .A3(KEYINPUT62), .A4(new_n1146), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1022), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1160), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n991), .B1(new_n1152), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n825), .A2(new_n828), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT125), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n1172), .A2(new_n984), .B1(G2067), .B2(new_n724), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n987), .A2(new_n980), .ZN(new_n1174));
  XOR2_X1   g749(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1175));
  XNOR2_X1  g750(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1173), .A2(new_n980), .B1(new_n986), .B2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n974), .A2(new_n979), .A3(G1996), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1178), .A2(KEYINPUT46), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n980), .B1(new_n981), .B2(new_n878), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(KEYINPUT46), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT47), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1177), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n970), .B1(new_n1170), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1184), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1148), .A2(KEYINPUT62), .A3(new_n1021), .A4(new_n1020), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1187), .B(new_n1166), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1092), .A2(new_n1096), .A3(new_n1093), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1096), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(KEYINPUT60), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1192), .A2(new_n1194), .A3(new_n1119), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1127), .A2(KEYINPUT119), .A3(new_n1130), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1136), .B1(new_n1135), .B2(new_n1126), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1140), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1150), .B1(new_n1200), .B2(new_n1082), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1188), .B1(new_n1201), .B2(new_n1022), .ZN(new_n1202));
  OAI211_X1 g777(.A(KEYINPUT127), .B(new_n1186), .C1(new_n1202), .C2(new_n991), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1185), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g779(.A1(new_n900), .A2(new_n901), .ZN(new_n1206));
  NOR4_X1   g780(.A1(G401), .A2(G229), .A3(new_n461), .A4(G227), .ZN(new_n1207));
  AND3_X1   g781(.A1(new_n1206), .A2(new_n960), .A3(new_n1207), .ZN(G308));
  NAND3_X1  g782(.A1(new_n1206), .A2(new_n960), .A3(new_n1207), .ZN(G225));
endmodule


