//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  INV_X1    g0003(.A(G244), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G50), .B2(G226), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n205), .B(new_n217), .C1(G116), .C2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(KEYINPUT1), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OR3_X1    g0022(.A1(new_n218), .A2(KEYINPUT1), .A3(new_n221), .ZN(new_n223));
  INV_X1    g0023(.A(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n215), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n230), .A2(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(KEYINPUT64), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n231), .A2(G50), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  OR3_X1    g0034(.A1(new_n233), .A2(new_n220), .A3(new_n234), .ZN(new_n235));
  AND4_X1   g0035(.A1(new_n222), .A2(new_n223), .A3(new_n228), .A4(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT67), .B(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n249), .B(KEYINPUT68), .Z(new_n250));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G274), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT69), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G222), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G223), .A2(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n234), .B1(G33), .B2(G41), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n268), .B(new_n269), .C1(G77), .C2(new_n264), .ZN(new_n270));
  INV_X1    g0070(.A(G226), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n257), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n259), .B(new_n270), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G200), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  OAI21_X1  g0076(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n220), .A2(G33), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n277), .B1(new_n278), .B2(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n234), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n219), .B2(G20), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n283), .A2(new_n285), .B1(G50), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n219), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G50), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n287), .B(new_n291), .C1(KEYINPUT71), .C2(KEYINPUT9), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(KEYINPUT71), .B2(KEYINPUT9), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n287), .A2(new_n291), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n294), .A2(KEYINPUT71), .A3(KEYINPUT9), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n275), .B1(new_n276), .B2(new_n274), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n274), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n294), .C1(G179), .C2(new_n274), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n271), .A2(new_n265), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n264), .B(new_n302), .C1(G232), .C2(new_n265), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G97), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT72), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n303), .A2(KEYINPUT72), .A3(new_n304), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n269), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n272), .A2(G238), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n259), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n310), .B1(new_n309), .B2(new_n312), .ZN(new_n315));
  OAI21_X1  g0115(.A(G169), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT14), .ZN(new_n317));
  INV_X1    g0117(.A(new_n315), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n313), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT14), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(G169), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n317), .B(new_n321), .C1(new_n319), .C2(new_n322), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n280), .A2(new_n290), .B1(new_n220), .B2(G68), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n281), .A2(new_n203), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n285), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT11), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n286), .A2(G68), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT73), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n289), .A2(new_n215), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT12), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n327), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(G200), .B1(new_n314), .B2(new_n315), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n318), .A2(G190), .A3(new_n313), .ZN(new_n335));
  INV_X1    g0135(.A(new_n332), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n282), .A2(new_n289), .ZN(new_n339));
  INV_X1    g0139(.A(new_n286), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(new_n282), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  AND2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(G20), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n344), .B(KEYINPUT7), .C1(new_n345), .C2(G33), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT7), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n264), .B2(G20), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n215), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n229), .A2(new_n215), .ZN(new_n350));
  NOR2_X1   g0150(.A1(G58), .A2(G68), .ZN(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n279), .A2(G159), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n342), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n355), .A2(new_n285), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n260), .A2(KEYINPUT74), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT3), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n359), .A3(G33), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n220), .A3(new_n262), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT7), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n360), .A2(new_n347), .A3(new_n220), .A4(new_n262), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(G68), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n354), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(KEYINPUT16), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n341), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n272), .A2(G232), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n261), .A2(new_n207), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n265), .A2(G226), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n360), .B2(new_n262), .ZN(new_n371));
  NOR2_X1   g0171(.A1(G223), .A2(G1698), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n234), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n261), .B2(new_n255), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n259), .B(new_n368), .C1(new_n374), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G200), .ZN(new_n378));
  AOI211_X1 g0178(.A(new_n372), .B(new_n370), .C1(new_n360), .C2(new_n262), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n269), .B1(new_n379), .B2(new_n369), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n380), .A2(G190), .A3(new_n259), .A4(new_n368), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n367), .A2(KEYINPUT17), .A3(new_n378), .A4(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n366), .A2(new_n285), .A3(new_n355), .ZN(new_n383));
  INV_X1    g0183(.A(new_n341), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n383), .A2(new_n378), .A3(new_n381), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT17), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n355), .A2(new_n285), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n215), .B1(new_n361), .B2(KEYINPUT7), .ZN(new_n390));
  AOI211_X1 g0190(.A(new_n342), .B(new_n354), .C1(new_n390), .C2(new_n363), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n384), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n377), .A2(G169), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n380), .A2(G179), .A3(new_n259), .A4(new_n368), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT18), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n392), .A2(new_n395), .A3(KEYINPUT18), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(KEYINPUT75), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(new_n395), .A3(KEYINPUT18), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n388), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n265), .A2(G232), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n264), .B(new_n404), .C1(new_n216), .C2(new_n265), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(new_n269), .C1(G107), .C2(new_n264), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n259), .C1(new_n204), .C2(new_n273), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G200), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n282), .A2(new_n280), .B1(new_n220), .B2(new_n203), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT15), .B(G87), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(new_n281), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n285), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n289), .A2(new_n203), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n413), .C1(new_n203), .C2(new_n340), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n414), .A2(KEYINPUT70), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(KEYINPUT70), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n408), .B1(new_n276), .B2(new_n407), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n407), .A2(G179), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n407), .A2(new_n298), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(new_n414), .A3(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n301), .A2(new_n338), .A3(new_n403), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT79), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n360), .A2(new_n262), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n204), .A2(G1698), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT4), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(KEYINPUT3), .A2(G33), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n427), .B1(new_n343), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n426), .A2(new_n430), .B1(KEYINPUT4), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n264), .A2(G250), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G283), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(KEYINPUT78), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT78), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(G33), .B2(G283), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n434), .A2(new_n265), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n425), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n208), .B1(new_n262), .B2(new_n263), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n437), .A2(G33), .A3(G283), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n435), .A2(KEYINPUT78), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n441), .A2(G1698), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n429), .B1(new_n360), .B2(new_n262), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n428), .B1(new_n264), .B2(new_n427), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n444), .B(KEYINPUT79), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n269), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n256), .A2(G1), .ZN(new_n449));
  AND2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  NOR2_X1   g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G274), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n452), .A2(new_n376), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(G257), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n448), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n298), .ZN(new_n459));
  INV_X1    g0259(.A(new_n285), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n219), .A2(G33), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(KEYINPUT76), .A3(new_n288), .A4(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n288), .A2(new_n461), .A3(new_n234), .A4(new_n284), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT76), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G97), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n289), .A2(G97), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(KEYINPUT77), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT77), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n209), .B1(new_n462), .B2(new_n465), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(new_n468), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT6), .ZN(new_n475));
  INV_X1    g0275(.A(G107), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n209), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(G97), .A2(G107), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(KEYINPUT6), .A3(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n481), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n346), .A2(new_n348), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(new_n476), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n285), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n474), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n448), .A2(new_n322), .A3(new_n457), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n459), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT81), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT81), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n459), .A2(new_n490), .A3(new_n486), .A4(new_n487), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n448), .A2(G190), .A3(new_n457), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n470), .A2(new_n473), .B1(new_n484), .B2(new_n285), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G200), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n448), .B2(new_n457), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT80), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n458), .A2(G200), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT80), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n493), .A4(new_n492), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n489), .A2(new_n491), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT23), .B1(new_n220), .B2(G107), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT23), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n476), .A3(G20), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n502), .B(new_n504), .C1(new_n505), .C2(new_n281), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT83), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n261), .A2(G20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G116), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(KEYINPUT83), .A3(new_n504), .A4(new_n502), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n264), .A2(new_n220), .A3(G87), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT22), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n426), .A2(KEYINPUT22), .A3(new_n220), .A4(G87), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT24), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n512), .A2(new_n516), .A3(KEYINPUT24), .A4(new_n515), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n285), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n462), .A2(new_n465), .A3(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n289), .A2(new_n476), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n523), .B(KEYINPUT25), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n456), .A2(G264), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n360), .A2(new_n262), .B1(new_n210), .B2(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n208), .A2(new_n265), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n529), .B1(G33), .B2(G294), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n454), .B(new_n527), .C1(new_n530), .C2(new_n376), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n298), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(G179), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n289), .A2(new_n505), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n463), .A2(new_n505), .ZN(new_n536));
  AOI21_X1  g0336(.A(G20), .B1(new_n261), .B2(G97), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n438), .B2(new_n436), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n284), .A2(new_n234), .B1(G20), .B2(new_n505), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n538), .A2(KEYINPUT20), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT20), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n535), .B(new_n536), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n456), .A2(G270), .ZN(new_n543));
  INV_X1    g0343(.A(G303), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n264), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n265), .A2(G264), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n360), .B2(new_n262), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n210), .A2(new_n265), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n454), .B(new_n543), .C1(new_n549), .C2(new_n376), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n276), .ZN(new_n551));
  AOI211_X1 g0351(.A(new_n542), .B(new_n551), .C1(G200), .C2(new_n550), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(G169), .A3(new_n542), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT21), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n549), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n455), .B1(new_n556), .B2(new_n269), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n557), .A2(G179), .A3(new_n543), .A4(new_n542), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n550), .A2(new_n542), .A3(KEYINPUT21), .A4(G169), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n534), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n410), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n462), .A2(new_n465), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n288), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n220), .A2(new_n566), .B1(new_n478), .B2(new_n207), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT19), .B1(new_n509), .B2(G97), .ZN(new_n568));
  AOI21_X1  g0368(.A(G20), .B1(new_n360), .B2(new_n262), .ZN(new_n569));
  AOI211_X1 g0369(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(G68), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n563), .B(new_n565), .C1(new_n570), .C2(new_n460), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n376), .B1(G250), .B2(new_n449), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n256), .A2(G1), .A3(G274), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n261), .A2(new_n505), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n360), .A2(new_n262), .B1(new_n216), .B2(new_n265), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n204), .A2(G1698), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n322), .B(new_n574), .C1(new_n578), .C2(new_n376), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n216), .A2(new_n265), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n426), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n575), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n376), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n572), .A2(new_n573), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n298), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n571), .A2(new_n579), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G200), .B1(new_n583), .B2(new_n584), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n426), .A2(new_n220), .A3(G68), .ZN(new_n588));
  INV_X1    g0388(.A(new_n567), .ZN(new_n589));
  INV_X1    g0389(.A(new_n568), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n564), .B1(new_n591), .B2(new_n285), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n462), .A2(new_n465), .A3(G87), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT82), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n462), .A2(new_n465), .A3(KEYINPUT82), .A4(G87), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(G190), .B(new_n574), .C1(new_n578), .C2(new_n376), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n587), .A2(new_n592), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n586), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n531), .A2(G200), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n526), .B(new_n601), .C1(new_n276), .C2(new_n531), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n501), .A2(new_n561), .A3(new_n600), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n424), .A2(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n420), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n337), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n388), .B1(new_n333), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n392), .A2(new_n395), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT18), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n399), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n297), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(new_n300), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT84), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n560), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n555), .A2(new_n558), .A3(KEYINPUT84), .A4(new_n559), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n526), .A2(new_n533), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n501), .A2(new_n620), .A3(new_n600), .A4(new_n602), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n489), .A2(new_n491), .A3(new_n600), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n448), .A2(new_n322), .A3(new_n457), .ZN(new_n624));
  AOI21_X1  g0424(.A(G169), .B1(new_n448), .B2(new_n457), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(new_n600), .A3(new_n627), .A4(new_n486), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n623), .A2(new_n586), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n614), .B1(new_n424), .B2(new_n630), .ZN(G369));
  NOR2_X1   g0431(.A1(new_n224), .A2(G20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n234), .ZN(new_n633));
  OR3_X1    g0433(.A1(new_n633), .A2(KEYINPUT85), .A3(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT85), .B1(new_n633), .B2(KEYINPUT27), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(G213), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT86), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(KEYINPUT86), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G343), .ZN(new_n641));
  INV_X1    g0441(.A(new_n542), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT87), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(new_n552), .ZN(new_n645));
  INV_X1    g0445(.A(new_n644), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n645), .A2(new_n560), .B1(new_n618), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G330), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n641), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n619), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n602), .B1(new_n526), .B2(new_n641), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n619), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n560), .A2(new_n641), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(new_n651), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n655), .A2(new_n658), .ZN(G399));
  NOR2_X1   g0459(.A1(new_n225), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n478), .A2(new_n207), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G116), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(G1), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n233), .B2(new_n661), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT88), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT28), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n641), .B1(new_n621), .B2(new_n629), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT29), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n501), .A2(new_n620), .A3(new_n600), .A4(new_n602), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n628), .A2(new_n586), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(KEYINPUT26), .B2(new_n622), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n650), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT90), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n670), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n586), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n489), .A2(new_n491), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n497), .A2(new_n500), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n679), .A2(new_n602), .A3(new_n680), .A4(new_n600), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n534), .A2(new_n560), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n678), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n622), .A2(new_n627), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT91), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n626), .A2(new_n600), .A3(new_n486), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT26), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n622), .A2(KEYINPUT91), .A3(new_n627), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n650), .B1(new_n684), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT29), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n677), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT89), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(KEYINPUT30), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n527), .B1(new_n530), .B2(new_n376), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n557), .A3(G179), .A4(new_n543), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n583), .A2(new_n584), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n448), .A2(new_n457), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n696), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n448), .A2(new_n457), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n697), .A2(new_n550), .A3(new_n322), .ZN(new_n704));
  INV_X1    g0504(.A(new_n696), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n703), .A2(new_n704), .A3(new_n700), .A4(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n458), .A2(new_n322), .A3(new_n531), .A4(new_n550), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n702), .B(new_n706), .C1(new_n700), .C2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n708), .A2(new_n709), .A3(new_n650), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n708), .B2(new_n650), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n603), .A2(new_n650), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n694), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n667), .B1(new_n715), .B2(G1), .ZN(G364));
  NOR2_X1   g0516(.A1(G13), .A2(G33), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n647), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(G355), .B(KEYINPUT92), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n226), .A3(new_n264), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n253), .A2(new_n256), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n426), .A2(new_n225), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G45), .B2(new_n233), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n723), .B1(G116), .B2(new_n226), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n234), .B1(G20), .B2(new_n298), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n719), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n632), .A2(G45), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n661), .A2(G1), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(G20), .A2(G179), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT93), .Z(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n276), .A3(G200), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT96), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(KEYINPUT33), .B(G317), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n276), .A2(new_n495), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(KEYINPUT97), .B(G326), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n740), .A2(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G283), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n276), .A2(G20), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT95), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n322), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n495), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n276), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n735), .A2(new_n754), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n746), .B1(new_n747), .B2(new_n752), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n735), .A2(new_n276), .A3(new_n495), .ZN(new_n757));
  INV_X1    g0557(.A(G311), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n220), .B1(new_n754), .B2(new_n322), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n264), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n742), .A2(G20), .A3(new_n322), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n544), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT98), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n750), .A2(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G329), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR4_X1   g0570(.A1(new_n756), .A2(new_n759), .A3(new_n762), .A4(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n760), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n740), .A2(G68), .B1(G97), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n763), .B1(new_n744), .B2(G50), .ZN(new_n774));
  INV_X1    g0574(.A(new_n764), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G87), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n751), .A2(G107), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n773), .A2(new_n774), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n768), .A2(KEYINPUT32), .A3(new_n779), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n757), .A2(new_n203), .B1(new_n755), .B2(new_n229), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT32), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n767), .B2(G159), .ZN(new_n784));
  NOR4_X1   g0584(.A1(new_n778), .A2(new_n780), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n728), .B1(new_n771), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n721), .A2(new_n730), .A3(new_n733), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n647), .A2(G330), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(new_n648), .A3(new_n732), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n789), .ZN(G396));
  AND2_X1   g0590(.A1(new_n670), .A2(new_n676), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n650), .A2(new_n414), .ZN(new_n792));
  AND3_X1   g0592(.A1(new_n421), .A2(KEYINPUT99), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(KEYINPUT99), .B1(new_n421), .B2(new_n792), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n793), .A2(new_n794), .B1(new_n420), .B2(new_n641), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n791), .A2(new_n796), .B1(new_n675), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(KEYINPUT100), .B2(new_n714), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n713), .B(KEYINPUT100), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n732), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n740), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n802), .A2(new_n747), .B1(new_n544), .B2(new_n743), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n760), .A2(new_n209), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n752), .A2(new_n207), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n763), .B1(new_n476), .B2(new_n764), .C1(new_n757), .C2(new_n505), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n807), .B1(new_n761), .B2(new_n755), .C1(new_n758), .C2(new_n768), .ZN(new_n808));
  INV_X1    g0608(.A(new_n755), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n740), .A2(G150), .B1(G143), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n811), .B2(new_n743), .C1(new_n779), .C2(new_n757), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n751), .A2(G68), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n229), .C2(new_n760), .ZN(new_n815));
  INV_X1    g0615(.A(new_n426), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n767), .B2(G132), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n290), .B2(new_n764), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n808), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n728), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n796), .A2(new_n717), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n728), .A2(new_n717), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n203), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n733), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n801), .A2(new_n824), .ZN(G384));
  NAND2_X1  g0625(.A1(new_n392), .A2(new_n640), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n826), .A2(new_n608), .A3(new_n827), .A4(new_n385), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n366), .A2(new_n285), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT16), .B1(new_n364), .B2(new_n365), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n384), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n395), .B2(new_n640), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n832), .A2(new_n385), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n828), .B1(new_n833), .B2(new_n827), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n640), .ZN(new_n835));
  OAI211_X1 g0635(.A(KEYINPUT38), .B(new_n834), .C1(new_n402), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT38), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n392), .A2(new_n395), .A3(KEYINPUT75), .A4(KEYINPUT18), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n401), .A2(new_n610), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n385), .B(KEYINPUT17), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n828), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n827), .B1(new_n832), .B2(new_n385), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n837), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n836), .A2(new_n845), .A3(KEYINPUT103), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n841), .A2(new_n844), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT103), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n333), .B(new_n337), .C1(new_n336), .C2(new_n641), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n323), .A2(new_n332), .A3(new_n650), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n712), .A3(new_n795), .ZN(new_n854));
  OR3_X1    g0654(.A1(new_n850), .A2(new_n854), .A3(KEYINPUT40), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n826), .A2(new_n608), .A3(new_n385), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(new_n827), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n826), .B1(new_n840), .B2(new_n611), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n837), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n836), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT40), .B1(new_n854), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n423), .A2(new_n712), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT104), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n862), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(G330), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n846), .A2(KEYINPUT39), .A3(new_n849), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n333), .A2(new_n650), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n640), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n612), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n850), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n641), .B(new_n797), .C1(new_n621), .C2(new_n629), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n650), .A2(new_n420), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n876), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n875), .A2(new_n882), .A3(new_n853), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n872), .A2(new_n874), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n866), .B(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n677), .A2(new_n423), .A3(new_n693), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n614), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n885), .B(new_n887), .Z(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n219), .B2(new_n632), .ZN(new_n889));
  OAI21_X1  g0689(.A(G77), .B1(new_n229), .B2(new_n215), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n233), .A2(new_n890), .B1(G50), .B2(new_n215), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(G1), .A3(new_n224), .ZN(new_n892));
  OAI211_X1 g0692(.A(G20), .B(new_n375), .C1(new_n481), .C2(KEYINPUT35), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n505), .B(new_n893), .C1(KEYINPUT35), .C2(new_n481), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT101), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT36), .Z(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(new_n892), .A3(new_n896), .ZN(G367));
  OAI22_X1  g0697(.A1(new_n752), .A2(new_n203), .B1(new_n229), .B2(new_n764), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n760), .A2(new_n215), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n744), .A2(G143), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n264), .B1(new_n755), .B2(new_n278), .C1(new_n290), .C2(new_n757), .ZN(new_n901));
  NOR4_X1   g0701(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n902), .B1(new_n811), .B2(new_n768), .C1(new_n779), .C2(new_n802), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n740), .A2(G294), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n809), .A2(G303), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n775), .A2(KEYINPUT46), .A3(G116), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n757), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(G283), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n751), .A2(G97), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT46), .B1(new_n775), .B2(G116), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n744), .B2(G311), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n767), .A2(G317), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n909), .A2(new_n910), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n816), .B1(new_n476), .B2(new_n760), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n903), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT47), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n728), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n592), .A2(new_n597), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n650), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n600), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n586), .B2(new_n920), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n922), .A2(new_n720), .ZN(new_n923));
  INV_X1    g0723(.A(new_n725), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n729), .B1(new_n226), .B2(new_n410), .C1(new_n240), .C2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n918), .A2(new_n733), .A3(new_n923), .A4(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n501), .B1(new_n493), .B2(new_n641), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n650), .A2(new_n626), .A3(new_n486), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n658), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT44), .Z(new_n933));
  NOR2_X1   g0733(.A1(new_n658), .A2(new_n931), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n655), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n653), .B(new_n656), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n648), .B(new_n938), .Z(new_n939));
  AND2_X1   g0739(.A1(new_n715), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n654), .A3(new_n935), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n715), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n660), .B(KEYINPUT41), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n731), .A2(G1), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n657), .A2(new_n930), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT105), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n679), .B1(new_n931), .B2(new_n619), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n954), .A2(new_n641), .B1(new_n949), .B2(KEYINPUT42), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT106), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n654), .A2(new_n931), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n953), .B1(new_n952), .B2(new_n955), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n958), .B1(new_n957), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n927), .B1(new_n948), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(G387));
  INV_X1    g0766(.A(new_n728), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n740), .A2(G311), .B1(G317), .B2(new_n809), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n544), .B2(new_n757), .C1(new_n753), .C2(new_n743), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT48), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n747), .B2(new_n760), .C1(new_n761), .C2(new_n764), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n971), .A2(new_n972), .B1(G116), .B2(new_n751), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n767), .A2(new_n745), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n973), .A2(new_n974), .A3(new_n816), .A4(new_n975), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n910), .B1(new_n215), .B2(new_n757), .C1(new_n768), .C2(new_n278), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n426), .B1(new_n779), .B2(new_n743), .C1(new_n802), .C2(new_n282), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(new_n562), .C2(new_n772), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n290), .B2(new_n755), .C1(new_n203), .C2(new_n764), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n967), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n282), .A2(KEYINPUT50), .A3(G50), .ZN(new_n982));
  INV_X1    g0782(.A(new_n663), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(G68), .A2(G77), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT50), .B1(new_n282), .B2(G50), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n984), .A2(new_n256), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n725), .B(new_n987), .C1(new_n245), .C2(new_n256), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n226), .A3(new_n264), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G107), .C2(new_n226), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT107), .Z(new_n991));
  AOI211_X1 g0791(.A(new_n732), .B(new_n981), .C1(new_n729), .C2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n653), .A2(new_n720), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n992), .A2(new_n993), .B1(new_n946), .B2(new_n939), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n660), .B1(new_n715), .B2(new_n939), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n940), .B2(new_n995), .ZN(G393));
  NAND3_X1  g0796(.A1(new_n936), .A2(KEYINPUT109), .A3(new_n655), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n937), .A2(new_n941), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n998), .B2(KEYINPUT109), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n942), .B(new_n660), .C1(new_n999), .C2(new_n940), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n946), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n930), .A2(new_n720), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT110), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n729), .B1(new_n209), .B2(new_n226), .C1(new_n924), .C2(new_n249), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT111), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n767), .A2(G143), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n203), .B2(new_n760), .C1(new_n282), .C2(new_n757), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n764), .A2(new_n215), .ZN(new_n1008));
  NOR4_X1   g0808(.A1(new_n1007), .A2(new_n816), .A3(new_n805), .A4(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n278), .A2(new_n743), .B1(new_n755), .B2(new_n779), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT51), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(new_n290), .C2(new_n802), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT112), .Z(new_n1013));
  AOI22_X1  g0813(.A1(G311), .A2(new_n809), .B1(new_n744), .B2(G317), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n763), .B1(new_n747), .B2(new_n764), .C1(new_n768), .C2(new_n753), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n777), .B1(new_n761), .B2(new_n757), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n505), .B2(new_n760), .C1(new_n544), .C2(new_n802), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n967), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  OR4_X1    g0821(.A1(new_n732), .A2(new_n1003), .A3(new_n1005), .A4(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1000), .A2(new_n1001), .A3(new_n1022), .ZN(G390));
  NAND3_X1  g0823(.A1(new_n423), .A2(G330), .A3(new_n712), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n886), .A2(new_n614), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT115), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT115), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n886), .A2(new_n1027), .A3(new_n614), .A4(new_n1024), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n871), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n860), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n877), .B1(new_n692), .B2(new_n797), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n851), .A2(KEYINPUT114), .A3(new_n852), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT114), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n641), .A2(new_n336), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n337), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n323), .C2(new_n332), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n852), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1034), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1033), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1030), .B(new_n1031), .C1(new_n1032), .C2(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n867), .A2(new_n869), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n853), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n880), .B1(new_n675), .B2(new_n797), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n879), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1042), .B1(new_n1045), .B2(new_n871), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n853), .A2(new_n712), .A3(G330), .A4(new_n795), .ZN(new_n1047));
  AND3_X1   g0847(.A1(new_n1041), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1047), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n712), .A2(G330), .A3(new_n795), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1040), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1032), .A2(new_n1047), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1043), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n1047), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1055), .A2(KEYINPUT116), .A3(new_n882), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT116), .B1(new_n1055), .B2(new_n882), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1029), .A2(new_n1050), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1047), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n622), .A2(KEYINPUT91), .A3(new_n627), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT91), .B1(new_n622), .B2(new_n627), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n689), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n501), .A2(new_n600), .A3(new_n602), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n586), .B1(new_n1066), .B2(new_n682), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n641), .B(new_n797), .C1(new_n1065), .C2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n877), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1040), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1070), .A2(new_n871), .A3(new_n860), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n882), .A2(new_n853), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n870), .B1(new_n1072), .B2(new_n1030), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1061), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1041), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1060), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1059), .A2(new_n660), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1074), .A2(new_n946), .A3(new_n1075), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT119), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1042), .A2(new_n717), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n822), .A2(new_n282), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n763), .B1(new_n743), .B2(new_n747), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n814), .B1(new_n505), .B2(new_n755), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(new_n740), .C2(G107), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n908), .A2(G97), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G77), .A2(new_n772), .B1(new_n775), .B2(G87), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n767), .A2(G294), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n752), .A2(new_n290), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n767), .A2(G125), .B1(G159), .B2(new_n772), .ZN(new_n1091));
  XOR2_X1   g0891(.A(KEYINPUT54), .B(G143), .Z(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n264), .C1(new_n757), .C2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1090), .B(new_n1094), .C1(G132), .C2(new_n809), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n744), .A2(G128), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n811), .C2(new_n802), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n764), .A2(new_n278), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT117), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT53), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1089), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT118), .Z(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n728), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1081), .A2(new_n733), .A3(new_n1082), .A4(new_n1103), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1079), .A2(new_n1080), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1080), .B1(new_n1079), .B2(new_n1104), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(KEYINPUT120), .B1(new_n1078), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1059), .A2(new_n660), .A3(new_n1077), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT120), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(new_n1106), .C2(new_n1105), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(G378));
  INV_X1    g0912(.A(G330), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n855), .B2(new_n861), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n297), .A2(new_n300), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1117), .B1(new_n297), .B2(new_n300), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n640), .A2(new_n294), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1121), .B(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1045), .A2(new_n875), .B1(new_n612), .B2(new_n873), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n872), .ZN(new_n1126));
  AND4_X1   g0926(.A1(new_n872), .A2(new_n1124), .A3(new_n874), .A4(new_n883), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1115), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1124), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n884), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1125), .A2(new_n872), .A3(new_n1124), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n1114), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1128), .A2(KEYINPUT57), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(KEYINPUT121), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT121), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1026), .A2(new_n1136), .A3(new_n1028), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1133), .B1(new_n1138), .B2(new_n1059), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT122), .B1(new_n1139), .B2(new_n661), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1026), .A2(new_n1136), .A3(new_n1028), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1136), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1141), .A2(new_n1142), .B1(new_n1060), .B2(new_n1076), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1133), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT122), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n1146), .A3(new_n660), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT57), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1140), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1124), .A2(new_n717), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n752), .A2(new_n229), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n740), .A2(G97), .B1(G283), .B2(new_n767), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n505), .B2(new_n743), .C1(new_n410), .C2(new_n757), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G107), .C2(new_n809), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n360), .A2(new_n255), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1158), .B(new_n899), .C1(G77), .C2(new_n775), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n262), .A3(new_n1159), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT58), .Z(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n290), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n757), .A2(new_n811), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G125), .A2(new_n744), .B1(new_n809), .B2(G128), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n278), .B2(new_n760), .C1(new_n764), .C2(new_n1093), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G132), .C2(new_n740), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT59), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G33), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(G41), .B1(new_n767), .B2(G124), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n779), .C2(new_n752), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1162), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n728), .B1(new_n1161), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n822), .A2(new_n290), .ZN(new_n1174));
  AND4_X1   g0974(.A1(new_n733), .A2(new_n1153), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1148), .B2(new_n946), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1152), .A2(new_n1176), .ZN(G375));
  NAND2_X1  g0977(.A1(new_n1040), .A2(new_n717), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n822), .A2(new_n215), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1154), .A2(new_n816), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT123), .Z(new_n1181));
  AOI22_X1  g0981(.A1(new_n740), .A2(new_n1092), .B1(G50), .B2(new_n772), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n767), .A2(G128), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n755), .A2(new_n811), .B1(new_n779), .B2(new_n764), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G132), .B2(new_n744), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n757), .A2(new_n278), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n752), .A2(new_n203), .B1(new_n209), .B2(new_n764), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G303), .B2(new_n767), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n744), .A2(G294), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n264), .B1(new_n772), .B2(new_n562), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n740), .A2(G116), .B1(G283), .B2(new_n809), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n757), .A2(new_n476), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n1186), .A2(new_n1187), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n728), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1178), .A2(new_n733), .A3(new_n1179), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1053), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1055), .A2(new_n882), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT116), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1055), .A2(KEYINPUT116), .A3(new_n882), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1198), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1197), .B1(new_n1203), .B2(new_n947), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT124), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT124), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1206), .B(new_n1197), .C1(new_n1203), .C2(new_n947), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1134), .A2(new_n1203), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(new_n944), .A3(new_n1060), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(G381));
  NAND4_X1  g1011(.A1(new_n965), .A2(new_n1001), .A3(new_n1022), .A4(new_n1000), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1212), .A2(G396), .A3(G393), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G381), .A2(G384), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1109), .A2(new_n1079), .A3(new_n1104), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(G375), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(G407));
  INV_X1    g1017(.A(G343), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  NAND3_X1  g1020(.A1(new_n1152), .A2(G378), .A3(new_n1176), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1215), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n944), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1176), .B1(new_n1149), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1221), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1218), .A2(G213), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1058), .B1(new_n1028), .B2(new_n1026), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n660), .B(new_n1060), .C1(new_n1229), .C2(KEYINPUT60), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1209), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1208), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(G384), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1208), .B(G384), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1218), .A2(G213), .A3(G2897), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1235), .A2(KEYINPUT125), .A3(new_n1236), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT125), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1239), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1228), .A2(new_n1240), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1226), .A2(new_n1227), .A3(new_n1243), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT62), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT62), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1226), .A2(new_n1243), .A3(new_n1249), .A4(new_n1227), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1245), .A2(new_n1247), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  XOR2_X1   g1051(.A(G393), .B(G396), .Z(new_n1252));
  AND2_X1   g1052(.A1(new_n1252), .A2(KEYINPUT126), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n948), .A2(new_n964), .ZN(new_n1254));
  OAI21_X1  g1054(.A(G390), .B1(new_n1254), .B2(new_n927), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1255), .B2(new_n1212), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1255), .A2(new_n1212), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1252), .B(KEYINPUT126), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1251), .A2(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1226), .A2(new_n1227), .B1(new_n1243), .B2(new_n1239), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1240), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1258), .A2(new_n1212), .A3(new_n1255), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1257), .B2(new_n1253), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT63), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1246), .A2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1226), .A2(KEYINPUT63), .A3(new_n1243), .A4(new_n1227), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1262), .A2(new_n1264), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1260), .A2(new_n1268), .ZN(G405));
  AND3_X1   g1069(.A1(new_n1152), .A2(G378), .A3(new_n1176), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1215), .B1(new_n1152), .B2(new_n1176), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1270), .A2(new_n1271), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G375), .A2(new_n1222), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1238), .A3(new_n1221), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT127), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n1264), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1243), .B1(new_n1221), .B2(new_n1273), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1270), .A2(new_n1271), .A3(new_n1237), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT127), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1259), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1278), .A2(new_n1283), .ZN(G402));
endmodule


