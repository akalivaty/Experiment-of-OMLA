//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT1), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G127gat), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G134gat), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT66), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT66), .B1(new_n208), .B2(new_n210), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT67), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n206), .B(new_n215), .C1(new_n211), .C2(new_n212), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n208), .A2(new_n210), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT68), .B(G120gat), .Z(new_n219));
  OAI211_X1 g018(.A(new_n218), .B(new_n205), .C1(new_n219), .C2(new_n203), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT27), .B(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT28), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G169gat), .ZN(new_n231));
  INV_X1    g030(.A(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n230), .B1(KEYINPUT26), .B2(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(KEYINPUT26), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n234), .A2(new_n235), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT28), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n228), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G190gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT23), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(G169gat), .B2(G176gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n246), .A3(new_n229), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n244), .A2(new_n246), .A3(new_n249), .A4(new_n229), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n251), .B(new_n250), .C1(new_n243), .C2(new_n247), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n221), .A2(new_n238), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n255), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(new_n217), .A3(new_n220), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G227gat), .ZN(new_n260));
  INV_X1    g059(.A(G233gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n202), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n259), .A2(new_n202), .A3(new_n263), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n256), .A2(new_n258), .A3(new_n262), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT33), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G15gat), .B(G43gat), .Z(new_n270));
  XNOR2_X1  g069(.A(G71gat), .B(G99gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n265), .B(new_n266), .C1(new_n269), .C2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n267), .B2(new_n268), .ZN(new_n275));
  INV_X1    g074(.A(new_n266), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(new_n264), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n267), .A2(KEYINPUT32), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n278), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT36), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT78), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT70), .B(KEYINPUT29), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287));
  INV_X1    g086(.A(G211gat), .ZN(new_n288));
  INV_X1    g087(.A(G218gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n287), .B1(KEYINPUT22), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G211gat), .B(G218gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n286), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n293), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n292), .B(new_n287), .C1(KEYINPUT22), .C2(new_n290), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(KEYINPUT77), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT3), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G141gat), .B(G148gat), .Z(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  INV_X1    g101(.A(G162gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT2), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(KEYINPUT74), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G155gat), .B(G162gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n301), .A2(KEYINPUT74), .A3(new_n306), .A4(new_n304), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n284), .B1(new_n300), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n285), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n297), .A2(new_n298), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n299), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n285), .B1(new_n297), .B2(KEYINPUT77), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n308), .A2(new_n309), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(KEYINPUT78), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n311), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G228gat), .A2(G233gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n315), .A2(KEYINPUT29), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n324), .A2(KEYINPUT79), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n312), .B1(new_n324), .B2(KEYINPUT79), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n323), .B1(new_n314), .B2(new_n315), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n322), .A2(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G22gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n329), .A2(new_n330), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n329), .B2(new_n330), .ZN(new_n335));
  XNOR2_X1  g134(.A(G78gat), .B(G106gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT31), .B(G50gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI22_X1  g138(.A1(new_n332), .A2(new_n333), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n329), .A2(new_n330), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n341), .A2(new_n334), .A3(new_n331), .A4(new_n338), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n221), .A2(new_n320), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n217), .A2(new_n310), .A3(new_n220), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT5), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT75), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n221), .A2(new_n313), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n217), .A2(new_n310), .A3(KEYINPUT4), .A4(new_n220), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n351), .A2(new_n353), .A3(new_n344), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n344), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n217), .A2(new_n310), .A3(new_n220), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n310), .B1(new_n217), .B2(new_n220), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT5), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n349), .A2(new_n355), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n353), .A2(new_n344), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n351), .A2(new_n364), .A3(new_n354), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n351), .B2(new_n354), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n363), .B(new_n348), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT0), .ZN(new_n370));
  XNOR2_X1  g169(.A(G57gat), .B(G85gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n362), .A2(new_n372), .A3(new_n367), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n368), .A2(KEYINPUT6), .A3(new_n373), .ZN(new_n378));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n238), .A2(new_n255), .A3(KEYINPUT69), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT69), .B1(new_n238), .B2(new_n255), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n380), .B1(new_n383), .B2(new_n285), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT71), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n257), .B2(new_n380), .ZN(new_n386));
  AOI211_X1 g185(.A(KEYINPUT71), .B(new_n379), .C1(new_n238), .C2(new_n255), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n315), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT69), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n257), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT72), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n238), .A2(new_n255), .A3(KEYINPUT69), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n380), .A4(new_n393), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n381), .A2(new_n382), .A3(new_n379), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n238), .B2(new_n255), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT72), .B1(new_n396), .B2(new_n380), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n297), .A2(new_n298), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G8gat), .B(G36gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  NAND3_X1  g202(.A1(new_n389), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n384), .B2(new_n388), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n398), .A2(new_n315), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT37), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT37), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n400), .A3(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n403), .B(KEYINPUT73), .Z(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n411), .A2(KEYINPUT38), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n377), .A2(new_n378), .A3(new_n404), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT82), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT83), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n408), .B1(new_n389), .B2(new_n400), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(new_n403), .ZN(new_n419));
  INV_X1    g218(.A(new_n403), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n257), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n392), .B1(new_n422), .B2(new_n379), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n391), .A2(new_n380), .A3(new_n393), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n315), .B1(new_n425), .B2(new_n394), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n391), .A2(new_n285), .A3(new_n393), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n379), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n386), .A2(new_n387), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n399), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT83), .B(new_n420), .C1(new_n431), .C2(new_n408), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n419), .A2(new_n432), .A3(new_n409), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT38), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n412), .B1(new_n431), .B2(new_n408), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n435), .A2(new_n407), .B1(new_n431), .B2(new_n403), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n378), .A4(new_n377), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n416), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n345), .A2(new_n344), .A3(new_n346), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n441), .A2(KEYINPUT81), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(KEYINPUT81), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT39), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n353), .B1(new_n365), .B2(new_n366), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n356), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n447), .A3(new_n356), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n372), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n440), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n356), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(KEYINPUT39), .A3(new_n443), .A4(new_n442), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n452), .A2(KEYINPUT40), .A3(new_n372), .A4(new_n448), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n453), .A3(new_n374), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n410), .B1(new_n426), .B2(new_n430), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n404), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT30), .B1(new_n431), .B2(new_n403), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n343), .B1(new_n439), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n377), .A2(new_n378), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n459), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n340), .A2(new_n342), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n283), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n343), .A2(new_n281), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(new_n463), .A3(new_n470), .A4(new_n459), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n278), .B(new_n279), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(new_n459), .A3(new_n466), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT35), .B1(new_n473), .B2(new_n464), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G71gat), .B(G78gat), .Z(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G64gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G57gat), .ZN(new_n481));
  INV_X1    g280(.A(G57gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G64gat), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT91), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT91), .B1(new_n481), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n479), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n482), .A2(KEYINPUT93), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G57gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n493), .A3(G64gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n481), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n489), .A2(new_n479), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(new_n209), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n330), .A2(G15gat), .ZN(new_n503));
  INV_X1    g302(.A(G15gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G22gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n503), .B2(new_n505), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n508), .A2(new_n509), .A3(G1gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT88), .B1(new_n511), .B2(G1gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  INV_X1    g312(.A(G1gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT16), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n504), .A2(G22gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n330), .A2(G15gat), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT87), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n516), .B1(new_n519), .B2(new_n507), .ZN(new_n520));
  OAI21_X1  g319(.A(G8gat), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n514), .A3(new_n507), .ZN(new_n522));
  INV_X1    g321(.A(G8gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n508), .A2(new_n509), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n522), .B(new_n523), .C1(new_n524), .C2(new_n516), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(KEYINPUT21), .B2(new_n497), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n502), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n302), .ZN(new_n530));
  XNOR2_X1  g329(.A(G183gat), .B(G211gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n528), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT99), .ZN(new_n534));
  INV_X1    g333(.A(G29gat), .ZN(new_n535));
  INV_X1    g334(.A(G36gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT14), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(G29gat), .B2(G36gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n540), .B1(G29gat), .B2(G36gat), .ZN(new_n541));
  INV_X1    g340(.A(G50gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(G43gat), .ZN(new_n543));
  INV_X1    g342(.A(G43gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G50gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n545), .A3(KEYINPUT15), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT85), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n540), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n537), .A2(new_n539), .A3(KEYINPUT85), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n544), .A2(G50gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n542), .A2(G43gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G29gat), .A2(G36gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n546), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n552), .A2(new_n558), .A3(KEYINPUT86), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT86), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n546), .A2(new_n557), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT15), .B1(new_n543), .B2(new_n545), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n537), .A2(new_n539), .A3(KEYINPUT85), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT85), .B1(new_n537), .B2(new_n539), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n560), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(KEYINPUT17), .B(new_n548), .C1(new_n559), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(KEYINPUT96), .A3(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(G85gat), .A3(G92gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT8), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(G99gat), .B2(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n573), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT98), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT98), .B1(new_n588), .B2(new_n583), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(new_n574), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n580), .B1(new_n593), .B2(new_n576), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n594), .A2(new_n573), .B1(new_n589), .B2(new_n587), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT86), .B1(new_n552), .B2(new_n558), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n563), .A2(new_n566), .A3(new_n560), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n547), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(KEYINPUT17), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n534), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n548), .B1(new_n559), .B2(new_n567), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n606), .A2(KEYINPUT99), .A3(new_n597), .A4(new_n568), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n604), .A2(new_n596), .B1(KEYINPUT41), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n608), .A2(new_n615), .A3(new_n611), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT95), .Z(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n615), .B1(new_n608), .B2(new_n611), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n621), .B1(new_n622), .B2(KEYINPUT100), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n614), .A2(new_n616), .A3(KEYINPUT100), .A4(new_n621), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n533), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI22_X1  g432(.A1(new_n490), .A2(new_n496), .B1(new_n591), .B2(new_n595), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT91), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n482), .A2(G64gat), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n480), .A2(G57gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT91), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n487), .B(KEYINPUT92), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n478), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n582), .A2(new_n590), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n594), .A2(new_n589), .A3(new_n587), .A4(new_n573), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n489), .A2(new_n495), .A3(new_n479), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n634), .A2(KEYINPUT101), .A3(new_n635), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n497), .A2(new_n596), .A3(KEYINPUT10), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n635), .A3(new_n647), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n633), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n634), .A2(new_n647), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n632), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n631), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n648), .A2(new_n649), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n632), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n656), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n661), .A3(new_n630), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n657), .A2(KEYINPUT102), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n664), .B(new_n631), .C1(new_n654), .C2(new_n656), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT90), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n604), .A2(new_n526), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n599), .A2(new_n600), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n669), .A2(new_n548), .A3(new_n521), .A4(new_n525), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(G229gat), .A2(G233gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT13), .Z(new_n673));
  AOI21_X1  g472(.A(new_n667), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  AOI211_X1 g474(.A(KEYINPUT90), .B(new_n675), .C1(new_n668), .C2(new_n670), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n526), .B1(new_n601), .B2(KEYINPUT17), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n606), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n679), .A2(KEYINPUT18), .A3(new_n672), .A4(new_n668), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n521), .A2(new_n525), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n568), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n672), .B(new_n668), .C1(new_n682), .C2(new_n602), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT18), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(G113gat), .B(G141gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G197gat), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT11), .B(G169gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT12), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n677), .A2(new_n680), .A3(new_n685), .A4(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n680), .B1(new_n674), .B2(new_n676), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT89), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n683), .A2(new_n693), .A3(new_n684), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n683), .B2(new_n684), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n690), .B(KEYINPUT84), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n691), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AND4_X1   g497(.A1(new_n477), .A2(new_n627), .A3(new_n666), .A4(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n464), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT103), .B(G1gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1324gat));
  XOR2_X1   g501(.A(KEYINPUT16), .B(G8gat), .Z(new_n703));
  AND3_X1   g502(.A1(new_n699), .A2(new_n465), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n523), .B1(new_n699), .B2(new_n465), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(KEYINPUT42), .B2(new_n704), .ZN(G1325gat));
  NAND3_X1  g506(.A1(new_n699), .A2(new_n504), .A3(new_n472), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n699), .A2(new_n282), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n709), .B2(new_n504), .ZN(G1326gat));
  NAND2_X1  g509(.A1(new_n699), .A2(new_n343), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NAND2_X1  g512(.A1(new_n624), .A2(new_n625), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n468), .B2(new_n476), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n528), .B(new_n532), .Z(new_n716));
  INV_X1    g515(.A(new_n698), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n663), .A2(new_n665), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n535), .A3(new_n464), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT45), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  INV_X1    g522(.A(new_n467), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n415), .A2(KEYINPUT82), .B1(new_n433), .B2(KEYINPUT38), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n460), .B1(new_n725), .B2(new_n438), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n726), .B2(new_n343), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n475), .B1(new_n727), .B2(new_n283), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n723), .B1(new_n728), .B2(new_n714), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n477), .A2(KEYINPUT44), .A3(new_n626), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(new_n719), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n732), .A2(new_n464), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n722), .B1(new_n733), .B2(new_n535), .ZN(G1328gat));
  AOI21_X1  g533(.A(new_n536), .B1(new_n732), .B2(new_n465), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n536), .A3(new_n465), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT46), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n735), .A2(new_n737), .ZN(G1329gat));
  NAND4_X1  g537(.A1(new_n731), .A2(G43gat), .A3(new_n282), .A4(new_n719), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n472), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n544), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g542(.A1(new_n729), .A2(new_n730), .A3(new_n343), .A4(new_n719), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n542), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n745), .B2(new_n744), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n720), .A2(new_n542), .A3(new_n343), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(KEYINPUT48), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(G50gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n748), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(G1331gat));
  NAND3_X1  g553(.A1(new_n627), .A2(new_n718), .A3(new_n717), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT105), .Z(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(new_n477), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n464), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n491), .A2(new_n493), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1332gat));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n756), .A2(new_n477), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT106), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n465), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT49), .B(G64gat), .Z(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(G1333gat));
  NAND4_X1  g567(.A1(new_n762), .A2(G71gat), .A3(new_n282), .A4(new_n764), .ZN(new_n769));
  INV_X1    g568(.A(G71gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n763), .B2(new_n281), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1334gat));
  NAND3_X1  g573(.A1(new_n762), .A2(new_n343), .A3(new_n764), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g575(.A1(new_n716), .A2(new_n698), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n666), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n731), .A2(new_n464), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n576), .B1(new_n780), .B2(KEYINPUT108), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(KEYINPUT108), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n715), .A2(new_n777), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(new_n576), .A3(new_n464), .A4(new_n718), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n786), .ZN(G1336gat));
  NAND3_X1  g586(.A1(new_n731), .A2(new_n465), .A3(new_n779), .ZN(new_n788));
  INV_X1    g587(.A(new_n593), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n459), .A2(G92gat), .A3(new_n666), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n795));
  AND4_X1   g594(.A1(new_n477), .A2(new_n626), .A3(new_n777), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n715), .B2(new_n777), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n788), .A2(new_n789), .B1(new_n798), .B2(new_n791), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n799), .B2(new_n793), .ZN(G1337gat));
  XNOR2_X1  g599(.A(KEYINPUT111), .B(G99gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n731), .A2(new_n282), .A3(new_n779), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(KEYINPUT110), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(KEYINPUT110), .B2(new_n802), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n785), .A2(new_n472), .A3(new_n718), .A4(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n466), .A2(G106gat), .A3(new_n666), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n785), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n729), .A2(new_n730), .A3(new_n343), .A4(new_n779), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G106gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n808), .B1(new_n796), .B2(new_n797), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT113), .B1(new_n815), .B2(KEYINPUT53), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817));
  AOI211_X1 g616(.A(new_n817), .B(new_n810), .C1(new_n812), .C2(new_n814), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n816), .B2(new_n818), .ZN(G1339gat));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n630), .B1(new_n654), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n650), .A2(new_n633), .A3(new_n653), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n660), .A2(new_n822), .A3(KEYINPUT54), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n662), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n660), .A2(new_n822), .A3(KEYINPUT54), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n631), .B1(new_n660), .B2(KEYINPUT54), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n698), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n685), .A2(new_n690), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n692), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n668), .A2(new_n670), .A3(new_n675), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n668), .A2(new_n670), .A3(KEYINPUT114), .A4(new_n675), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n672), .B1(new_n679), .B2(new_n668), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n689), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n678), .A2(new_n606), .B1(new_n604), .B2(new_n526), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n835), .B(new_n836), .C1(new_n672), .C2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(KEYINPUT115), .A3(new_n689), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n832), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n718), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n626), .B1(new_n830), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n825), .A2(new_n845), .A3(new_n829), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n714), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n533), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n716), .A2(new_n714), .A3(new_n666), .A4(new_n717), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n343), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n465), .A2(new_n463), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n281), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n717), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n853), .A2(new_n463), .A3(new_n473), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n203), .A3(new_n698), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT116), .ZN(G1340gat));
  OAI21_X1  g662(.A(G120gat), .B1(new_n858), .B2(new_n666), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(new_n219), .A3(new_n718), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1341gat));
  OAI21_X1  g665(.A(G127gat), .B1(new_n858), .B2(new_n533), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n860), .A2(new_n209), .A3(new_n716), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT117), .ZN(G1342gat));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n626), .A3(new_n857), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G134gat), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n860), .A2(new_n207), .A3(new_n626), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT56), .ZN(new_n876));
  OR3_X1    g675(.A1(new_n874), .A2(KEYINPUT119), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT119), .B1(new_n874), .B2(new_n876), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1343gat));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n852), .B2(new_n343), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n466), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n827), .B2(new_n828), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n821), .A2(KEYINPUT121), .A3(new_n823), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n826), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n698), .A3(new_n825), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n843), .A2(KEYINPUT115), .A3(new_n689), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT115), .B1(new_n843), .B2(new_n689), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n691), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n891), .B2(new_n666), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n718), .A2(new_n845), .A3(KEYINPUT120), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n887), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n849), .B1(new_n894), .B2(new_n714), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n851), .B1(new_n895), .B2(new_n716), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n880), .B1(new_n882), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n282), .A2(new_n856), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n698), .A2(G141gat), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n283), .A2(new_n343), .ZN(new_n903));
  NOR4_X1   g702(.A1(new_n853), .A2(new_n463), .A3(new_n903), .A4(new_n465), .ZN(new_n904));
  AOI21_X1  g703(.A(G141gat), .B1(new_n904), .B2(new_n698), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT122), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT58), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT122), .B(new_n908), .C1(new_n902), .C2(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1344gat));
  NOR4_X1   g709(.A1(new_n533), .A2(new_n626), .A3(new_n718), .A4(new_n698), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n714), .ZN(new_n912));
  INV_X1    g711(.A(new_n849), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n914), .B2(new_n533), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n881), .B1(new_n915), .B2(new_n466), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n852), .A2(new_n882), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n898), .A2(new_n718), .ZN(new_n920));
  OAI211_X1 g719(.A(KEYINPUT59), .B(G148gat), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n897), .A2(KEYINPUT59), .A3(new_n920), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n904), .B2(new_n718), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n921), .B(new_n922), .C1(G148gat), .C2(new_n924), .ZN(G1345gat));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n302), .A3(new_n716), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n897), .A2(new_n533), .A3(new_n899), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(new_n302), .ZN(G1346gat));
  AOI21_X1  g727(.A(G162gat), .B1(new_n904), .B2(new_n626), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n714), .A2(new_n303), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n900), .B2(new_n930), .ZN(G1347gat));
  NAND2_X1  g730(.A1(new_n465), .A2(new_n463), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(new_n281), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n854), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n231), .A3(new_n717), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n464), .B1(new_n850), .B2(new_n851), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n465), .A3(new_n469), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(new_n717), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n935), .B1(new_n231), .B2(new_n938), .ZN(G1348gat));
  OAI21_X1  g738(.A(new_n232), .B1(new_n937), .B2(new_n666), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT123), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n934), .A2(new_n232), .A3(new_n666), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n934), .B2(new_n533), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n716), .A2(new_n222), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n937), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n854), .A2(new_n626), .A3(new_n933), .ZN(new_n948));
  XNOR2_X1  g747(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n948), .A2(G190gat), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n948), .B2(G190gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n626), .A2(new_n223), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n950), .A2(new_n951), .B1(new_n937), .B2(new_n952), .ZN(G1351gat));
  INV_X1    g752(.A(new_n936), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(new_n903), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(new_n459), .ZN(new_n957));
  AOI21_X1  g756(.A(G197gat), .B1(new_n957), .B2(new_n698), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n282), .A2(new_n932), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n918), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n698), .A2(G197gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1352gat));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n718), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G204gat), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n459), .A2(G204gat), .A3(new_n666), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT62), .B1(new_n956), .B2(new_n965), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n956), .A2(KEYINPUT62), .A3(new_n965), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(G1353gat));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT57), .B1(new_n896), .B2(new_n343), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n852), .A2(new_n882), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n716), .B(new_n959), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  OAI21_X1  g772(.A(G211gat), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n972), .A2(new_n973), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n918), .A2(KEYINPUT126), .A3(new_n716), .A4(new_n959), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n978), .A2(new_n976), .A3(new_n969), .A4(G211gat), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n533), .A2(G211gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n955), .A2(new_n465), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n955), .A2(new_n983), .A3(new_n465), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g785(.A(KEYINPUT127), .B1(new_n977), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n976), .ZN(new_n988));
  OAI21_X1  g787(.A(KEYINPUT63), .B1(new_n988), .B2(new_n974), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n989), .A2(new_n990), .A3(new_n979), .A4(new_n985), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n987), .A2(new_n991), .ZN(G1354gat));
  NAND3_X1  g791(.A1(new_n957), .A2(new_n289), .A3(new_n626), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n960), .A2(new_n626), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n993), .B1(new_n995), .B2(new_n289), .ZN(G1355gat));
endmodule


