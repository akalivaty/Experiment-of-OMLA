

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XOR2_X1 U322 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n291) );
  XNOR2_X1 U323 ( .A(KEYINPUT4), .B(KEYINPUT93), .ZN(n290) );
  XNOR2_X1 U324 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U325 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n293) );
  XNOR2_X1 U326 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n292) );
  XNOR2_X1 U327 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U328 ( .A(n295), .B(n294), .Z(n305) );
  XOR2_X1 U329 ( .A(KEYINPUT81), .B(G134GAT), .Z(n297) );
  XNOR2_X1 U330 ( .A(KEYINPUT80), .B(G127GAT), .ZN(n296) );
  XNOR2_X1 U331 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U332 ( .A(KEYINPUT0), .B(n298), .Z(n381) );
  XOR2_X1 U333 ( .A(G155GAT), .B(KEYINPUT3), .Z(n300) );
  XNOR2_X1 U334 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n299) );
  XNOR2_X1 U335 ( .A(n300), .B(n299), .ZN(n403) );
  XOR2_X1 U336 ( .A(n403), .B(KEYINPUT1), .Z(n302) );
  NAND2_X1 U337 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U338 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U339 ( .A(n381), .B(n303), .ZN(n304) );
  XNOR2_X1 U340 ( .A(n305), .B(n304), .ZN(n313) );
  XOR2_X1 U341 ( .A(G57GAT), .B(G148GAT), .Z(n307) );
  XNOR2_X1 U342 ( .A(G141GAT), .B(G1GAT), .ZN(n306) );
  XNOR2_X1 U343 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U344 ( .A(G85GAT), .B(G120GAT), .Z(n309) );
  XNOR2_X1 U345 ( .A(G29GAT), .B(G113GAT), .ZN(n308) );
  XNOR2_X1 U346 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U347 ( .A(n311), .B(n310), .Z(n312) );
  XOR2_X1 U348 ( .A(n313), .B(n312), .Z(n481) );
  XOR2_X1 U349 ( .A(G57GAT), .B(KEYINPUT13), .Z(n363) );
  XOR2_X1 U350 ( .A(n363), .B(KEYINPUT33), .Z(n318) );
  XOR2_X1 U351 ( .A(G148GAT), .B(G106GAT), .Z(n315) );
  XNOR2_X1 U352 ( .A(G204GAT), .B(G78GAT), .ZN(n314) );
  XNOR2_X1 U353 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U354 ( .A(KEYINPUT72), .B(n316), .Z(n408) );
  XNOR2_X1 U355 ( .A(n408), .B(KEYINPUT31), .ZN(n317) );
  XNOR2_X1 U356 ( .A(n318), .B(n317), .ZN(n323) );
  XNOR2_X1 U357 ( .A(G99GAT), .B(G71GAT), .ZN(n319) );
  XNOR2_X1 U358 ( .A(n319), .B(G120GAT), .ZN(n394) );
  XOR2_X1 U359 ( .A(n394), .B(KEYINPUT32), .Z(n321) );
  NAND2_X1 U360 ( .A1(G230GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U361 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U362 ( .A(n323), .B(n322), .Z(n325) );
  XOR2_X1 U363 ( .A(G85GAT), .B(G92GAT), .Z(n344) );
  XOR2_X1 U364 ( .A(G176GAT), .B(G64GAT), .Z(n418) );
  XNOR2_X1 U365 ( .A(n344), .B(n418), .ZN(n324) );
  XNOR2_X1 U366 ( .A(n325), .B(n324), .ZN(n568) );
  XOR2_X1 U367 ( .A(G141GAT), .B(G22GAT), .Z(n400) );
  XOR2_X1 U368 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n327) );
  XNOR2_X1 U369 ( .A(G197GAT), .B(KEYINPUT70), .ZN(n326) );
  XNOR2_X1 U370 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U371 ( .A(n400), .B(n328), .Z(n330) );
  NAND2_X1 U372 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U373 ( .A(n330), .B(n329), .ZN(n332) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n331) );
  XNOR2_X1 U375 ( .A(n331), .B(G8GAT), .ZN(n367) );
  XOR2_X1 U376 ( .A(n332), .B(n367), .Z(n340) );
  XOR2_X1 U377 ( .A(G43GAT), .B(G29GAT), .Z(n334) );
  XNOR2_X1 U378 ( .A(KEYINPUT68), .B(G50GAT), .ZN(n333) );
  XNOR2_X1 U379 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U380 ( .A(n335), .B(KEYINPUT8), .Z(n337) );
  XNOR2_X1 U381 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n336) );
  XNOR2_X1 U382 ( .A(n337), .B(n336), .ZN(n358) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(G15GAT), .ZN(n338) );
  XNOR2_X1 U384 ( .A(n338), .B(G113GAT), .ZN(n382) );
  XNOR2_X1 U385 ( .A(n358), .B(n382), .ZN(n339) );
  XNOR2_X1 U386 ( .A(n340), .B(n339), .ZN(n563) );
  XOR2_X1 U387 ( .A(n563), .B(KEYINPUT71), .Z(n511) );
  INV_X1 U388 ( .A(n511), .ZN(n547) );
  NOR2_X1 U389 ( .A1(n568), .A2(n547), .ZN(n341) );
  XOR2_X1 U390 ( .A(KEYINPUT73), .B(n341), .Z(n455) );
  XOR2_X1 U391 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n343) );
  XNOR2_X1 U392 ( .A(G106GAT), .B(KEYINPUT65), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U394 ( .A(n344), .B(G162GAT), .Z(n346) );
  XNOR2_X1 U395 ( .A(G99GAT), .B(G218GAT), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U397 ( .A(n348), .B(n347), .ZN(n350) );
  AND2_X1 U398 ( .A1(G232GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U399 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U400 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n352) );
  XNOR2_X1 U401 ( .A(G134GAT), .B(KEYINPUT75), .ZN(n351) );
  XNOR2_X1 U402 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U403 ( .A(n354), .B(n353), .ZN(n360) );
  XOR2_X1 U404 ( .A(KEYINPUT67), .B(KEYINPUT76), .Z(n356) );
  XNOR2_X1 U405 ( .A(G190GAT), .B(KEYINPUT9), .ZN(n355) );
  XNOR2_X1 U406 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U407 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U408 ( .A(n360), .B(n359), .ZN(n557) );
  INV_X1 U409 ( .A(n557), .ZN(n534) );
  XOR2_X1 U410 ( .A(G155GAT), .B(G78GAT), .Z(n362) );
  XNOR2_X1 U411 ( .A(G127GAT), .B(G71GAT), .ZN(n361) );
  XNOR2_X1 U412 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U413 ( .A(n364), .B(n363), .Z(n366) );
  XNOR2_X1 U414 ( .A(G15GAT), .B(G183GAT), .ZN(n365) );
  XNOR2_X1 U415 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U416 ( .A(n367), .B(KEYINPUT12), .Z(n369) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U418 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U419 ( .A(n371), .B(n370), .Z(n379) );
  XOR2_X1 U420 ( .A(KEYINPUT79), .B(G64GAT), .Z(n373) );
  XNOR2_X1 U421 ( .A(G22GAT), .B(G211GAT), .ZN(n372) );
  XNOR2_X1 U422 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U423 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n375) );
  XNOR2_X1 U424 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n374) );
  XNOR2_X1 U425 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U426 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U427 ( .A(n379), .B(n378), .Z(n572) );
  INV_X1 U428 ( .A(n572), .ZN(n554) );
  NOR2_X1 U429 ( .A1(n534), .A2(n554), .ZN(n380) );
  XNOR2_X1 U430 ( .A(n380), .B(KEYINPUT16), .ZN(n439) );
  XOR2_X1 U431 ( .A(G176GAT), .B(KEYINPUT82), .Z(n384) );
  XNOR2_X1 U432 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U433 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U434 ( .A(G43GAT), .B(KEYINPUT20), .Z(n386) );
  NAND2_X1 U435 ( .A1(G227GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U436 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U437 ( .A(n388), .B(n387), .Z(n396) );
  XOR2_X1 U438 ( .A(G183GAT), .B(KEYINPUT83), .Z(n390) );
  XNOR2_X1 U439 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n389) );
  XNOR2_X1 U440 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U441 ( .A(n391), .B(KEYINPUT17), .Z(n393) );
  XNOR2_X1 U442 ( .A(KEYINPUT84), .B(G190GAT), .ZN(n392) );
  XNOR2_X1 U443 ( .A(n393), .B(n392), .ZN(n415) );
  XNOR2_X1 U444 ( .A(n415), .B(n394), .ZN(n395) );
  XOR2_X1 U445 ( .A(n396), .B(n395), .Z(n485) );
  XOR2_X1 U446 ( .A(n485), .B(KEYINPUT85), .Z(n428) );
  XOR2_X1 U447 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n398) );
  XNOR2_X1 U448 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n397) );
  XNOR2_X1 U449 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U450 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U451 ( .A1(G228GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U452 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U453 ( .A(n404), .B(n403), .Z(n406) );
  XNOR2_X1 U454 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n405) );
  XNOR2_X1 U455 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U456 ( .A(n408), .B(n407), .ZN(n413) );
  XOR2_X1 U457 ( .A(KEYINPUT21), .B(G218GAT), .Z(n410) );
  XNOR2_X1 U458 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n409) );
  XNOR2_X1 U459 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(n411), .ZN(n414) );
  INV_X1 U461 ( .A(n414), .ZN(n412) );
  XOR2_X1 U462 ( .A(n413), .B(n412), .Z(n543) );
  XNOR2_X1 U463 ( .A(KEYINPUT28), .B(n543), .ZN(n489) );
  INV_X1 U464 ( .A(n489), .ZN(n510) );
  XOR2_X1 U465 ( .A(n415), .B(n414), .Z(n426) );
  XOR2_X1 U466 ( .A(G204GAT), .B(G8GAT), .Z(n417) );
  XNOR2_X1 U467 ( .A(G169GAT), .B(G36GAT), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U469 ( .A(KEYINPUT94), .B(n418), .Z(n420) );
  XNOR2_X1 U470 ( .A(G92GAT), .B(KEYINPUT76), .ZN(n419) );
  XNOR2_X1 U471 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U472 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U474 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U475 ( .A(n426), .B(n425), .Z(n461) );
  XNOR2_X1 U476 ( .A(n461), .B(KEYINPUT27), .ZN(n433) );
  INV_X1 U477 ( .A(n481), .ZN(n542) );
  NAND2_X1 U478 ( .A1(n433), .A2(n542), .ZN(n507) );
  NOR2_X1 U479 ( .A1(n510), .A2(n507), .ZN(n427) );
  NAND2_X1 U480 ( .A1(n428), .A2(n427), .ZN(n438) );
  INV_X1 U481 ( .A(n485), .ZN(n545) );
  NAND2_X1 U482 ( .A1(n545), .A2(n461), .ZN(n429) );
  NAND2_X1 U483 ( .A1(n543), .A2(n429), .ZN(n430) );
  XOR2_X1 U484 ( .A(KEYINPUT25), .B(n430), .Z(n435) );
  NOR2_X1 U485 ( .A1(n545), .A2(n543), .ZN(n432) );
  XNOR2_X1 U486 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n431) );
  XOR2_X1 U487 ( .A(n432), .B(n431), .Z(n562) );
  NAND2_X1 U488 ( .A1(n433), .A2(n562), .ZN(n434) );
  NAND2_X1 U489 ( .A1(n435), .A2(n434), .ZN(n436) );
  NAND2_X1 U490 ( .A1(n481), .A2(n436), .ZN(n437) );
  NAND2_X1 U491 ( .A1(n438), .A2(n437), .ZN(n451) );
  NAND2_X1 U492 ( .A1(n439), .A2(n451), .ZN(n440) );
  XOR2_X1 U493 ( .A(KEYINPUT96), .B(n440), .Z(n469) );
  NAND2_X1 U494 ( .A1(n455), .A2(n469), .ZN(n449) );
  NOR2_X1 U495 ( .A1(n481), .A2(n449), .ZN(n441) );
  XOR2_X1 U496 ( .A(G1GAT), .B(n441), .Z(n442) );
  XNOR2_X1 U497 ( .A(KEYINPUT34), .B(n442), .ZN(G1324GAT) );
  INV_X1 U498 ( .A(n461), .ZN(n537) );
  NOR2_X1 U499 ( .A1(n537), .A2(n449), .ZN(n443) );
  XOR2_X1 U500 ( .A(G8GAT), .B(n443), .Z(G1325GAT) );
  XOR2_X1 U501 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n445) );
  XNOR2_X1 U502 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n447) );
  NOR2_X1 U504 ( .A1(n485), .A2(n449), .ZN(n446) );
  XOR2_X1 U505 ( .A(n447), .B(n446), .Z(n448) );
  XNOR2_X1 U506 ( .A(KEYINPUT97), .B(n448), .ZN(G1326GAT) );
  NOR2_X1 U507 ( .A1(n489), .A2(n449), .ZN(n450) );
  XOR2_X1 U508 ( .A(G22GAT), .B(n450), .Z(G1327GAT) );
  XOR2_X1 U509 ( .A(G29GAT), .B(KEYINPUT39), .Z(n459) );
  XNOR2_X1 U510 ( .A(n557), .B(KEYINPUT36), .ZN(n578) );
  NAND2_X1 U511 ( .A1(n554), .A2(n451), .ZN(n452) );
  NOR2_X1 U512 ( .A1(n578), .A2(n452), .ZN(n454) );
  XOR2_X1 U513 ( .A(KEYINPUT100), .B(KEYINPUT37), .Z(n453) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n479) );
  NAND2_X1 U515 ( .A1(n479), .A2(n455), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n456), .B(KEYINPUT101), .ZN(n457) );
  XNOR2_X1 U517 ( .A(KEYINPUT38), .B(n457), .ZN(n465) );
  NAND2_X1 U518 ( .A1(n465), .A2(n542), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U520 ( .A(KEYINPUT102), .B(n460), .ZN(G1328GAT) );
  NAND2_X1 U521 ( .A1(n465), .A2(n461), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U523 ( .A1(n465), .A2(n545), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT40), .ZN(n464) );
  XNOR2_X1 U525 ( .A(G43GAT), .B(n464), .ZN(G1330GAT) );
  XOR2_X1 U526 ( .A(G50GAT), .B(KEYINPUT103), .Z(n467) );
  NAND2_X1 U527 ( .A1(n465), .A2(n510), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n467), .B(n466), .ZN(G1331GAT) );
  XNOR2_X1 U529 ( .A(KEYINPUT41), .B(n568), .ZN(n550) );
  NOR2_X1 U530 ( .A1(n563), .A2(n550), .ZN(n468) );
  XOR2_X1 U531 ( .A(KEYINPUT105), .B(n468), .Z(n480) );
  NAND2_X1 U532 ( .A1(n480), .A2(n469), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n481), .A2(n476), .ZN(n472) );
  XOR2_X1 U534 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n470) );
  XNOR2_X1 U535 ( .A(G57GAT), .B(n470), .ZN(n471) );
  XNOR2_X1 U536 ( .A(n472), .B(n471), .ZN(G1332GAT) );
  NOR2_X1 U537 ( .A1(n537), .A2(n476), .ZN(n473) );
  XOR2_X1 U538 ( .A(KEYINPUT106), .B(n473), .Z(n474) );
  XNOR2_X1 U539 ( .A(G64GAT), .B(n474), .ZN(G1333GAT) );
  NOR2_X1 U540 ( .A1(n485), .A2(n476), .ZN(n475) );
  XOR2_X1 U541 ( .A(G71GAT), .B(n475), .Z(G1334GAT) );
  NOR2_X1 U542 ( .A1(n489), .A2(n476), .ZN(n478) );
  XNOR2_X1 U543 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n477) );
  XNOR2_X1 U544 ( .A(n478), .B(n477), .ZN(G1335GAT) );
  NAND2_X1 U545 ( .A1(n480), .A2(n479), .ZN(n488) );
  NOR2_X1 U546 ( .A1(n481), .A2(n488), .ZN(n482) );
  XOR2_X1 U547 ( .A(G85GAT), .B(n482), .Z(G1336GAT) );
  NOR2_X1 U548 ( .A1(n537), .A2(n488), .ZN(n484) );
  XNOR2_X1 U549 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n484), .B(n483), .ZN(G1337GAT) );
  NOR2_X1 U551 ( .A1(n485), .A2(n488), .ZN(n486) );
  XOR2_X1 U552 ( .A(KEYINPUT108), .B(n486), .Z(n487) );
  XNOR2_X1 U553 ( .A(G99GAT), .B(n487), .ZN(G1338GAT) );
  NOR2_X1 U554 ( .A1(n489), .A2(n488), .ZN(n491) );
  XNOR2_X1 U555 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U557 ( .A(G106GAT), .B(n492), .ZN(G1339GAT) );
  XNOR2_X1 U558 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n506) );
  INV_X1 U559 ( .A(n550), .ZN(n529) );
  NAND2_X1 U560 ( .A1(n563), .A2(n529), .ZN(n494) );
  XNOR2_X1 U561 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n493) );
  XNOR2_X1 U562 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U563 ( .A1(n495), .A2(n554), .ZN(n496) );
  NOR2_X1 U564 ( .A1(n534), .A2(n496), .ZN(n498) );
  XNOR2_X1 U565 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n497) );
  XNOR2_X1 U566 ( .A(n498), .B(n497), .ZN(n504) );
  NOR2_X1 U567 ( .A1(n554), .A2(n578), .ZN(n499) );
  XOR2_X1 U568 ( .A(KEYINPUT45), .B(n499), .Z(n500) );
  NOR2_X1 U569 ( .A1(n568), .A2(n500), .ZN(n501) );
  XOR2_X1 U570 ( .A(KEYINPUT112), .B(n501), .Z(n502) );
  NOR2_X1 U571 ( .A1(n511), .A2(n502), .ZN(n503) );
  NOR2_X1 U572 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n538) );
  NOR2_X1 U574 ( .A1(n538), .A2(n507), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n545), .A2(n522), .ZN(n508) );
  XOR2_X1 U576 ( .A(KEYINPUT113), .B(n508), .Z(n509) );
  NOR2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n517) );
  NAND2_X1 U578 ( .A1(n517), .A2(n511), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U580 ( .A(G120GAT), .B(KEYINPUT49), .Z(n514) );
  NAND2_X1 U581 ( .A1(n517), .A2(n529), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(G1341GAT) );
  NAND2_X1 U583 ( .A1(n572), .A2(n517), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n515), .B(KEYINPUT50), .ZN(n516) );
  XNOR2_X1 U585 ( .A(G127GAT), .B(n516), .ZN(G1342GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n519) );
  NAND2_X1 U587 ( .A1(n517), .A2(n534), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(n521) );
  XOR2_X1 U589 ( .A(G134GAT), .B(KEYINPUT114), .Z(n520) );
  XNOR2_X1 U590 ( .A(n521), .B(n520), .ZN(G1343GAT) );
  XOR2_X1 U591 ( .A(G141GAT), .B(KEYINPUT117), .Z(n525) );
  NAND2_X1 U592 ( .A1(n562), .A2(n522), .ZN(n523) );
  XOR2_X1 U593 ( .A(KEYINPUT116), .B(n523), .Z(n535) );
  NAND2_X1 U594 ( .A1(n563), .A2(n535), .ZN(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(G1344GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n527) );
  XNOR2_X1 U597 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n526) );
  XNOR2_X1 U598 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U599 ( .A(KEYINPUT118), .B(n528), .Z(n531) );
  NAND2_X1 U600 ( .A1(n529), .A2(n535), .ZN(n530) );
  XNOR2_X1 U601 ( .A(n531), .B(n530), .ZN(G1345GAT) );
  NAND2_X1 U602 ( .A1(n535), .A2(n572), .ZN(n532) );
  XNOR2_X1 U603 ( .A(n532), .B(KEYINPUT120), .ZN(n533) );
  XNOR2_X1 U604 ( .A(G155GAT), .B(n533), .ZN(G1346GAT) );
  NAND2_X1 U605 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n536), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U607 ( .A(KEYINPUT54), .ZN(n540) );
  NOR2_X1 U608 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n561) );
  NAND2_X1 U611 ( .A1(n561), .A2(n543), .ZN(n544) );
  XNOR2_X1 U612 ( .A(KEYINPUT55), .B(n544), .ZN(n546) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n556) );
  NOR2_X1 U614 ( .A1(n547), .A2(n556), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1348GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n556), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(n553), .ZN(G1349GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n556), .ZN(n555) );
  XOR2_X1 U622 ( .A(G183GAT), .B(n555), .Z(G1350GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(G190GAT), .B(n560), .Z(G1351GAT) );
  XOR2_X1 U627 ( .A(G197GAT), .B(KEYINPUT59), .Z(n565) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n577) );
  INV_X1 U629 ( .A(n577), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n573), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U635 ( .A1(n573), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(n571), .ZN(G1353GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

