//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n566,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(KEYINPUT3), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n473), .A4(new_n462), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n471), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G101), .A3(new_n473), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n468), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(G160));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n462), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT70), .Z(new_n482));
  INV_X1    g057(.A(G100), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n483), .A2(new_n473), .A3(KEYINPUT71), .ZN(new_n484));
  AOI21_X1  g059(.A(KEYINPUT71), .B1(new_n483), .B2(new_n473), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G112), .B2(new_n473), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n479), .A2(new_n473), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n482), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT72), .Z(G162));
  AND2_X1   g065(.A1(new_n473), .A2(G138), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n472), .A2(new_n462), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n473), .A3(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n465), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n472), .A2(G126), .A3(G2105), .A4(new_n462), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n473), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT73), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n496), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n501), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n503), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT75), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n511), .A2(new_n513), .B1(new_n510), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n521), .B(new_n522), .C1(new_n518), .C2(new_n517), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT76), .B(G88), .Z(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G62), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n516), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n519), .A2(new_n512), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(G651), .B1(G50), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n527), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(new_n520), .A2(new_n523), .A3(G89), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT78), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n535), .A2(KEYINPUT78), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g116(.A1(G63), .A2(G651), .ZN(new_n542));
  OR3_X1    g117(.A1(new_n516), .A2(KEYINPUT77), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(KEYINPUT77), .B1(new_n516), .B2(new_n542), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n543), .A2(new_n544), .B1(G51), .B2(new_n531), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  NAND2_X1  g122(.A1(new_n531), .A2(G52), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n525), .B2(G90), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n516), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n524), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n531), .A2(G43), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n561), .B1(new_n556), .B2(new_n557), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT80), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(new_n531), .A2(G53), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n524), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n516), .A2(KEYINPUT81), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n521), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G65), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n550), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  OR2_X1    g158(.A1(new_n521), .A2(G74), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(G49), .B2(new_n531), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n520), .A2(new_n523), .A3(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n516), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n590), .A2(KEYINPUT82), .A3(G651), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n550), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n520), .A2(new_n523), .A3(G86), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n531), .A2(G48), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n591), .A2(new_n594), .A3(new_n595), .A4(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n525), .A2(G85), .ZN(new_n598));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n516), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G47), .B2(new_n531), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT83), .B1(new_n524), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n520), .A2(new_n523), .A3(new_n607), .A4(G92), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n531), .A2(G54), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n577), .A2(G66), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n574), .B2(new_n576), .ZN(new_n618));
  INV_X1    g193(.A(new_n615), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT84), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n616), .A2(G651), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n611), .A2(new_n612), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n604), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n604), .B1(new_n624), .B2(G868), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n581), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(G868), .B2(new_n581), .ZN(G280));
  XNOR2_X1  g204(.A(KEYINPUT85), .B(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n624), .B1(G860), .B2(new_n630), .ZN(G148));
  INV_X1    g206(.A(new_n563), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n624), .A2(new_n630), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT86), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n633), .B1(new_n635), .B2(G868), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n475), .A2(new_n473), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n638), .A2(new_n465), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n480), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n487), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n473), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G2096), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n642), .A2(new_n649), .ZN(G156));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n653), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2100), .Z(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n648), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT88), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n679), .A2(new_n680), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(new_n684), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT89), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  NOR2_X1   g272(.A1(G29), .A2(G35), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G162), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT29), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G2090), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G32), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT98), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n480), .A2(G141), .ZN(new_n707));
  INV_X1    g282(.A(G105), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n638), .ZN(new_n709));
  AOI211_X1 g284(.A(new_n706), .B(new_n709), .C1(G129), .C2(new_n487), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n703), .B1(new_n710), .B2(new_n702), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT30), .B(G28), .ZN(new_n714));
  OR2_X1    g289(.A1(KEYINPUT31), .A2(G11), .ZN(new_n715));
  NAND2_X1  g290(.A1(KEYINPUT31), .A2(G11), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n714), .A2(new_n702), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n647), .B2(new_n702), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n480), .A2(G139), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n465), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n723), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n719), .B(new_n722), .C1(new_n473), .C2(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G33), .B(new_n725), .S(G29), .Z(new_n726));
  AOI21_X1  g301(.A(new_n718), .B1(new_n726), .B2(G2072), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G2072), .B2(new_n726), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G19), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n563), .B2(new_n729), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1341), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n729), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT100), .B(G1961), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR4_X1   g311(.A1(new_n713), .A2(new_n728), .A3(new_n732), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n702), .A2(G26), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT28), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n487), .A2(G128), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT95), .ZN(new_n741));
  OR2_X1    g316(.A1(G104), .A2(G2105), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n742), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n480), .A2(G140), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT94), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2067), .ZN(new_n749));
  INV_X1    g324(.A(G34), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n750), .A2(KEYINPUT24), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n702), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G160), .B2(new_n702), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT97), .ZN(new_n755));
  INV_X1    g330(.A(G2084), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n729), .A2(G20), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT23), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n581), .B2(new_n729), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n702), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n702), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2078), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n737), .A2(new_n749), .A3(new_n757), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n701), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n755), .A2(new_n756), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT101), .ZN(new_n769));
  NOR2_X1   g344(.A1(G4), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n624), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1348), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(G168), .A2(G16), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(KEYINPUT99), .C1(G16), .C2(G21), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(KEYINPUT99), .B2(new_n774), .ZN(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n767), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n729), .A2(G22), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G166), .B2(new_n729), .ZN(new_n781));
  INV_X1    g356(.A(G1971), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n729), .A2(G6), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G305), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT32), .B(G1981), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n785), .A2(new_n787), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n783), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n729), .A2(G23), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n585), .A2(new_n586), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n729), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT92), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT33), .B(G1976), .Z(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT93), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  OR3_X1    g372(.A1(new_n790), .A2(new_n797), .A3(KEYINPUT34), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT34), .B1(new_n790), .B2(new_n797), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n702), .A2(G25), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n480), .A2(G131), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n487), .A2(G119), .ZN(new_n802));
  INV_X1    g377(.A(G95), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n803), .A2(new_n473), .A3(KEYINPUT90), .ZN(new_n804));
  AOI21_X1  g379(.A(KEYINPUT90), .B1(new_n803), .B2(new_n473), .ZN(new_n805));
  OAI221_X1 g380(.A(G2104), .B1(G107), .B2(new_n473), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n801), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n800), .B1(new_n808), .B2(new_n702), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT91), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G1986), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n729), .A2(G24), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G290), .B2(G16), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n812), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n813), .B2(new_n815), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n798), .A2(new_n799), .A3(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT36), .Z(new_n819));
  NOR2_X1   g394(.A1(new_n779), .A2(new_n819), .ZN(G311));
  INV_X1    g395(.A(G311), .ZN(G150));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  INV_X1    g397(.A(G67), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n516), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n824), .A2(G651), .B1(G55), .B2(new_n531), .ZN(new_n825));
  INV_X1    g400(.A(G93), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n524), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT102), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n562), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n525), .A2(G81), .B1(new_n556), .B2(new_n557), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n825), .B(KEYINPUT102), .C1(new_n826), .C2(new_n524), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n828), .B(new_n827), .C1(new_n560), .C2(new_n562), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT38), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n624), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT103), .B(G860), .Z(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n841), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n827), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(G145));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n504), .A2(new_n505), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n747), .B(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(new_n807), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n807), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n710), .B(new_n725), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n487), .A2(G130), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n473), .A2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G142), .B2(new_n480), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(new_n640), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n853), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n852), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G160), .B(new_n647), .ZN(new_n863));
  XNOR2_X1  g438(.A(G162), .B(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n850), .A2(new_n860), .A3(new_n851), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n862), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(KEYINPUT104), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  AOI211_X1 g444(.A(new_n869), .B(new_n864), .C1(new_n862), .C2(new_n865), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n847), .B(new_n866), .C1(new_n868), .C2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g447(.A(G868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n827), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n835), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n623), .A2(G299), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n621), .A2(new_n612), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT10), .B1(new_n606), .B2(new_n608), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n882), .A3(new_n581), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n878), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n878), .B2(new_n883), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n635), .A2(new_n875), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n877), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n891));
  XOR2_X1   g466(.A(G303), .B(G305), .Z(new_n892));
  XNOR2_X1  g467(.A(G290), .B(new_n792), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n891), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n878), .B(new_n883), .C1(new_n877), .C2(new_n889), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n890), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n890), .B2(new_n902), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n899), .A2(new_n891), .A3(new_n900), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n874), .B1(new_n906), .B2(new_n873), .ZN(G295));
  OAI21_X1  g482(.A(new_n874), .B1(new_n906), .B2(new_n873), .ZN(G331));
  NOR2_X1   g483(.A1(new_n623), .A2(G299), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n581), .B1(new_n879), .B2(new_n882), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT41), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n885), .ZN(new_n912));
  NAND2_X1  g487(.A1(G286), .A2(G301), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n540), .A2(G171), .A3(new_n541), .A4(new_n545), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n913), .A2(new_n833), .A3(new_n834), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n916), .A2(new_n835), .A3(KEYINPUT107), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT107), .B1(new_n916), .B2(new_n835), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n835), .ZN(new_n921));
  AND4_X1   g496(.A1(new_n878), .A2(new_n921), .A3(new_n883), .A4(new_n915), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n894), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n847), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n887), .A2(KEYINPUT108), .B1(new_n915), .B2(new_n921), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n912), .B2(KEYINPUT108), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n916), .A2(new_n835), .A3(KEYINPUT107), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n931), .A2(new_n878), .A3(new_n883), .A4(new_n915), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n894), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n925), .A2(new_n933), .A3(KEYINPUT43), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n922), .B1(new_n912), .B2(new_n919), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n936), .B2(new_n894), .ZN(new_n937));
  INV_X1    g512(.A(new_n894), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n931), .A2(new_n915), .B1(new_n911), .B2(new_n885), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n939), .B2(new_n922), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n935), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n942), .A2(KEYINPUT44), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n925), .B2(new_n933), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT108), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n921), .A2(new_n915), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n911), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n932), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n938), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(KEYINPUT109), .A3(new_n937), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n945), .A2(new_n952), .A3(KEYINPUT43), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n937), .A2(new_n935), .A3(new_n940), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n954), .A2(KEYINPUT44), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n953), .A2(new_n955), .A3(KEYINPUT110), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT110), .B1(new_n953), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n943), .B1(new_n956), .B2(new_n957), .ZN(G397));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n504), .B2(new_n505), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n468), .A2(G40), .A3(new_n474), .A4(new_n476), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n747), .A2(G2067), .ZN(new_n965));
  INV_X1    g540(.A(G2067), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n744), .A2(new_n966), .A3(new_n746), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n710), .B(G1996), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n808), .A2(new_n811), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n808), .A2(new_n811), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(G290), .A2(G1986), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n598), .A2(new_n813), .A3(new_n602), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n964), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(G303), .A2(G8), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT55), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT45), .B(new_n959), .C1(new_n504), .C2(new_n505), .ZN(new_n980));
  INV_X1    g555(.A(new_n963), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n498), .A2(new_n502), .A3(KEYINPUT73), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n506), .B1(new_n504), .B2(new_n505), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n961), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n982), .B(KEYINPUT112), .C1(new_n985), .C2(new_n986), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n782), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n963), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n959), .B1(new_n503), .B2(new_n507), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n994), .A2(G2090), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n979), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT114), .B(G86), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n520), .A2(new_n523), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT115), .B1(new_n1002), .B2(new_n596), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n594), .A2(new_n591), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(KEYINPUT115), .A3(new_n596), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1000), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G305), .A2(G1981), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n999), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1008), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1006), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1011), .A2(new_n1004), .A3(new_n1003), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1010), .B(KEYINPUT49), .C1(new_n1012), .C2(new_n1000), .ZN(new_n1013));
  OAI21_X1  g588(.A(G8), .B1(new_n960), .B2(new_n963), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n792), .A2(G1976), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1019), .A3(new_n1015), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G288), .A2(new_n1018), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n1021), .B2(new_n1014), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT113), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1021), .A2(new_n1014), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n1019), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1016), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n981), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(new_n985), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(G2090), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n997), .B1(new_n991), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n979), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n963), .B1(new_n960), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n961), .A2(G1384), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n983), .B2(new_n984), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI211_X1 g619(.A(KEYINPUT117), .B(new_n1041), .C1(new_n983), .C2(new_n984), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n777), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1030), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n756), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G286), .A2(new_n997), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n998), .A2(new_n1029), .A3(new_n1037), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT63), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(KEYINPUT118), .A3(new_n1053), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1028), .B(KEYINPUT116), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1049), .A2(KEYINPUT63), .A3(new_n1050), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1058), .A2(KEYINPUT119), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1028), .B(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1056), .A2(new_n1057), .A3(new_n1062), .A4(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1016), .A2(new_n1018), .A3(new_n792), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1014), .B1(new_n1069), .B2(new_n1010), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1037), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1058), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1956), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n994), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n980), .A2(new_n981), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n993), .B2(new_n961), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n581), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT57), .B1(new_n573), .B2(new_n580), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1348), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1033), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n960), .A2(new_n963), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n966), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1084), .B1(new_n1089), .B2(new_n623), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1074), .A2(new_n1078), .A3(new_n1082), .A4(new_n1081), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1089), .A2(KEYINPUT60), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n1088), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1094), .A2(KEYINPUT121), .A3(new_n624), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT121), .B1(new_n1094), .B2(new_n624), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1086), .A2(new_n623), .A3(KEYINPUT60), .A4(new_n1088), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT120), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1093), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1996), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1087), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  AOI22_X1  g678(.A1(new_n1076), .A2(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n632), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1084), .A2(KEYINPUT61), .A3(new_n1091), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1092), .B1(new_n1100), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1040), .B1(new_n503), .B2(new_n507), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT117), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1039), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1118), .A2(new_n777), .B1(new_n756), .B2(new_n1047), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n997), .B1(new_n1119), .B2(G168), .ZN(new_n1120));
  AOI21_X1  g695(.A(G168), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1114), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1046), .A2(G168), .A3(new_n1048), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(new_n1114), .A3(G8), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT122), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n998), .A2(new_n1029), .A3(new_n1037), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1129));
  INV_X1    g704(.A(G2078), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(KEYINPUT53), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G1961), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1033), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(G2078), .B1(new_n989), .B2(new_n990), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1131), .B(new_n1133), .C1(new_n1134), .C2(KEYINPUT53), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G171), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n993), .A2(new_n961), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT112), .B1(new_n1137), .B2(new_n982), .ZN(new_n1138));
  INV_X1    g713(.A(new_n990), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1130), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT53), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1140), .A2(new_n1141), .B1(new_n1132), .B2(new_n1033), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1130), .A2(KEYINPUT123), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1141), .B1(KEYINPUT123), .B2(new_n1130), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n982), .A2(new_n962), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1136), .B1(new_n1146), .B2(G171), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1128), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1124), .A2(G8), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT51), .B1(new_n1150), .B2(new_n1121), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(new_n1125), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1113), .A2(new_n1127), .A3(new_n1149), .A4(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1148), .B1(new_n1146), .B2(G171), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1142), .A2(KEYINPUT124), .A3(G301), .A4(new_n1131), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1135), .B2(G171), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1155), .A2(new_n1159), .A3(KEYINPUT125), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1068), .B(new_n1072), .C1(new_n1154), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1151), .A2(new_n1152), .A3(new_n1125), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1152), .B1(new_n1151), .B2(new_n1125), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1127), .A2(KEYINPUT62), .A3(new_n1153), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1128), .A2(new_n1136), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT126), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1169), .A2(new_n1170), .A3(new_n1174), .A4(new_n1171), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n977), .B1(new_n1165), .B2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n975), .A2(new_n963), .A3(new_n962), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT48), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n973), .B2(new_n964), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n969), .A2(new_n710), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n964), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n964), .A2(new_n1101), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(KEYINPUT46), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT127), .Z(new_n1186));
  OAI211_X1 g761(.A(new_n1182), .B(new_n1186), .C1(KEYINPUT46), .C2(new_n1184), .ZN(new_n1187));
  XOR2_X1   g762(.A(new_n1187), .B(KEYINPUT47), .Z(new_n1188));
  NAND2_X1  g763(.A1(new_n969), .A2(new_n970), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n967), .B1(new_n1189), .B2(new_n971), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1180), .B(new_n1188), .C1(new_n964), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1177), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g767(.A(G227), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1194), .A2(G319), .ZN(new_n1195));
  NOR3_X1   g769(.A1(G229), .A2(G401), .A3(new_n1195), .ZN(new_n1196));
  OAI211_X1 g770(.A(new_n1196), .B(new_n871), .C1(new_n941), .C2(new_n934), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


