

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U325 ( .A(n314), .B(n313), .ZN(n318) );
  XNOR2_X1 U326 ( .A(n312), .B(n294), .ZN(n313) );
  XNOR2_X1 U327 ( .A(n340), .B(n339), .ZN(n343) );
  XOR2_X1 U328 ( .A(n326), .B(n325), .Z(n561) );
  XNOR2_X1 U329 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n447), .B(n446), .ZN(n448) );
  AND2_X1 U331 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U332 ( .A(G8GAT), .B(G183GAT), .Z(n294) );
  XOR2_X1 U333 ( .A(n424), .B(n357), .Z(n295) );
  NOR2_X1 U334 ( .A1(n578), .A2(n370), .ZN(n371) );
  XNOR2_X1 U335 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n298) );
  XNOR2_X1 U336 ( .A(n439), .B(n293), .ZN(n440) );
  XNOR2_X1 U337 ( .A(n312), .B(n298), .ZN(n301) );
  XNOR2_X1 U338 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U339 ( .A(n441), .B(n440), .ZN(n442) );
  NOR2_X1 U340 ( .A1(n568), .A2(n472), .ZN(n436) );
  XNOR2_X1 U341 ( .A(KEYINPUT37), .B(KEYINPUT106), .ZN(n479) );
  XNOR2_X1 U342 ( .A(n480), .B(n479), .ZN(n522) );
  XOR2_X1 U343 ( .A(n451), .B(n450), .Z(n528) );
  XNOR2_X1 U344 ( .A(n459), .B(G190GAT), .ZN(n460) );
  XNOR2_X1 U345 ( .A(n482), .B(G43GAT), .ZN(n483) );
  XNOR2_X1 U346 ( .A(n484), .B(n483), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n297) );
  XNOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n312) );
  XOR2_X1 U350 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XNOR2_X1 U351 ( .A(n439), .B(KEYINPUT32), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n299), .B(KEYINPUT33), .ZN(n300) );
  XOR2_X1 U353 ( .A(n301), .B(n300), .Z(n307) );
  XOR2_X1 U354 ( .A(G204GAT), .B(G64GAT), .Z(n303) );
  XNOR2_X1 U355 ( .A(G176GAT), .B(G92GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n378) );
  XNOR2_X1 U357 ( .A(G148GAT), .B(G106GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n304), .B(G78GAT), .ZN(n429) );
  XNOR2_X1 U359 ( .A(n378), .B(n429), .ZN(n305) );
  XOR2_X1 U360 ( .A(G99GAT), .B(G85GAT), .Z(n327) );
  XNOR2_X1 U361 ( .A(n305), .B(n327), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n309) );
  AND2_X1 U363 ( .A1(G230GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n575) );
  XNOR2_X1 U365 ( .A(KEYINPUT41), .B(n575), .ZN(n556) );
  XNOR2_X1 U366 ( .A(KEYINPUT108), .B(n556), .ZN(n541) );
  XOR2_X1 U367 ( .A(G22GAT), .B(G155GAT), .Z(n424) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(KEYINPUT70), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n310), .B(G15GAT), .ZN(n357) );
  NAND2_X1 U370 ( .A1(G231GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n295), .B(n311), .ZN(n314) );
  XOR2_X1 U372 ( .A(G78GAT), .B(KEYINPUT82), .Z(n316) );
  XNOR2_X1 U373 ( .A(G127GAT), .B(KEYINPUT14), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U375 ( .A(n318), .B(n317), .Z(n326) );
  XOR2_X1 U376 ( .A(G211GAT), .B(KEYINPUT15), .Z(n320) );
  XNOR2_X1 U377 ( .A(KEYINPUT12), .B(KEYINPUT80), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U379 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n322) );
  XNOR2_X1 U380 ( .A(G71GAT), .B(G64GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U383 ( .A(G134GAT), .B(KEYINPUT78), .Z(n396) );
  XOR2_X1 U384 ( .A(G36GAT), .B(G190GAT), .Z(n382) );
  XOR2_X1 U385 ( .A(n327), .B(n382), .Z(n329) );
  NAND2_X1 U386 ( .A1(G232GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n396), .B(n330), .ZN(n340) );
  XOR2_X1 U389 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n332) );
  XNOR2_X1 U390 ( .A(G218GAT), .B(KEYINPUT75), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U392 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n334) );
  XNOR2_X1 U393 ( .A(KEYINPUT79), .B(KEYINPUT76), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U395 ( .A(n336), .B(n335), .Z(n338) );
  INV_X1 U396 ( .A(G92GAT), .ZN(n337) );
  XNOR2_X1 U397 ( .A(G50GAT), .B(G162GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n341), .B(KEYINPUT74), .ZN(n418) );
  XNOR2_X1 U399 ( .A(n418), .B(G106GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U401 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n345) );
  XNOR2_X1 U402 ( .A(G43GAT), .B(G29GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U404 ( .A(KEYINPUT7), .B(n346), .ZN(n365) );
  INV_X1 U405 ( .A(n365), .ZN(n347) );
  XOR2_X2 U406 ( .A(n348), .B(n347), .Z(n564) );
  XNOR2_X1 U407 ( .A(n564), .B(KEYINPUT36), .ZN(n584) );
  NOR2_X1 U408 ( .A1(n561), .A2(n584), .ZN(n349) );
  XOR2_X1 U409 ( .A(KEYINPUT45), .B(n349), .Z(n350) );
  NOR2_X1 U410 ( .A1(n350), .A2(n575), .ZN(n351) );
  XNOR2_X1 U411 ( .A(KEYINPUT114), .B(n351), .ZN(n368) );
  XOR2_X1 U412 ( .A(KEYINPUT67), .B(G22GAT), .Z(n353) );
  XNOR2_X1 U413 ( .A(G113GAT), .B(G141GAT), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U415 ( .A(n354), .B(G36GAT), .Z(n356) );
  XOR2_X1 U416 ( .A(G169GAT), .B(G8GAT), .Z(n385) );
  XNOR2_X1 U417 ( .A(n385), .B(G50GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n361) );
  XOR2_X1 U419 ( .A(n357), .B(KEYINPUT66), .Z(n359) );
  NAND2_X1 U420 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U422 ( .A(n361), .B(n360), .Z(n367) );
  XOR2_X1 U423 ( .A(KEYINPUT30), .B(G197GAT), .Z(n363) );
  XNOR2_X1 U424 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U426 ( .A(n365), .B(n364), .Z(n366) );
  XOR2_X1 U427 ( .A(n367), .B(n366), .Z(n511) );
  INV_X1 U428 ( .A(n511), .ZN(n571) );
  NAND2_X1 U429 ( .A1(n368), .A2(n571), .ZN(n376) );
  INV_X1 U430 ( .A(n561), .ZN(n578) );
  NOR2_X1 U431 ( .A1(n571), .A2(n556), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n369), .B(KEYINPUT46), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(KEYINPUT112), .ZN(n372) );
  NAND2_X1 U434 ( .A1(n372), .A2(n564), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n373), .B(KEYINPUT113), .ZN(n374) );
  XNOR2_X1 U436 ( .A(KEYINPUT47), .B(n374), .ZN(n375) );
  NAND2_X1 U437 ( .A1(n376), .A2(n375), .ZN(n377) );
  XOR2_X1 U438 ( .A(n377), .B(KEYINPUT48), .Z(n535) );
  XOR2_X1 U439 ( .A(KEYINPUT95), .B(n378), .Z(n380) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U442 ( .A(n382), .B(n381), .Z(n387) );
  XOR2_X1 U443 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n384) );
  XNOR2_X1 U444 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n443) );
  XNOR2_X1 U446 ( .A(n385), .B(n443), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U448 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n389) );
  XNOR2_X1 U449 ( .A(G218GAT), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U451 ( .A(G197GAT), .B(n390), .Z(n427) );
  XOR2_X1 U452 ( .A(n391), .B(n427), .Z(n526) );
  INV_X1 U453 ( .A(n526), .ZN(n495) );
  XOR2_X1 U454 ( .A(n495), .B(KEYINPUT122), .Z(n392) );
  NOR2_X1 U455 ( .A1(n535), .A2(n392), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n393), .B(KEYINPUT54), .ZN(n416) );
  XOR2_X1 U457 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n395) );
  XNOR2_X1 U458 ( .A(G141GAT), .B(KEYINPUT92), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n430) );
  XOR2_X1 U460 ( .A(n430), .B(G85GAT), .Z(n398) );
  XNOR2_X1 U461 ( .A(G162GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n398), .B(n397), .ZN(n411) );
  XOR2_X1 U463 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n400) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(KEYINPUT6), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U466 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n402) );
  XNOR2_X1 U467 ( .A(G1GAT), .B(G120GAT), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U469 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U470 ( .A(G57GAT), .B(G148GAT), .Z(n406) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U472 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U473 ( .A(G155GAT), .B(n407), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U476 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n413) );
  XNOR2_X1 U477 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n412) );
  XNOR2_X1 U478 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U479 ( .A(G113GAT), .B(n414), .ZN(n450) );
  XOR2_X1 U480 ( .A(n415), .B(n450), .Z(n491) );
  INV_X1 U481 ( .A(n491), .ZN(n524) );
  NAND2_X1 U482 ( .A1(n416), .A2(n524), .ZN(n417) );
  XNOR2_X1 U483 ( .A(n417), .B(KEYINPUT64), .ZN(n568) );
  XOR2_X1 U484 ( .A(n418), .B(KEYINPUT90), .Z(n420) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U486 ( .A(n420), .B(n419), .ZN(n434) );
  XOR2_X1 U487 ( .A(KEYINPUT89), .B(KEYINPUT93), .Z(n422) );
  XNOR2_X1 U488 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U490 ( .A(n423), .B(KEYINPUT22), .Z(n426) );
  XNOR2_X1 U491 ( .A(n424), .B(G204GAT), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U493 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U496 ( .A(n434), .B(n433), .Z(n472) );
  XNOR2_X1 U497 ( .A(KEYINPUT55), .B(KEYINPUT123), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n452) );
  XOR2_X1 U499 ( .A(G190GAT), .B(G99GAT), .Z(n438) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G134GAT), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n441) );
  XOR2_X1 U502 ( .A(n442), .B(KEYINPUT20), .Z(n449) );
  XNOR2_X1 U503 ( .A(n443), .B(KEYINPUT88), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT87), .B(G176GAT), .Z(n445) );
  XNOR2_X1 U505 ( .A(G169GAT), .B(G15GAT), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U507 ( .A(n528), .ZN(n536) );
  NAND2_X1 U508 ( .A1(n452), .A2(n536), .ZN(n566) );
  NOR2_X1 U509 ( .A1(n541), .A2(n566), .ZN(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n453) );
  XNOR2_X1 U511 ( .A(n453), .B(G176GAT), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  NOR2_X1 U513 ( .A1(n561), .A2(n566), .ZN(n458) );
  INV_X1 U514 ( .A(G183GAT), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n456), .B(KEYINPUT124), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(G1350GAT) );
  NOR2_X1 U517 ( .A1(n564), .A2(n566), .ZN(n461) );
  INV_X1 U518 ( .A(KEYINPUT58), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XNOR2_X1 U520 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n464) );
  NOR2_X1 U521 ( .A1(n528), .A2(n526), .ZN(n462) );
  NOR2_X1 U522 ( .A1(n472), .A2(n462), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n495), .B(KEYINPUT27), .ZN(n471) );
  NAND2_X1 U525 ( .A1(n472), .A2(n528), .ZN(n465) );
  XOR2_X1 U526 ( .A(n465), .B(KEYINPUT26), .Z(n569) );
  NAND2_X1 U527 ( .A1(n471), .A2(n569), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U529 ( .A(KEYINPUT97), .B(n468), .Z(n469) );
  NAND2_X1 U530 ( .A1(n469), .A2(n524), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(KEYINPUT98), .ZN(n476) );
  NAND2_X1 U532 ( .A1(n491), .A2(n471), .ZN(n534) );
  NOR2_X1 U533 ( .A1(n536), .A2(n534), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n472), .B(KEYINPUT28), .ZN(n473) );
  XOR2_X1 U535 ( .A(n473), .B(KEYINPUT65), .Z(n501) );
  INV_X1 U536 ( .A(n501), .ZN(n538) );
  NAND2_X1 U537 ( .A1(n474), .A2(n538), .ZN(n475) );
  NAND2_X1 U538 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U539 ( .A(KEYINPUT99), .B(n477), .ZN(n488) );
  NOR2_X1 U540 ( .A1(n488), .A2(n584), .ZN(n478) );
  NAND2_X1 U541 ( .A1(n561), .A2(n478), .ZN(n480) );
  NOR2_X1 U542 ( .A1(n571), .A2(n575), .ZN(n489) );
  NAND2_X1 U543 ( .A1(n522), .A2(n489), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n481), .B(KEYINPUT38), .ZN(n509) );
  NOR2_X1 U545 ( .A1(n528), .A2(n509), .ZN(n484) );
  XNOR2_X1 U546 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n482) );
  XOR2_X1 U547 ( .A(KEYINPUT101), .B(KEYINPUT34), .Z(n493) );
  NAND2_X1 U548 ( .A1(n578), .A2(n564), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n485), .B(KEYINPUT16), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n486), .B(KEYINPUT84), .ZN(n487) );
  NOR2_X1 U551 ( .A1(n488), .A2(n487), .ZN(n512) );
  NAND2_X1 U552 ( .A1(n512), .A2(n489), .ZN(n490) );
  XOR2_X1 U553 ( .A(KEYINPUT100), .B(n490), .Z(n502) );
  NAND2_X1 U554 ( .A1(n491), .A2(n502), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NAND2_X1 U557 ( .A1(n502), .A2(n495), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n498) );
  NAND2_X1 U560 ( .A1(n502), .A2(n536), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n500) );
  XOR2_X1 U562 ( .A(G15GAT), .B(KEYINPUT102), .Z(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n504) );
  NAND2_X1 U565 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G22GAT), .B(n505), .ZN(G1327GAT) );
  NOR2_X1 U568 ( .A1(n509), .A2(n524), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(KEYINPUT39), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G29GAT), .B(n507), .ZN(G1328GAT) );
  NOR2_X1 U571 ( .A1(n526), .A2(n509), .ZN(n508) );
  XOR2_X1 U572 ( .A(G36GAT), .B(n508), .Z(G1329GAT) );
  NOR2_X1 U573 ( .A1(n538), .A2(n509), .ZN(n510) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n510), .Z(G1331GAT) );
  NOR2_X1 U575 ( .A1(n541), .A2(n511), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n512), .A2(n523), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n524), .A2(n518), .ZN(n513) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n513), .Z(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n526), .A2(n518), .ZN(n515) );
  XOR2_X1 U581 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U582 ( .A1(n528), .A2(n518), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  NOR2_X1 U585 ( .A1(n538), .A2(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(n521), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n531) );
  NOR2_X1 U590 ( .A1(n524), .A2(n531), .ZN(n525) );
  XOR2_X1 U591 ( .A(G85GAT), .B(n525), .Z(G1336GAT) );
  NOR2_X1 U592 ( .A1(n526), .A2(n531), .ZN(n527) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n527), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n531), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(G1338GAT) );
  NOR2_X1 U597 ( .A1(n538), .A2(n531), .ZN(n532) );
  XOR2_X1 U598 ( .A(KEYINPUT44), .B(n532), .Z(n533) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n553) );
  NAND2_X1 U601 ( .A1(n553), .A2(n536), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT115), .B(n537), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n549) );
  NOR2_X1 U604 ( .A1(n571), .A2(n549), .ZN(n540) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n540), .Z(G1340GAT) );
  NOR2_X1 U606 ( .A1(n549), .A2(n541), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n543) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT116), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U611 ( .A1(n561), .A2(n549), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U614 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  NOR2_X1 U615 ( .A1(n564), .A2(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  NAND2_X1 U619 ( .A1(n553), .A2(n569), .ZN(n563) );
  NOR2_X1 U620 ( .A1(n571), .A2(n563), .ZN(n554) );
  XOR2_X1 U621 ( .A(G141GAT), .B(n554), .Z(n555) );
  XNOR2_X1 U622 ( .A(KEYINPUT120), .B(n555), .ZN(G1344GAT) );
  NOR2_X1 U623 ( .A1(n563), .A2(n556), .ZN(n560) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n558) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n563), .ZN(n562) );
  XOR2_X1 U629 ( .A(G155GAT), .B(n562), .Z(G1346GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NOR2_X1 U632 ( .A1(n571), .A2(n566), .ZN(n567) );
  XOR2_X1 U633 ( .A(G169GAT), .B(n567), .Z(G1348GAT) );
  INV_X1 U634 ( .A(n568), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n583) );
  NOR2_X1 U636 ( .A1(n571), .A2(n583), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U641 ( .A(n583), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT125), .Z(n582) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(n586), .B(n585), .Z(G1355GAT) );
endmodule

