

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772;

  XNOR2_X1 U367 ( .A(n387), .B(KEYINPUT79), .ZN(n352) );
  NOR2_X1 U368 ( .A1(G953), .A2(G237), .ZN(n575) );
  XOR2_X1 U369 ( .A(KEYINPUT18), .B(KEYINPUT81), .Z(n344) );
  NAND2_X2 U370 ( .A1(n487), .A2(n489), .ZN(n488) );
  NOR2_X2 U371 ( .A1(n660), .A2(n772), .ZN(n644) );
  XNOR2_X2 U372 ( .A(n518), .B(G101), .ZN(n522) );
  NOR2_X1 U373 ( .A1(n652), .A2(G902), .ZN(n527) );
  XNOR2_X2 U374 ( .A(n536), .B(n537), .ZN(n756) );
  XNOR2_X2 U375 ( .A(n558), .B(G140), .ZN(n536) );
  NAND2_X1 U376 ( .A1(n355), .A2(n353), .ZN(n681) );
  AND2_X1 U377 ( .A1(n358), .A2(n356), .ZN(n355) );
  NAND2_X1 U378 ( .A1(n354), .A2(KEYINPUT48), .ZN(n353) );
  XNOR2_X1 U379 ( .A(n382), .B(n431), .ZN(n360) );
  INV_X1 U380 ( .A(n611), .ZN(n597) );
  OR2_X2 U381 ( .A1(n345), .A2(n560), .ZN(n452) );
  NOR2_X2 U382 ( .A1(n724), .A2(G902), .ZN(n535) );
  INV_X1 U383 ( .A(G146), .ZN(n507) );
  INV_X1 U384 ( .A(KEYINPUT64), .ZN(n493) );
  INV_X4 U385 ( .A(G953), .ZN(n763) );
  NOR2_X1 U386 ( .A1(n722), .A2(G953), .ZN(n723) );
  NAND2_X1 U387 ( .A1(n360), .A2(n357), .ZN(n356) );
  INV_X1 U388 ( .A(n360), .ZN(n354) );
  NOR2_X1 U389 ( .A1(n359), .A2(n371), .ZN(n358) );
  AND2_X1 U390 ( .A1(n393), .A2(n392), .ZN(n391) );
  AND2_X1 U391 ( .A1(n367), .A2(n417), .ZN(n357) );
  NAND2_X1 U392 ( .A1(n408), .A2(n406), .ZN(n769) );
  NAND2_X1 U393 ( .A1(n500), .A2(n678), .ZN(n371) );
  AND2_X1 U394 ( .A1(n409), .A2(n411), .ZN(n408) );
  NAND2_X1 U395 ( .A1(n423), .A2(n422), .ZN(n425) );
  NAND2_X1 U396 ( .A1(n418), .A2(n424), .ZN(n422) );
  AND2_X1 U397 ( .A1(n420), .A2(n419), .ZN(n423) );
  NOR2_X1 U398 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U399 ( .A1(n625), .A2(n432), .ZN(n656) );
  AND2_X1 U400 ( .A1(n472), .A2(n471), .ZN(n697) );
  XNOR2_X1 U401 ( .A(n624), .B(n473), .ZN(n472) );
  NOR2_X1 U402 ( .A1(n638), .A2(n685), .ZN(n639) );
  XNOR2_X1 U403 ( .A(n348), .B(n551), .ZN(n692) );
  NOR2_X1 U404 ( .A1(n591), .A2(n401), .ZN(n405) );
  NAND2_X1 U405 ( .A1(n351), .A2(n349), .ZN(n348) );
  NAND2_X1 U406 ( .A1(n597), .A2(n400), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n688), .B(KEYINPUT104), .ZN(n591) );
  NAND2_X1 U408 ( .A1(n466), .A2(n350), .ZN(n349) );
  XOR2_X1 U409 ( .A(n733), .B(n732), .Z(n509) );
  XNOR2_X1 U410 ( .A(n582), .B(n479), .ZN(n586) );
  NAND2_X1 U411 ( .A1(n467), .A2(n469), .ZN(n465) );
  XNOR2_X1 U412 ( .A(n412), .B(n533), .ZN(n724) );
  XNOR2_X1 U413 ( .A(n494), .B(n752), .ZN(n345) );
  XNOR2_X1 U414 ( .A(n546), .B(n545), .ZN(n741) );
  XNOR2_X1 U415 ( .A(n756), .B(n540), .ZN(n546) );
  XNOR2_X1 U416 ( .A(n365), .B(KEYINPUT91), .ZN(n449) );
  XNOR2_X1 U417 ( .A(n389), .B(n559), .ZN(n497) );
  XNOR2_X1 U418 ( .A(n363), .B(n508), .ZN(n567) );
  XNOR2_X1 U419 ( .A(n520), .B(n519), .ZN(n521) );
  INV_X2 U420 ( .A(G128), .ZN(n347) );
  INV_X2 U421 ( .A(G125), .ZN(n361) );
  XOR2_X1 U422 ( .A(G122), .B(KEYINPUT16), .Z(n559) );
  XOR2_X1 U423 ( .A(G902), .B(KEYINPUT15), .Z(n560) );
  XOR2_X1 U424 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n544) );
  XNOR2_X1 U425 ( .A(n345), .B(KEYINPUT55), .ZN(n647) );
  INV_X1 U426 ( .A(n346), .ZN(n398) );
  NAND2_X1 U427 ( .A1(n372), .A2(n346), .ZN(n618) );
  XNOR2_X2 U428 ( .A(n347), .B(G143), .ZN(n363) );
  AND2_X1 U429 ( .A1(n686), .A2(n364), .ZN(n350) );
  NAND2_X1 U430 ( .A1(n465), .A2(n686), .ZN(n351) );
  NAND2_X1 U431 ( .A1(n352), .A2(n701), .ZN(n428) );
  NAND2_X1 U432 ( .A1(n352), .A2(n632), .ZN(n583) );
  NOR2_X1 U433 ( .A1(n367), .A2(n417), .ZN(n359) );
  XNOR2_X2 U434 ( .A(n361), .B(G146), .ZN(n558) );
  NAND2_X1 U435 ( .A1(n697), .A2(n628), .ZN(n416) );
  NAND2_X1 U436 ( .A1(n636), .A2(n627), .ZN(n641) );
  INV_X1 U437 ( .A(n623), .ZN(n362) );
  XNOR2_X1 U438 ( .A(n596), .B(KEYINPUT1), .ZN(n691) );
  AND2_X1 U439 ( .A1(n378), .A2(n645), .ZN(n388) );
  NOR2_X1 U440 ( .A1(n681), .A2(n646), .ZN(n485) );
  NAND2_X1 U441 ( .A1(n549), .A2(G221), .ZN(n550) );
  INV_X1 U442 ( .A(KEYINPUT76), .ZN(n473) );
  INV_X1 U443 ( .A(n677), .ZN(n500) );
  INV_X1 U444 ( .A(KEYINPUT45), .ZN(n474) );
  NAND2_X1 U445 ( .A1(n478), .A2(n477), .ZN(n602) );
  INV_X1 U446 ( .A(n586), .ZN(n478) );
  XNOR2_X1 U447 ( .A(n621), .B(n622), .ZN(n636) );
  XOR2_X1 U448 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n577) );
  XOR2_X1 U449 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n574) );
  XOR2_X1 U450 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n542) );
  INV_X1 U451 ( .A(n454), .ZN(n471) );
  NOR2_X1 U452 ( .A1(G902), .A2(G237), .ZN(n528) );
  INV_X1 U453 ( .A(n589), .ZN(n499) );
  INV_X1 U454 ( .A(KEYINPUT69), .ZN(n551) );
  XNOR2_X1 U455 ( .A(n524), .B(n525), .ZN(n506) );
  INV_X1 U456 ( .A(G134), .ZN(n508) );
  XNOR2_X1 U457 ( .A(n379), .B(n563), .ZN(n565) );
  XNOR2_X1 U458 ( .A(n562), .B(n380), .ZN(n379) );
  INV_X1 U459 ( .A(KEYINPUT98), .ZN(n380) );
  XNOR2_X1 U460 ( .A(G116), .B(G107), .ZN(n564) );
  XNOR2_X1 U461 ( .A(n496), .B(n495), .ZN(n494) );
  XNOR2_X1 U462 ( .A(n557), .B(n556), .ZN(n496) );
  NOR2_X1 U463 ( .A1(KEYINPUT85), .A2(n679), .ZN(n680) );
  INV_X1 U464 ( .A(KEYINPUT39), .ZN(n462) );
  XNOR2_X1 U465 ( .A(n608), .B(n381), .ZN(n458) );
  INV_X1 U466 ( .A(KEYINPUT110), .ZN(n381) );
  XNOR2_X1 U467 ( .A(n581), .B(G475), .ZN(n479) );
  NOR2_X1 U468 ( .A1(G902), .A2(n731), .ZN(n582) );
  XNOR2_X1 U469 ( .A(n570), .B(G478), .ZN(n477) );
  AND2_X1 U470 ( .A1(n692), .A2(n596), .ZN(n552) );
  NOR2_X2 U471 ( .A1(n399), .A2(n398), .ZN(n619) );
  BUF_X1 U472 ( .A(n688), .Z(n454) );
  NAND2_X1 U473 ( .A1(n464), .A2(n463), .ZN(n685) );
  NOR2_X1 U474 ( .A1(G952), .A2(n763), .ZN(n745) );
  INV_X1 U475 ( .A(KEYINPUT46), .ZN(n431) );
  XNOR2_X1 U476 ( .A(n607), .B(KEYINPUT47), .ZN(n429) );
  XNOR2_X1 U477 ( .A(n434), .B(n433), .ZN(n549) );
  INV_X1 U478 ( .A(KEYINPUT20), .ZN(n433) );
  NOR2_X1 U479 ( .A1(n560), .A2(n435), .ZN(n434) );
  INV_X1 U480 ( .A(G234), .ZN(n435) );
  INV_X1 U481 ( .A(KEYINPUT68), .ZN(n383) );
  AND2_X1 U482 ( .A1(n644), .A2(n385), .ZN(n384) );
  INV_X1 U483 ( .A(KEYINPUT44), .ZN(n385) );
  INV_X1 U484 ( .A(KEYINPUT48), .ZN(n417) );
  XNOR2_X1 U485 ( .A(n567), .B(n517), .ZN(n757) );
  XNOR2_X1 U486 ( .A(G104), .B(G122), .ZN(n573) );
  XNOR2_X1 U487 ( .A(n530), .B(G101), .ZN(n427) );
  INV_X1 U488 ( .A(KEYINPUT80), .ZN(n529) );
  XNOR2_X1 U489 ( .A(n757), .B(n507), .ZN(n412) );
  NAND2_X1 U490 ( .A1(n560), .A2(KEYINPUT2), .ZN(n483) );
  XNOR2_X1 U491 ( .A(n555), .B(n554), .ZN(n556) );
  INV_X1 U492 ( .A(KEYINPUT90), .ZN(n554) );
  NAND2_X1 U493 ( .A1(n763), .A2(G224), .ZN(n555) );
  NAND2_X1 U494 ( .A1(G234), .A2(G237), .ZN(n511) );
  AND2_X1 U495 ( .A1(n620), .A2(n686), .ZN(n451) );
  INV_X1 U496 ( .A(G902), .ZN(n468) );
  XNOR2_X1 U497 ( .A(G128), .B(G137), .ZN(n538) );
  INV_X1 U498 ( .A(KEYINPUT31), .ZN(n415) );
  NAND2_X1 U499 ( .A1(n404), .A2(n498), .ZN(n387) );
  XNOR2_X1 U500 ( .A(n405), .B(n376), .ZN(n404) );
  AND2_X1 U501 ( .A1(n552), .A2(n499), .ZN(n498) );
  NOR2_X1 U502 ( .A1(n401), .A2(n604), .ZN(n400) );
  XNOR2_X1 U503 ( .A(n460), .B(n569), .ZN(n459) );
  XOR2_X1 U504 ( .A(n648), .B(n647), .Z(n510) );
  XNOR2_X1 U505 ( .A(n455), .B(KEYINPUT86), .ZN(n721) );
  NAND2_X1 U506 ( .A1(n407), .A2(n410), .ZN(n406) );
  NOR2_X1 U507 ( .A1(n601), .A2(n638), .ZN(n675) );
  XNOR2_X1 U508 ( .A(n457), .B(KEYINPUT36), .ZN(n601) );
  NAND2_X1 U509 ( .A1(n458), .A2(n370), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n602), .B(n476), .ZN(n666) );
  INV_X1 U511 ( .A(KEYINPUT105), .ZN(n476) );
  INV_X1 U512 ( .A(n477), .ZN(n584) );
  NAND2_X1 U513 ( .A1(n397), .A2(n369), .ZN(n448) );
  NAND2_X1 U514 ( .A1(n503), .A2(n502), .ZN(n501) );
  INV_X1 U515 ( .A(n745), .ZN(n502) );
  XNOR2_X1 U516 ( .A(n504), .B(n377), .ZN(n503) );
  AND2_X1 U517 ( .A1(n548), .A2(n468), .ZN(n364) );
  AND2_X1 U518 ( .A1(G210), .A2(n561), .ZN(n365) );
  OR2_X1 U519 ( .A1(n617), .A2(n616), .ZN(n366) );
  INV_X1 U520 ( .A(n706), .ZN(n626) );
  INV_X1 U521 ( .A(n700), .ZN(n401) );
  AND2_X1 U522 ( .A1(n430), .A2(n429), .ZN(n367) );
  OR2_X1 U523 ( .A1(n700), .A2(n402), .ZN(n368) );
  INV_X1 U524 ( .A(n548), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n547), .B(KEYINPUT25), .ZN(n548) );
  AND2_X1 U526 ( .A1(n623), .A2(n685), .ZN(n369) );
  AND2_X1 U527 ( .A1(n597), .A2(n700), .ZN(n370) );
  AND2_X1 U528 ( .A1(n403), .A2(n368), .ZN(n372) );
  AND2_X1 U529 ( .A1(n368), .A2(n366), .ZN(n373) );
  XOR2_X1 U530 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n374) );
  XOR2_X1 U531 ( .A(KEYINPUT88), .B(KEYINPUT33), .Z(n375) );
  XNOR2_X1 U532 ( .A(KEYINPUT30), .B(KEYINPUT106), .ZN(n376) );
  XOR2_X1 U533 ( .A(n652), .B(KEYINPUT62), .Z(n377) );
  INV_X1 U534 ( .A(KEYINPUT101), .ZN(n446) );
  BUF_X1 U535 ( .A(n730), .Z(n740) );
  XOR2_X1 U536 ( .A(n363), .B(n558), .Z(n495) );
  INV_X1 U537 ( .A(n641), .ZN(n397) );
  INV_X1 U538 ( .A(n567), .ZN(n460) );
  XNOR2_X1 U539 ( .A(n767), .B(n383), .ZN(n386) );
  NAND2_X1 U540 ( .A1(n386), .A2(n384), .ZN(n378) );
  NAND2_X1 U541 ( .A1(n391), .A2(n394), .ZN(n390) );
  XNOR2_X1 U542 ( .A(n566), .B(n459), .ZN(n736) );
  NAND2_X1 U543 ( .A1(n390), .A2(n633), .ZN(n414) );
  NAND2_X1 U544 ( .A1(n706), .A2(KEYINPUT101), .ZN(n443) );
  XNOR2_X1 U545 ( .A(n414), .B(KEYINPUT87), .ZN(n475) );
  NAND2_X1 U546 ( .A1(n769), .A2(n771), .ZN(n382) );
  NAND2_X1 U547 ( .A1(n388), .A2(n475), .ZN(n450) );
  NAND2_X1 U548 ( .A1(n438), .A2(n437), .ZN(n447) );
  XNOR2_X1 U549 ( .A(n427), .B(n389), .ZN(n532) );
  XNOR2_X2 U550 ( .A(n426), .B(G107), .ZN(n389) );
  NAND2_X1 U551 ( .A1(n439), .A2(n413), .ZN(n392) );
  NAND2_X1 U552 ( .A1(n442), .A2(n413), .ZN(n393) );
  NAND2_X1 U553 ( .A1(n396), .A2(n395), .ZN(n394) );
  INV_X1 U554 ( .A(n442), .ZN(n395) );
  NOR2_X1 U555 ( .A1(n439), .A2(n413), .ZN(n396) );
  INV_X1 U556 ( .A(n448), .ZN(n653) );
  NAND2_X1 U557 ( .A1(n403), .A2(n373), .ZN(n399) );
  INV_X1 U558 ( .A(n604), .ZN(n402) );
  NAND2_X1 U559 ( .A1(n611), .A2(n604), .ZN(n403) );
  INV_X1 U560 ( .A(n585), .ZN(n407) );
  NAND2_X1 U561 ( .A1(n585), .A2(n374), .ZN(n409) );
  XNOR2_X2 U562 ( .A(n428), .B(n462), .ZN(n585) );
  NOR2_X1 U563 ( .A1(n602), .A2(n374), .ZN(n410) );
  NAND2_X1 U564 ( .A1(n602), .A2(n374), .ZN(n411) );
  XNOR2_X1 U565 ( .A(n412), .B(n505), .ZN(n652) );
  INV_X1 U566 ( .A(KEYINPUT102), .ZN(n413) );
  INV_X1 U567 ( .A(n438), .ZN(n668) );
  XNOR2_X2 U568 ( .A(n416), .B(n415), .ZN(n438) );
  AND2_X1 U569 ( .A1(n421), .A2(n632), .ZN(n419) );
  NAND2_X1 U570 ( .A1(n445), .A2(KEYINPUT101), .ZN(n444) );
  XOR2_X2 U571 ( .A(G131), .B(KEYINPUT71), .Z(n571) );
  INV_X1 U572 ( .A(n716), .ZN(n418) );
  NAND2_X1 U573 ( .A1(n716), .A2(n631), .ZN(n420) );
  NAND2_X1 U574 ( .A1(n629), .A2(n631), .ZN(n421) );
  NOR2_X1 U575 ( .A1(n629), .A2(n631), .ZN(n424) );
  XNOR2_X2 U576 ( .A(n425), .B(KEYINPUT35), .ZN(n767) );
  XNOR2_X2 U577 ( .A(G104), .B(G110), .ZN(n426) );
  NOR2_X1 U578 ( .A1(n664), .A2(n675), .ZN(n430) );
  INV_X1 U579 ( .A(n552), .ZN(n432) );
  INV_X1 U580 ( .A(n560), .ZN(n646) );
  XNOR2_X2 U581 ( .A(n497), .B(n436), .ZN(n752) );
  XNOR2_X1 U582 ( .A(n506), .B(n436), .ZN(n505) );
  XNOR2_X2 U583 ( .A(n521), .B(n522), .ZN(n436) );
  INV_X1 U584 ( .A(n656), .ZN(n437) );
  NAND2_X1 U585 ( .A1(n448), .A2(n440), .ZN(n439) );
  NAND2_X1 U586 ( .A1(n447), .A2(n441), .ZN(n440) );
  AND2_X1 U587 ( .A1(n626), .A2(n446), .ZN(n441) );
  NAND2_X1 U588 ( .A1(n444), .A2(n443), .ZN(n442) );
  INV_X1 U589 ( .A(n447), .ZN(n445) );
  XNOR2_X2 U590 ( .A(n452), .B(n449), .ZN(n611) );
  XNOR2_X2 U591 ( .A(n450), .B(n474), .ZN(n746) );
  NAND2_X1 U592 ( .A1(n730), .A2(G475), .ZN(n734) );
  XNOR2_X2 U593 ( .A(n488), .B(n493), .ZN(n730) );
  NAND2_X1 U594 ( .A1(n730), .A2(G210), .ZN(n649) );
  NAND2_X1 U595 ( .A1(n628), .A2(n451), .ZN(n621) );
  XNOR2_X2 U596 ( .A(n619), .B(KEYINPUT0), .ZN(n628) );
  XNOR2_X2 U597 ( .A(n453), .B(n375), .ZN(n716) );
  NAND2_X1 U598 ( .A1(n472), .A2(n599), .ZN(n453) );
  XNOR2_X2 U599 ( .A(G113), .B(KEYINPUT72), .ZN(n518) );
  NAND2_X1 U600 ( .A1(n684), .A2(n683), .ZN(n455) );
  XNOR2_X1 U601 ( .A(n456), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U602 ( .A1(n735), .A2(n745), .ZN(n456) );
  INV_X1 U603 ( .A(n746), .ZN(n486) );
  XNOR2_X1 U604 ( .A(n461), .B(n651), .ZN(G51) );
  NOR2_X2 U605 ( .A1(n650), .A2(n745), .ZN(n461) );
  NAND2_X1 U606 ( .A1(n364), .A2(n466), .ZN(n463) );
  INV_X1 U607 ( .A(n465), .ZN(n464) );
  INV_X1 U608 ( .A(n741), .ZN(n466) );
  NAND2_X1 U609 ( .A1(n741), .A2(n470), .ZN(n467) );
  NAND2_X1 U610 ( .A1(n470), .A2(G902), .ZN(n469) );
  XNOR2_X1 U611 ( .A(n481), .B(n480), .ZN(n731) );
  INV_X1 U612 ( .A(n756), .ZN(n480) );
  XNOR2_X1 U613 ( .A(n580), .B(n482), .ZN(n481) );
  XNOR2_X1 U614 ( .A(n572), .B(G113), .ZN(n482) );
  NAND2_X1 U615 ( .A1(n484), .A2(n483), .ZN(n487) );
  NAND2_X1 U616 ( .A1(n486), .A2(n485), .ZN(n484) );
  NAND2_X1 U617 ( .A1(n491), .A2(n490), .ZN(n489) );
  NOR2_X1 U618 ( .A1(n746), .A2(n681), .ZN(n679) );
  INV_X1 U619 ( .A(n681), .ZN(n490) );
  NOR2_X1 U620 ( .A1(n746), .A2(n492), .ZN(n491) );
  INV_X1 U621 ( .A(KEYINPUT2), .ZN(n492) );
  XNOR2_X1 U622 ( .A(n501), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U623 ( .A1(n730), .A2(G472), .ZN(n504) );
  XNOR2_X1 U624 ( .A(n734), .B(n509), .ZN(n735) );
  XNOR2_X1 U625 ( .A(n649), .B(n510), .ZN(n650) );
  XNOR2_X2 U626 ( .A(G116), .B(G119), .ZN(n520) );
  INV_X1 U627 ( .A(KEYINPUT3), .ZN(n519) );
  XNOR2_X1 U628 ( .A(n529), .B(G140), .ZN(n530) );
  XNOR2_X1 U629 ( .A(n571), .B(n516), .ZN(n517) );
  INV_X1 U630 ( .A(G469), .ZN(n534) );
  XNOR2_X1 U631 ( .A(n741), .B(KEYINPUT122), .ZN(n742) );
  XNOR2_X1 U632 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U633 ( .A(n511), .B(KEYINPUT14), .ZN(n512) );
  NAND2_X1 U634 ( .A1(G952), .A2(n512), .ZN(n715) );
  NOR2_X1 U635 ( .A1(G953), .A2(n715), .ZN(n617) );
  NAND2_X1 U636 ( .A1(G902), .A2(n512), .ZN(n513) );
  XOR2_X1 U637 ( .A(KEYINPUT92), .B(n513), .Z(n514) );
  NAND2_X1 U638 ( .A1(G953), .A2(n514), .ZN(n615) );
  NOR2_X1 U639 ( .A1(G900), .A2(n615), .ZN(n515) );
  NOR2_X1 U640 ( .A1(n617), .A2(n515), .ZN(n589) );
  XOR2_X1 U641 ( .A(G137), .B(KEYINPUT4), .Z(n516) );
  XNOR2_X1 U642 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n523) );
  XNOR2_X1 U643 ( .A(n523), .B(KEYINPUT78), .ZN(n524) );
  NAND2_X1 U644 ( .A1(n575), .A2(G210), .ZN(n525) );
  XNOR2_X1 U645 ( .A(G472), .B(KEYINPUT94), .ZN(n526) );
  XNOR2_X2 U646 ( .A(n527), .B(n526), .ZN(n688) );
  INV_X1 U647 ( .A(n591), .ZN(n634) );
  XNOR2_X1 U648 ( .A(n528), .B(KEYINPUT77), .ZN(n561) );
  NAND2_X1 U649 ( .A1(G214), .A2(n561), .ZN(n700) );
  NAND2_X1 U650 ( .A1(G227), .A2(n763), .ZN(n531) );
  XNOR2_X1 U651 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X2 U652 ( .A(n535), .B(n534), .ZN(n596) );
  XOR2_X1 U653 ( .A(KEYINPUT10), .B(KEYINPUT70), .Z(n537) );
  XOR2_X1 U654 ( .A(G110), .B(G119), .Z(n539) );
  XNOR2_X1 U655 ( .A(n539), .B(n538), .ZN(n540) );
  NAND2_X1 U656 ( .A1(G234), .A2(n763), .ZN(n541) );
  XNOR2_X1 U657 ( .A(n542), .B(n541), .ZN(n568) );
  NAND2_X1 U658 ( .A1(n568), .A2(G221), .ZN(n543) );
  XNOR2_X1 U659 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U660 ( .A1(n549), .A2(G217), .ZN(n547) );
  XOR2_X1 U661 ( .A(n550), .B(KEYINPUT21), .Z(n686) );
  XNOR2_X1 U662 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n553) );
  XNOR2_X1 U663 ( .A(n344), .B(n553), .ZN(n557) );
  XOR2_X1 U664 ( .A(n597), .B(KEYINPUT38), .Z(n701) );
  XOR2_X1 U665 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n563) );
  XNOR2_X1 U666 ( .A(G122), .B(KEYINPUT99), .ZN(n562) );
  XNOR2_X1 U667 ( .A(n565), .B(n564), .ZN(n566) );
  NAND2_X1 U668 ( .A1(G217), .A2(n568), .ZN(n569) );
  NOR2_X1 U669 ( .A1(G902), .A2(n736), .ZN(n570) );
  XNOR2_X1 U670 ( .A(G143), .B(n571), .ZN(n572) );
  XNOR2_X1 U671 ( .A(n574), .B(n573), .ZN(n579) );
  NAND2_X1 U672 ( .A1(G214), .A2(n575), .ZN(n576) );
  XNOR2_X1 U673 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U674 ( .A(n579), .B(n578), .Z(n580) );
  XNOR2_X1 U675 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n581) );
  NAND2_X1 U676 ( .A1(n584), .A2(n586), .ZN(n661) );
  NOR2_X1 U677 ( .A1(n585), .A2(n661), .ZN(n677) );
  NOR2_X1 U678 ( .A1(n586), .A2(n477), .ZN(n632) );
  NOR2_X1 U679 ( .A1(n611), .A2(n583), .ZN(n664) );
  NAND2_X1 U680 ( .A1(n586), .A2(n477), .ZN(n704) );
  NAND2_X1 U681 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U682 ( .A1(n704), .A2(n705), .ZN(n588) );
  XNOR2_X1 U683 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n587) );
  XNOR2_X1 U684 ( .A(n588), .B(n587), .ZN(n717) );
  NOR2_X1 U685 ( .A1(n589), .A2(n685), .ZN(n590) );
  NAND2_X1 U686 ( .A1(n590), .A2(n686), .ZN(n598) );
  NOR2_X1 U687 ( .A1(n598), .A2(n591), .ZN(n592) );
  XNOR2_X1 U688 ( .A(KEYINPUT28), .B(n592), .ZN(n593) );
  NAND2_X1 U689 ( .A1(n593), .A2(n596), .ZN(n605) );
  NOR2_X1 U690 ( .A1(n717), .A2(n605), .ZN(n595) );
  XNOR2_X1 U691 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n594) );
  XNOR2_X1 U692 ( .A(n595), .B(n594), .ZN(n771) );
  INV_X1 U693 ( .A(n691), .ZN(n623) );
  XOR2_X1 U694 ( .A(KEYINPUT89), .B(n623), .Z(n638) );
  NOR2_X1 U695 ( .A1(n598), .A2(n666), .ZN(n600) );
  XOR2_X1 U696 ( .A(KEYINPUT6), .B(n688), .Z(n627) );
  INV_X1 U697 ( .A(n627), .ZN(n599) );
  NAND2_X1 U698 ( .A1(n600), .A2(n599), .ZN(n608) );
  NAND2_X1 U699 ( .A1(n661), .A2(n602), .ZN(n603) );
  XOR2_X1 U700 ( .A(KEYINPUT100), .B(n603), .Z(n706) );
  XNOR2_X1 U701 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n604) );
  NOR2_X1 U702 ( .A1(n618), .A2(n605), .ZN(n606) );
  XNOR2_X1 U703 ( .A(n606), .B(KEYINPUT83), .ZN(n665) );
  NOR2_X1 U704 ( .A1(n706), .A2(n665), .ZN(n607) );
  NOR2_X1 U705 ( .A1(n362), .A2(n608), .ZN(n609) );
  NAND2_X1 U706 ( .A1(n609), .A2(n700), .ZN(n610) );
  XNOR2_X1 U707 ( .A(n610), .B(KEYINPUT43), .ZN(n612) );
  NAND2_X1 U708 ( .A1(n612), .A2(n611), .ZN(n678) );
  XOR2_X1 U709 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n614) );
  XNOR2_X1 U710 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n613) );
  XNOR2_X1 U711 ( .A(n614), .B(n613), .ZN(n622) );
  INV_X1 U712 ( .A(n704), .ZN(n620) );
  NOR2_X1 U713 ( .A1(G898), .A2(n615), .ZN(n616) );
  NAND2_X1 U714 ( .A1(n692), .A2(n691), .ZN(n624) );
  NAND2_X1 U715 ( .A1(n454), .A2(n628), .ZN(n625) );
  INV_X1 U716 ( .A(n628), .ZN(n629) );
  XOR2_X1 U717 ( .A(KEYINPUT34), .B(KEYINPUT82), .Z(n630) );
  XNOR2_X1 U718 ( .A(KEYINPUT73), .B(n630), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n767), .A2(KEYINPUT44), .ZN(n633) );
  NOR2_X1 U720 ( .A1(n634), .A2(n685), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U722 ( .A1(n362), .A2(n637), .ZN(n660) );
  XNOR2_X1 U723 ( .A(n639), .B(KEYINPUT103), .ZN(n640) );
  XNOR2_X1 U724 ( .A(KEYINPUT32), .B(n642), .ZN(n772) );
  NAND2_X1 U725 ( .A1(KEYINPUT68), .A2(n644), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n643), .A2(KEYINPUT44), .ZN(n645) );
  XOR2_X1 U727 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n648) );
  XNOR2_X1 U728 ( .A(KEYINPUT56), .B(KEYINPUT118), .ZN(n651) );
  XOR2_X1 U729 ( .A(G101), .B(n653), .Z(G3) );
  XOR2_X1 U730 ( .A(G104), .B(KEYINPUT111), .Z(n655) );
  INV_X1 U731 ( .A(n666), .ZN(n669) );
  NAND2_X1 U732 ( .A1(n656), .A2(n669), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(G6) );
  XOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n658) );
  INV_X1 U735 ( .A(n661), .ZN(n672) );
  NAND2_X1 U736 ( .A1(n656), .A2(n672), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U738 ( .A(G107), .B(n659), .ZN(G9) );
  XOR2_X1 U739 ( .A(G110), .B(n660), .Z(G12) );
  NOR2_X1 U740 ( .A1(n661), .A2(n665), .ZN(n663) );
  XNOR2_X1 U741 ( .A(G128), .B(KEYINPUT29), .ZN(n662) );
  XNOR2_X1 U742 ( .A(n663), .B(n662), .ZN(G30) );
  XOR2_X1 U743 ( .A(G143), .B(n664), .Z(G45) );
  NOR2_X1 U744 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U745 ( .A(G146), .B(n667), .Z(G48) );
  NAND2_X1 U746 ( .A1(n668), .A2(n669), .ZN(n670) );
  XNOR2_X1 U747 ( .A(n670), .B(KEYINPUT112), .ZN(n671) );
  XNOR2_X1 U748 ( .A(G113), .B(n671), .ZN(G15) );
  XOR2_X1 U749 ( .A(G116), .B(KEYINPUT113), .Z(n674) );
  NAND2_X1 U750 ( .A1(n668), .A2(n672), .ZN(n673) );
  XNOR2_X1 U751 ( .A(n674), .B(n673), .ZN(G18) );
  XNOR2_X1 U752 ( .A(G125), .B(n675), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n676), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U754 ( .A(G134), .B(n677), .Z(G36) );
  XNOR2_X1 U755 ( .A(G140), .B(n678), .ZN(G42) );
  XNOR2_X1 U756 ( .A(n680), .B(KEYINPUT2), .ZN(n684) );
  NAND2_X1 U757 ( .A1(n490), .A2(n746), .ZN(n682) );
  NAND2_X1 U758 ( .A1(KEYINPUT85), .A2(n682), .ZN(n683) );
  NOR2_X1 U759 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U760 ( .A(KEYINPUT49), .B(n687), .ZN(n689) );
  NAND2_X1 U761 ( .A1(n689), .A2(n454), .ZN(n690) );
  XNOR2_X1 U762 ( .A(KEYINPUT114), .B(n690), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n692), .A2(n362), .ZN(n693) );
  XNOR2_X1 U764 ( .A(n693), .B(KEYINPUT50), .ZN(n694) );
  NOR2_X1 U765 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U767 ( .A(KEYINPUT51), .B(n698), .Z(n699) );
  NOR2_X1 U768 ( .A1(n717), .A2(n699), .ZN(n711) );
  NOR2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U770 ( .A(KEYINPUT115), .B(n702), .Z(n703) );
  NOR2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U774 ( .A1(n716), .A2(n709), .ZN(n710) );
  NOR2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U776 ( .A(n712), .B(KEYINPUT116), .ZN(n713) );
  XNOR2_X1 U777 ( .A(KEYINPUT52), .B(n713), .ZN(n714) );
  NOR2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U779 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U781 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U782 ( .A(n723), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U783 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n724), .B(KEYINPUT57), .ZN(n725) );
  XNOR2_X1 U785 ( .A(n726), .B(n725), .ZN(n728) );
  NAND2_X1 U786 ( .A1(G469), .A2(n740), .ZN(n727) );
  XNOR2_X1 U787 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U788 ( .A1(n745), .A2(n729), .ZN(G54) );
  XNOR2_X1 U789 ( .A(KEYINPUT59), .B(KEYINPUT66), .ZN(n733) );
  XNOR2_X1 U790 ( .A(n731), .B(KEYINPUT120), .ZN(n732) );
  XOR2_X1 U791 ( .A(n736), .B(KEYINPUT121), .Z(n738) );
  NAND2_X1 U792 ( .A1(G478), .A2(n740), .ZN(n737) );
  XNOR2_X1 U793 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U794 ( .A1(n745), .A2(n739), .ZN(G63) );
  NAND2_X1 U795 ( .A1(n740), .A2(G217), .ZN(n743) );
  NOR2_X1 U796 ( .A1(n745), .A2(n744), .ZN(G66) );
  OR2_X1 U797 ( .A1(G953), .A2(n746), .ZN(n750) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n747) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n747), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n748), .A2(G898), .ZN(n749) );
  NAND2_X1 U801 ( .A1(n750), .A2(n749), .ZN(n754) );
  NOR2_X1 U802 ( .A1(G898), .A2(n763), .ZN(n751) );
  NOR2_X1 U803 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U804 ( .A(n754), .B(n753), .ZN(n755) );
  XOR2_X1 U805 ( .A(KEYINPUT123), .B(n755), .Z(G69) );
  XNOR2_X1 U806 ( .A(n757), .B(n756), .ZN(n761) );
  INV_X1 U807 ( .A(n761), .ZN(n758) );
  XOR2_X1 U808 ( .A(G227), .B(n758), .Z(n759) );
  NAND2_X1 U809 ( .A1(n759), .A2(G900), .ZN(n760) );
  NAND2_X1 U810 ( .A1(n760), .A2(G953), .ZN(n766) );
  XOR2_X1 U811 ( .A(n761), .B(n490), .Z(n762) );
  XNOR2_X1 U812 ( .A(n762), .B(KEYINPUT124), .ZN(n764) );
  NAND2_X1 U813 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U814 ( .A1(n766), .A2(n765), .ZN(G72) );
  XNOR2_X1 U815 ( .A(n767), .B(G122), .ZN(n768) );
  XNOR2_X1 U816 ( .A(n768), .B(KEYINPUT125), .ZN(G24) );
  XNOR2_X1 U817 ( .A(n769), .B(G131), .ZN(n770) );
  XNOR2_X1 U818 ( .A(n770), .B(KEYINPUT126), .ZN(G33) );
  XNOR2_X1 U819 ( .A(G137), .B(n771), .ZN(G39) );
  XOR2_X1 U820 ( .A(n772), .B(G119), .Z(G21) );
endmodule

