//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n591, new_n592, new_n593, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  INV_X1    g041(.A(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(G2104), .ZN(new_n468));
  OAI22_X1  g043(.A1(new_n465), .A2(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n463), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n461), .A2(new_n462), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n464), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n463), .A2(KEYINPUT66), .A3(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n476), .B(new_n480), .C1(G136), .C2(new_n485), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n465), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(KEYINPUT4), .A2(G138), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n461), .B2(new_n462), .ZN(new_n491));
  AND2_X1   g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n464), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n461), .B2(new_n462), .ZN(new_n495));
  AND2_X1   g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n489), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  AND3_X1   g081(.A1(KEYINPUT67), .A2(KEYINPUT6), .A3(G651), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT6), .B1(KEYINPUT67), .B2(G651), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n507), .A2(new_n508), .B1(new_n501), .B2(new_n502), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT67), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT67), .A2(KEYINPUT6), .A3(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n506), .A2(new_n511), .A3(KEYINPUT68), .A4(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI21_X1  g096(.A(G543), .B1(new_n507), .B2(new_n508), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n509), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT5), .B(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G62), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n527), .B2(new_n500), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n520), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(new_n529), .ZN(G166));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n522), .A2(KEYINPUT69), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n515), .A2(new_n516), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n533), .A2(new_n534), .A3(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n531), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n539));
  INV_X1    g114(.A(G89), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(new_n509), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(G168));
  NAND2_X1  g117(.A1(new_n510), .A2(G90), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n544));
  OAI21_X1  g119(.A(G64), .B1(new_n501), .B2(new_n502), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n544), .B1(new_n547), .B2(G651), .ZN(new_n548));
  AOI211_X1 g123(.A(KEYINPUT70), .B(new_n525), .C1(new_n545), .C2(new_n546), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n543), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n532), .A2(new_n535), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n551), .A2(G52), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(G171));
  AND2_X1   g128(.A1(new_n551), .A2(G43), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n555), .A2(new_n525), .B1(new_n556), .B2(new_n509), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT71), .Z(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n509), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n533), .A2(new_n526), .A3(KEYINPUT72), .A4(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n522), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n517), .A2(new_n572), .A3(G53), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n503), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n569), .A2(new_n574), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(KEYINPUT73), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n550), .B2(new_n552), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n547), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT70), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n547), .A2(new_n544), .A3(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n551), .A2(G52), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n585), .A2(KEYINPUT73), .A3(new_n586), .A4(new_n543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G301));
  NAND2_X1  g164(.A1(G168), .A2(KEYINPUT74), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(new_n536), .B2(new_n541), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G286));
  INV_X1    g169(.A(G166), .ZN(G303));
  NAND2_X1  g170(.A1(new_n517), .A2(G49), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n533), .A2(G87), .A3(new_n526), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G288));
  AND2_X1   g174(.A1(G73), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n526), .B2(G61), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n525), .ZN(new_n602));
  INV_X1    g177(.A(G86), .ZN(new_n603));
  INV_X1    g178(.A(G48), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n509), .A2(new_n603), .B1(new_n522), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G305));
  AND2_X1   g182(.A1(new_n551), .A2(G47), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n609), .A2(new_n525), .B1(new_n610), .B2(new_n509), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G290));
  AOI21_X1  g188(.A(new_n534), .B1(new_n533), .B2(G543), .ZN(new_n614));
  AOI211_X1 g189(.A(KEYINPUT69), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n615));
  OAI21_X1  g190(.A(G54), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n509), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n533), .A2(new_n526), .A3(KEYINPUT10), .A4(G92), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  INV_X1    g197(.A(G66), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n503), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G651), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n616), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n588), .B2(G868), .ZN(G284));
  AOI21_X1  g203(.A(new_n627), .B1(new_n588), .B2(G868), .ZN(G321));
  NOR2_X1   g204(.A1(G299), .A2(G868), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n593), .B2(G868), .ZN(G297));
  AOI21_X1  g206(.A(new_n630), .B1(new_n593), .B2(G868), .ZN(G280));
  AND3_X1   g207(.A1(new_n616), .A2(new_n621), .A3(new_n625), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT75), .B(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(G860), .B2(new_n634), .ZN(G148));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g214(.A1(new_n477), .A2(new_n468), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT12), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT76), .B(G2100), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT77), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n478), .A2(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n464), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  INV_X1    g223(.A(G135), .ZN(new_n649));
  OAI221_X1 g224(.A(new_n646), .B1(new_n647), .B2(new_n648), .C1(new_n484), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n642), .A2(new_n643), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT78), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n645), .A2(new_n651), .A3(new_n653), .ZN(G156));
  XOR2_X1   g229(.A(KEYINPUT15), .B(G2435), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2438), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT80), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(KEYINPUT14), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G14), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n665), .A2(new_n668), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT81), .Z(G401));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(KEYINPUT17), .ZN(new_n680));
  INV_X1    g255(.A(new_n674), .ZN(new_n681));
  INV_X1    g256(.A(new_n675), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n681), .A2(new_n677), .A3(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(new_n676), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n679), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2096), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1956), .B(G2474), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1961), .B(G1966), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(KEYINPUT83), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  NOR3_X1   g275(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1991), .B(G1996), .Z(new_n707));
  AOI21_X1  g282(.A(new_n704), .B1(new_n700), .B2(new_n703), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n707), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n700), .A2(new_n703), .ZN(new_n711));
  INV_X1    g286(.A(new_n704), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n710), .B1(new_n713), .B2(new_n705), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n690), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n707), .B1(new_n706), .B2(new_n708), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n710), .A3(new_n705), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n716), .A2(new_n689), .A3(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n715), .A2(new_n718), .ZN(G229));
  NOR2_X1   g294(.A1(G16), .A2(G23), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT86), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n722));
  NAND2_X1  g297(.A1(G288), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(KEYINPUT87), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n721), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT33), .B(G1976), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(G22), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G166), .B2(new_n726), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G1971), .ZN(new_n732));
  NOR2_X1   g307(.A1(G6), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n606), .B2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT32), .B(G1981), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n731), .A2(G1971), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n729), .A2(new_n732), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n612), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G16), .B2(G24), .ZN(new_n741));
  INV_X1    g316(.A(G1986), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT84), .B(G29), .Z(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G25), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n485), .A2(G131), .ZN(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n748));
  INV_X1    g323(.A(G107), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G2105), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n478), .B2(G119), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(new_n745), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT35), .B(G1991), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT85), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n741), .A2(new_n742), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n739), .A2(new_n743), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT88), .B(KEYINPUT36), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AND3_X1   g338(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT26), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n764), .B(new_n766), .C1(new_n478), .C2(G129), .ZN(new_n767));
  INV_X1    g342(.A(G141), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n484), .B2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G29), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n771), .B2(G32), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n745), .A2(G27), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n745), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT99), .B(G2078), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n775), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n771), .A2(G33), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n783));
  NAND2_X1  g358(.A1(G103), .A2(G2104), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G2105), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n788));
  INV_X1    g363(.A(G139), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n787), .B1(new_n464), .B2(new_n788), .C1(new_n484), .C2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n782), .B1(new_n790), .B2(G29), .ZN(new_n791));
  INV_X1    g366(.A(G2072), .ZN(new_n792));
  OAI21_X1  g367(.A(KEYINPUT90), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(G160), .A2(G29), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT24), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(G34), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n744), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G2084), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n792), .B2(new_n791), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n633), .A2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G4), .B2(G16), .ZN(new_n804));
  INV_X1    g379(.A(G1348), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT100), .B(G1956), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n726), .A2(G20), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT23), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n569), .A2(new_n574), .A3(new_n578), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n726), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n781), .A2(new_n793), .A3(new_n802), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n745), .A2(G35), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n745), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT29), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2090), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n791), .A2(new_n792), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n558), .A2(G16), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G16), .B2(G19), .ZN(new_n820));
  INV_X1    g395(.A(G1341), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n817), .A2(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n744), .A2(G26), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT28), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n478), .A2(G128), .ZN(new_n825));
  NOR2_X1   g400(.A1(G104), .A2(G2105), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT89), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n828));
  INV_X1    g403(.A(G140), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n825), .B1(new_n827), .B2(new_n828), .C1(new_n484), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n824), .B1(new_n830), .B2(G29), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G2067), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n822), .B(new_n832), .C1(new_n821), .C2(new_n820), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n812), .A2(new_n816), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n804), .A2(new_n805), .ZN(new_n835));
  INV_X1    g410(.A(G1961), .ZN(new_n836));
  NOR2_X1   g411(.A1(G5), .A2(G16), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT97), .ZN(new_n838));
  INV_X1    g413(.A(G171), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(new_n726), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n835), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n810), .A2(new_n806), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n773), .A2(new_n774), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT91), .Z(new_n844));
  NAND4_X1  g419(.A1(new_n834), .A2(new_n841), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n726), .A2(G21), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G168), .B2(new_n726), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT92), .B(G1966), .Z(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT96), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n840), .A2(new_n836), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n847), .A2(new_n849), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G11), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT30), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n771), .B1(new_n856), .B2(G28), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT94), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n857), .A2(new_n858), .B1(new_n856), .B2(G28), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n650), .B2(new_n744), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT95), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n851), .A2(new_n852), .A3(new_n853), .A4(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT98), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n845), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n763), .A2(new_n866), .ZN(G150));
  INV_X1    g442(.A(G150), .ZN(G311));
  AOI22_X1  g443(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(new_n525), .ZN(new_n870));
  INV_X1    g445(.A(G55), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n532), .B2(new_n535), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n510), .A2(G93), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT101), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(G55), .B1(new_n614), .B2(new_n615), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n510), .A2(G93), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n870), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT103), .B(G860), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n874), .A2(new_n878), .ZN(new_n883));
  INV_X1    g458(.A(new_n870), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n558), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n879), .A2(KEYINPUT102), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n879), .B2(KEYINPUT102), .ZN(new_n891));
  AOI211_X1 g466(.A(new_n886), .B(new_n870), .C1(new_n874), .C2(new_n878), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT38), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n633), .A2(G559), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n880), .B1(new_n897), .B2(KEYINPUT39), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n882), .B1(new_n900), .B2(new_n901), .ZN(G145));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n498), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n489), .A2(KEYINPUT105), .A3(new_n493), .A4(new_n497), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n830), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(new_n752), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n752), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n769), .A2(new_n790), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n769), .A2(new_n790), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G118), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n914), .A2(new_n915), .B1(new_n917), .B2(G2105), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n478), .A2(G130), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G142), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n484), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n641), .B(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n913), .A2(new_n922), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n910), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n650), .B(G160), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(G162), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n908), .A2(new_n923), .A3(new_n909), .A4(new_n924), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n928), .B1(new_n926), .B2(new_n929), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n934), .B(new_n935), .ZN(G395));
  XNOR2_X1  g511(.A(new_n894), .B(new_n636), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n809), .A2(new_n626), .A3(KEYINPUT108), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n633), .B2(G299), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n633), .B2(G299), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n809), .A2(KEYINPUT109), .A3(new_n626), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n633), .A2(new_n942), .A3(G299), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT109), .B1(new_n809), .B2(new_n626), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT108), .B1(new_n809), .B2(new_n626), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n633), .A2(new_n939), .A3(G299), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n948), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(new_n949), .B2(new_n950), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n943), .A2(new_n957), .A3(new_n944), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n941), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n955), .B1(new_n959), .B2(new_n948), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n947), .B1(new_n937), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n612), .B(G166), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n725), .B(G305), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n964), .B(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT42), .Z(new_n967));
  AND2_X1   g542(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n947), .B(KEYINPUT111), .C1(new_n937), .C2(new_n960), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(G868), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n879), .A2(G868), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(G295));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n972), .ZN(G331));
  NAND3_X1  g549(.A1(new_n581), .A2(new_n587), .A3(G168), .ZN(new_n975));
  NAND3_X1  g550(.A1(G171), .A2(new_n592), .A3(new_n590), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n891), .A2(new_n892), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n885), .A2(new_n888), .A3(new_n886), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n975), .A2(new_n976), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n890), .A2(new_n981), .A3(new_n893), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(new_n960), .ZN(new_n984));
  INV_X1    g559(.A(new_n946), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n980), .B2(new_n982), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n966), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n978), .A2(new_n979), .A3(new_n977), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n981), .B1(new_n890), .B2(new_n893), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n946), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n966), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n990), .B(new_n991), .C1(new_n960), .C2(new_n983), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n987), .A2(new_n931), .A3(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT113), .B(KEYINPUT43), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n946), .B1(new_n983), .B2(new_n948), .ZN(new_n997));
  INV_X1    g572(.A(new_n959), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n998), .A2(new_n980), .A3(KEYINPUT41), .A4(new_n982), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n991), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n1000), .A2(new_n987), .A3(new_n931), .A4(new_n994), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n987), .A3(new_n931), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1006), .B(KEYINPUT44), .C1(new_n993), .C2(new_n995), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(G397));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  INV_X1    g584(.A(G40), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n469), .A2(new_n472), .A3(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1009), .B(new_n1011), .C1(new_n906), .C2(G1384), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT114), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n830), .B(G2067), .ZN(new_n1014));
  INV_X1    g589(.A(G1996), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n770), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1012), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1015), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n769), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n752), .B(new_n756), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1021), .B2(new_n1013), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G290), .A2(G1986), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT48), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1019), .B(KEYINPUT46), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1013), .B1(new_n769), .B2(new_n1014), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT47), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  OR3_X1    g606(.A1(new_n1020), .A2(new_n756), .A3(new_n752), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n830), .A2(G2067), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1031), .B1(new_n1013), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n519), .A2(new_n529), .A3(G8), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n469), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n470), .A2(new_n471), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G2105), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n1042), .A3(G40), .ZN(new_n1043));
  INV_X1    g618(.A(G1384), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n498), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1045), .B2(new_n1009), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n904), .A2(KEYINPUT45), .A3(new_n1044), .A4(new_n905), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1971), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(KEYINPUT50), .ZN(new_n1051));
  INV_X1    g626(.A(G2090), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n498), .A2(new_n1053), .A3(new_n1044), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1051), .A2(new_n1052), .A3(new_n1011), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1050), .A2(KEYINPUT119), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G8), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT119), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1039), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1055), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1971), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1061));
  OAI211_X1 g636(.A(G8), .B(new_n1038), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1050), .A2(new_n1055), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(new_n1065), .A3(G8), .A4(new_n1038), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G8), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n498), .A2(new_n1044), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(new_n1069), .B2(new_n1011), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT116), .A4(G1976), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n1072));
  INV_X1    g647(.A(G1976), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n725), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n601), .A2(new_n525), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n510), .A2(G86), .ZN(new_n1081));
  INV_X1    g656(.A(G1981), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n517), .A2(G48), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(G1981), .B1(new_n602), .B2(new_n605), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT49), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT118), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1011), .A2(new_n1044), .A3(new_n498), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1088), .A2(new_n1089), .A3(G8), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT118), .A3(new_n1086), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1079), .A2(KEYINPUT52), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1078), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1051), .A2(new_n1011), .A3(new_n1054), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n1044), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1011), .B(new_n1098), .C1(new_n1069), .C2(KEYINPUT45), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1097), .A2(new_n800), .B1(new_n1099), .B2(new_n848), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1100), .A2(new_n1068), .A3(G286), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1059), .A2(new_n1067), .A3(new_n1095), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1101), .A2(KEYINPUT63), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1064), .A2(G8), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1039), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1105), .A2(new_n1067), .A3(new_n1095), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G168), .A2(new_n1068), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT51), .B1(new_n1110), .B2(KEYINPUT123), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(new_n1112), .C1(new_n1100), .C2(new_n1068), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1112), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1099), .A2(new_n848), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1051), .A2(new_n800), .A3(new_n1011), .A4(new_n1054), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G168), .ZN(new_n1118));
  OAI211_X1 g693(.A(G8), .B(new_n1114), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1110), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT62), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1059), .A2(new_n1067), .A3(new_n1095), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1048), .B2(G2078), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1096), .A2(new_n836), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1125), .A2(G2078), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1046), .A2(new_n1128), .A3(new_n1098), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n588), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1113), .A2(new_n1119), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1123), .A2(new_n1124), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1067), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1138));
  OR2_X1    g713(.A1(G288), .A2(G1976), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1084), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1137), .A2(new_n1095), .B1(new_n1140), .B2(new_n1070), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1109), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1009), .B1(new_n906), .B2(G1384), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1143), .A2(new_n1047), .A3(new_n1011), .A4(new_n1128), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1126), .A2(new_n1144), .A3(G301), .A4(new_n1127), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n1131), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1133), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1130), .A2(new_n588), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1126), .A2(new_n1144), .A3(new_n1127), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT124), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(G171), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(KEYINPUT124), .ZN(new_n1152));
  OAI211_X1 g727(.A(KEYINPUT54), .B(new_n1148), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1147), .A2(new_n1124), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(G1956), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1096), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT56), .B(G2072), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1046), .A2(new_n1047), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n1162));
  AOI22_X1  g737(.A1(new_n567), .A2(new_n568), .B1(G651), .B2(new_n577), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n574), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n809), .A2(KEYINPUT57), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1161), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1089), .ZN(new_n1172));
  INV_X1    g747(.A(G2067), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1096), .A2(new_n805), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1174), .A2(new_n626), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1169), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1171), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n626), .B1(new_n1174), .B2(KEYINPUT60), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(KEYINPUT60), .B2(new_n1174), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1171), .A2(new_n1176), .A3(KEYINPUT61), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT58), .B(G1341), .ZN(new_n1183));
  OAI22_X1  g758(.A1(new_n1048), .A2(G1996), .B1(new_n1172), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n558), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1184), .A2(KEYINPUT59), .A3(new_n558), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n626), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1182), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1171), .A2(new_n1176), .A3(KEYINPUT122), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1161), .A2(new_n1170), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1192), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1178), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1142), .B1(new_n1156), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n612), .A2(new_n742), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1018), .B1(new_n1023), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1022), .A2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1035), .B1(new_n1199), .B2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g778(.A(G319), .ZN(new_n1205));
  NOR2_X1   g779(.A1(G227), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g780(.A(new_n1206), .B1(new_n670), .B2(new_n671), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1207), .B1(new_n715), .B2(new_n718), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1208), .B1(new_n932), .B2(new_n933), .ZN(new_n1209));
  INV_X1    g783(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g784(.A(KEYINPUT126), .B1(new_n1002), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n1212));
  AOI211_X1 g786(.A(new_n1212), .B(new_n1209), .C1(new_n996), .C2(new_n1001), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n1211), .A2(new_n1213), .ZN(G308));
  NAND2_X1  g788(.A1(new_n1002), .A2(new_n1210), .ZN(G225));
endmodule


