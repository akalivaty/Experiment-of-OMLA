//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT22), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(G137), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(G125), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n196), .B1(new_n200), .B2(new_n194), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT73), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n201), .A2(new_n202), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT73), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n206), .A3(new_n202), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT24), .B(G110), .Z(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G110), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n210), .B(KEYINPUT23), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(new_n212), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n208), .B(new_n216), .C1(new_n217), .C2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n217), .A3(new_n212), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT74), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n218), .A2(KEYINPUT74), .A3(new_n217), .A4(new_n212), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n223), .B(new_n224), .C1(new_n214), .C2(new_n215), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n201), .A2(new_n202), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n200), .A2(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n193), .B1(new_n220), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n220), .A2(new_n229), .A3(new_n193), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT75), .B(KEYINPUT25), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n231), .A2(new_n188), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n232), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n235), .A2(new_n230), .A3(G902), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT25), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n189), .B(new_n234), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n235), .A2(new_n230), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n189), .A2(G902), .ZN(new_n241));
  XOR2_X1   g055(.A(new_n241), .B(KEYINPUT76), .Z(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT77), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n239), .A2(new_n246), .A3(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(G472), .A2(G902), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT72), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT31), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT70), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n211), .B2(G116), .ZN(new_n255));
  INV_X1    g069(.A(G116), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT67), .A3(G119), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n255), .A2(new_n257), .B1(G116), .B2(new_n211), .ZN(new_n258));
  XOR2_X1   g072(.A(KEYINPUT2), .B(G113), .Z(new_n259));
  OR2_X1    g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(KEYINPUT68), .A3(new_n259), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT68), .B1(new_n258), .B2(new_n259), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G137), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT11), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(G137), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT11), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n266), .B(new_n271), .C1(new_n267), .C2(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G131), .ZN(new_n274));
  INV_X1    g088(.A(G131), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n269), .A2(new_n275), .A3(new_n270), .A4(new_n272), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(KEYINPUT66), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT66), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(new_n278), .A3(G131), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n202), .A2(G143), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G143), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G146), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n202), .A2(KEYINPUT64), .A3(G143), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(KEYINPUT0), .A2(G128), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n280), .A2(new_n284), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n286), .A2(new_n290), .B1(new_n291), .B2(new_n288), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n277), .A2(new_n279), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n209), .B1(new_n280), .B2(KEYINPUT1), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n286), .A2(new_n295), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n270), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n267), .A2(G137), .ZN(new_n300));
  OAI21_X1  g114(.A(G131), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n276), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n265), .A2(new_n293), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n265), .B1(new_n293), .B2(new_n302), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT28), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT28), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G237), .A2(G953), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G210), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n311), .B(KEYINPUT27), .Z(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT26), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(G101), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n253), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n252), .A2(KEYINPUT70), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n293), .A2(new_n302), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT30), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT69), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(KEYINPUT30), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n293), .A2(new_n302), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n304), .B1(new_n324), .B2(new_n264), .ZN(new_n325));
  INV_X1    g139(.A(new_n314), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n316), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n265), .B1(new_n319), .B2(new_n323), .ZN(new_n328));
  INV_X1    g142(.A(new_n316), .ZN(new_n329));
  NOR4_X1   g143(.A1(new_n328), .A2(new_n304), .A3(new_n314), .A4(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n315), .B(KEYINPUT71), .C1(new_n327), .C2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  AOI211_X1 g146(.A(KEYINPUT69), .B(new_n320), .C1(new_n293), .C2(new_n302), .ZN(new_n333));
  AND4_X1   g147(.A1(new_n293), .A2(new_n302), .A3(new_n321), .A4(new_n322), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n264), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n303), .A3(new_n326), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n329), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n325), .A2(new_n326), .A3(new_n316), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT71), .B1(new_n339), .B2(new_n315), .ZN(new_n340));
  OAI211_X1 g154(.A(KEYINPUT32), .B(new_n251), .C1(new_n332), .C2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n306), .A2(new_n326), .A3(KEYINPUT29), .A4(new_n308), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n309), .B2(new_n314), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n325), .A2(new_n326), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n188), .B(new_n342), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G472), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n315), .B1(new_n327), .B2(new_n330), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n331), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT32), .B1(new_n352), .B2(new_n251), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n248), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G110), .B(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n190), .A2(G227), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n357), .B(KEYINPUT78), .Z(new_n358));
  INV_X1    g172(.A(KEYINPUT12), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n277), .A2(new_n279), .ZN(new_n360));
  INV_X1    g174(.A(G107), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G104), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(KEYINPUT79), .A2(G107), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT79), .A2(G107), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G101), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT80), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n291), .A2(new_n296), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n371), .B1(new_n291), .B2(new_n294), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n373), .B(G104), .C1(new_n364), .C2(new_n365), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n367), .A2(G107), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n362), .A2(KEYINPUT3), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n374), .A2(new_n369), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n361), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT79), .A2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n367), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n362), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(G101), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n370), .A2(new_n372), .A3(new_n377), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n370), .A2(new_n377), .A3(new_n384), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n297), .ZN(new_n387));
  AOI211_X1 g201(.A(new_n359), .B(new_n360), .C1(new_n385), .C2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n383), .B1(new_n382), .B2(G101), .ZN(new_n391));
  AOI211_X1 g205(.A(KEYINPUT80), .B(new_n369), .C1(new_n381), .C2(new_n362), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n298), .B1(new_n393), .B2(new_n377), .ZN(new_n394));
  INV_X1    g208(.A(new_n385), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n360), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n387), .A2(KEYINPUT82), .A3(new_n385), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n399), .A2(new_n400), .A3(new_n359), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n399), .B2(new_n359), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n389), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n370), .A2(new_n377), .A3(new_n384), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT10), .A3(new_n298), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G101), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT4), .A3(new_n377), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n409), .A3(G101), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n292), .A3(new_n410), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n412));
  OAI211_X1 g226(.A(new_n405), .B(new_n411), .C1(new_n395), .C2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n397), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n358), .B1(new_n403), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n357), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n413), .A2(new_n397), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n188), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G469), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n357), .B1(new_n415), .B2(new_n420), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n387), .A2(KEYINPUT82), .A3(new_n385), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT82), .B1(new_n387), .B2(new_n385), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n427), .A2(new_n428), .A3(new_n360), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT83), .B1(new_n429), .B2(KEYINPUT12), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n399), .A2(new_n400), .A3(new_n359), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n388), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n426), .B1(new_n432), .B2(new_n419), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT84), .B(G469), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n188), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n424), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(KEYINPUT9), .B(G234), .Z(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G221), .B1(new_n438), .B2(G902), .ZN(new_n439));
  OAI21_X1  g253(.A(G214), .B1(G237), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n292), .A2(G125), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(G125), .B2(new_n297), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n190), .A2(G224), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n443), .B(new_n444), .Z(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT85), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n258), .A2(new_n259), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT68), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n256), .A2(KEYINPUT5), .A3(G119), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n258), .B2(KEYINPUT5), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n451), .A2(new_n261), .B1(new_n453), .B2(G113), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n404), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n264), .A2(new_n410), .A3(new_n408), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n448), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT86), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n456), .A3(new_n448), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT6), .A4(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n460), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n462), .A2(new_n457), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT86), .B1(new_n457), .B2(new_n463), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n445), .B(new_n461), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n453), .A2(G113), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n262), .B2(new_n263), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(new_n404), .A3(KEYINPUT87), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n454), .B1(new_n386), .B2(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n447), .A2(KEYINPUT8), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n447), .A2(KEYINPUT8), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n443), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n444), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n444), .A2(new_n477), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n443), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n474), .A2(new_n478), .A3(new_n460), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n188), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(KEYINPUT89), .A3(new_n188), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n466), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G210), .B1(G237), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n466), .A2(new_n484), .A3(new_n487), .A4(new_n485), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n441), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT96), .ZN(new_n492));
  INV_X1    g306(.A(G122), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n493), .A2(KEYINPUT92), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(KEYINPUT92), .ZN(new_n495));
  OAI21_X1  g309(.A(G116), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n256), .A2(G122), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n496), .B(new_n497), .C1(new_n365), .C2(new_n364), .ZN(new_n498));
  INV_X1    g312(.A(new_n496), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n497), .B(KEYINPUT14), .ZN(new_n500));
  OAI21_X1  g314(.A(G107), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n209), .B2(G143), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n283), .A2(KEYINPUT93), .A3(G128), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n209), .A2(G143), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n509), .A2(new_n267), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n505), .A2(new_n507), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT95), .ZN(new_n513));
  AOI21_X1  g327(.A(G134), .B1(new_n513), .B2(new_n508), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n498), .B(new_n501), .C1(new_n511), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n496), .A2(new_n497), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n366), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n498), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n267), .B1(new_n509), .B2(new_n510), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT13), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n505), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n505), .B2(new_n520), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT94), .A4(KEYINPUT13), .ZN(new_n524));
  AND4_X1   g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .A4(new_n507), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n518), .B(new_n519), .C1(new_n525), .C2(new_n267), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n438), .A2(new_n187), .A3(G953), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n515), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n515), .B2(new_n526), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n492), .B(new_n188), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT15), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n530), .A2(new_n531), .A3(G478), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n188), .B1(new_n528), .B2(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT96), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n530), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(G478), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n190), .A2(G952), .ZN(new_n538));
  NAND2_X1  g352(.A1(G234), .A2(G237), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT97), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT21), .B(G898), .Z(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(G902), .A3(G953), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G475), .ZN(new_n545));
  AOI21_X1  g359(.A(G143), .B1(new_n310), .B2(G214), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n310), .A2(G143), .A3(G214), .ZN(new_n548));
  NAND2_X1  g362(.A1(KEYINPUT18), .A2(G131), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n548), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT18), .B(G131), .C1(new_n551), .C2(new_n546), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n197), .A2(new_n199), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT91), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n200), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n202), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n550), .B(new_n552), .C1(new_n557), .C2(new_n227), .ZN(new_n558));
  OAI21_X1  g372(.A(G131), .B1(new_n551), .B2(new_n546), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n547), .A2(new_n275), .A3(new_n548), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n561), .B2(new_n559), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n558), .B1(new_n563), .B2(new_n208), .ZN(new_n564));
  XNOR2_X1  g378(.A(G113), .B(G122), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(new_n367), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n566), .B(new_n558), .C1(new_n563), .C2(new_n208), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n545), .B1(new_n570), .B2(new_n188), .ZN(new_n571));
  INV_X1    g385(.A(new_n569), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n226), .B1(new_n559), .B2(new_n560), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT19), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n553), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n200), .B(KEYINPUT91), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n202), .B(new_n575), .C1(new_n576), .C2(new_n574), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n566), .B1(new_n578), .B2(new_n558), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n545), .B(new_n188), .C1(new_n572), .C2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n578), .A2(new_n558), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n569), .B1(new_n583), .B2(new_n566), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT20), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n545), .A4(new_n188), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n571), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n537), .A2(KEYINPUT98), .A3(new_n544), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n515), .A2(new_n526), .ZN(new_n589));
  INV_X1    g403(.A(new_n527), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n515), .A2(new_n526), .A3(new_n527), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n492), .B1(new_n593), .B2(new_n188), .ZN(new_n594));
  INV_X1    g408(.A(new_n530), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n536), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n530), .A2(new_n531), .A3(G478), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(new_n587), .A3(new_n544), .A4(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n588), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n436), .A2(new_n439), .A3(new_n491), .A4(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n354), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n369), .ZN(G3));
  AOI21_X1  g418(.A(new_n250), .B1(new_n351), .B2(new_n331), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n188), .B1(new_n332), .B2(new_n340), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n606), .B2(G472), .ZN(new_n607));
  INV_X1    g421(.A(new_n439), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n424), .B2(new_n435), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n491), .A2(new_n248), .A3(new_n544), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n590), .B2(KEYINPUT99), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n593), .B(new_n612), .Z(new_n613));
  NAND2_X1  g427(.A1(new_n188), .A2(G478), .ZN(new_n614));
  INV_X1    g428(.A(new_n593), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(G902), .ZN(new_n616));
  OAI22_X1  g430(.A1(new_n613), .A2(new_n614), .B1(G478), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n587), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n607), .A2(new_n609), .A3(new_n610), .A4(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  INV_X1    g437(.A(new_n537), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n580), .A2(new_n581), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n571), .B1(new_n625), .B2(new_n582), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n607), .A2(new_n609), .A3(new_n610), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NAND2_X1  g445(.A1(new_n220), .A2(new_n229), .ZN(new_n632));
  INV_X1    g446(.A(new_n193), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n632), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n242), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n239), .A2(new_n636), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n491), .A2(new_n600), .A3(new_n588), .A4(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n607), .A3(new_n609), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT100), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(G12));
  INV_X1    g456(.A(new_n347), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n605), .B2(KEYINPUT32), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT32), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n332), .A2(new_n340), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n645), .B1(new_n646), .B2(new_n250), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n491), .A2(new_n637), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n541), .B1(G900), .B2(new_n543), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n628), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n648), .A2(new_n609), .A3(new_n649), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  XNOR2_X1  g468(.A(new_n650), .B(KEYINPUT101), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT39), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n609), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT40), .Z(new_n658));
  NOR2_X1   g472(.A1(new_n325), .A2(new_n314), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n304), .A2(new_n305), .ZN(new_n660));
  AOI21_X1  g474(.A(G902), .B1(new_n660), .B2(new_n314), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n353), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n665), .A2(new_n341), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n637), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n489), .A2(new_n490), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT38), .Z(new_n669));
  NOR2_X1   g483(.A1(new_n537), .A2(new_n587), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n440), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n658), .A2(new_n667), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  OAI211_X1 g488(.A(new_n609), .B(new_n649), .C1(new_n348), .C2(new_n353), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n620), .A2(new_n650), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(KEYINPUT102), .A3(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n648), .A2(new_n609), .A3(new_n649), .A4(new_n678), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  INV_X1    g498(.A(new_n248), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n644), .B2(new_n647), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n425), .B1(new_n403), .B2(new_n418), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n687), .B1(new_n688), .B2(G902), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n433), .A2(KEYINPUT103), .A3(new_n188), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n690), .A3(G469), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n439), .A3(new_n435), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT104), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n491), .A2(new_n544), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n691), .A2(new_n695), .A3(new_n439), .A4(new_n435), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n686), .A2(new_n693), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n619), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT41), .B(G113), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  AND3_X1   g514(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n701), .A2(new_n702), .A3(new_n686), .A4(new_n628), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT105), .B1(new_n697), .B2(new_n627), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  AND3_X1   g520(.A1(new_n691), .A2(new_n439), .A3(new_n435), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n648), .A2(new_n707), .A3(new_n638), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT106), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n211), .ZN(G21));
  NAND4_X1  g524(.A1(new_n693), .A2(new_n694), .A3(new_n670), .A4(new_n696), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n250), .B1(new_n339), .B2(new_n315), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n606), .B2(G472), .ZN(new_n713));
  INV_X1    g527(.A(new_n244), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n493), .ZN(G24));
  INV_X1    g531(.A(new_n637), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n718), .B(new_n712), .C1(new_n606), .C2(G472), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n707), .A3(new_n491), .A4(new_n678), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n423), .B2(G469), .ZN(new_n723));
  INV_X1    g537(.A(new_n358), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n724), .B1(new_n432), .B2(new_n414), .ZN(new_n725));
  INV_X1    g539(.A(new_n422), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n722), .A2(new_n188), .A3(G469), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n435), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n668), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n608), .A2(new_n441), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n730), .A2(KEYINPUT108), .A3(new_n731), .A4(new_n732), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n686), .A3(new_n678), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n647), .B(KEYINPUT109), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n244), .B1(new_n741), .B2(new_n644), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n737), .A2(new_n742), .A3(KEYINPUT42), .A4(new_n678), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  OR3_X1    g559(.A1(new_n416), .A2(new_n422), .A3(new_n728), .ZN(new_n746));
  INV_X1    g560(.A(G469), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n727), .B2(new_n188), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n748), .B2(new_n722), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n668), .B1(new_n749), .B2(new_n435), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT108), .B1(new_n750), .B2(new_n732), .ZN(new_n751));
  INV_X1    g565(.A(new_n736), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n686), .B(new_n652), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT110), .B(G134), .Z(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G36));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n727), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n725), .A2(KEYINPUT45), .A3(new_n726), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n758), .A3(G469), .ZN(new_n759));
  NAND2_X1  g573(.A1(G469), .A2(G902), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n760), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n435), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n439), .A3(new_n656), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n668), .A2(new_n441), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n617), .A2(new_n587), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT43), .Z(new_n771));
  INV_X1    g585(.A(new_n607), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n637), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n768), .A2(new_n769), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  NAND2_X1  g592(.A1(new_n765), .A2(new_n439), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n648), .A2(new_n248), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n678), .A3(new_n769), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT112), .Z(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n698), .A2(new_n716), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n705), .A2(new_n789), .A3(new_n708), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n719), .A2(new_n678), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n751), .B2(new_n752), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n753), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n537), .A2(new_n618), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n607), .A2(new_n609), .A3(new_n610), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n639), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n603), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n639), .A3(KEYINPUT113), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n769), .A2(new_n626), .A3(new_n650), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n624), .A2(new_n718), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n648), .A2(new_n800), .A3(new_n609), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n798), .A2(new_n621), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n793), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n790), .A2(new_n804), .A3(new_n744), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n720), .A2(new_n653), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n718), .A2(new_n439), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n665), .B2(new_n341), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n731), .A2(new_n671), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n650), .A4(new_n730), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n720), .A2(new_n653), .A3(KEYINPUT114), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n683), .A2(new_n808), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n806), .B1(new_n679), .B2(new_n682), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n812), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n788), .B1(new_n805), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT115), .ZN(new_n821));
  INV_X1    g635(.A(new_n805), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n720), .A2(new_n653), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n680), .A2(new_n681), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n680), .A2(new_n681), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n823), .B(new_n812), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n818), .A3(KEYINPUT116), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n817), .B1(new_n816), .B2(new_n812), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n822), .A2(KEYINPUT53), .A3(new_n828), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n834), .B(new_n788), .C1(new_n805), .C2(new_n819), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n821), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n830), .B1(KEYINPUT52), .B2(new_n814), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n799), .A2(new_n621), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT113), .B1(new_n795), .B2(new_n639), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n839), .A2(new_n603), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n753), .A3(new_n802), .A4(new_n792), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n788), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n739), .B(new_n677), .C1(new_n735), .C2(new_n736), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n742), .A2(new_n846), .B1(new_n738), .B2(new_n739), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n705), .A2(new_n789), .A3(new_n708), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n804), .A2(KEYINPUT117), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n832), .A2(new_n849), .A3(new_n804), .A4(new_n828), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n845), .A2(new_n851), .B1(new_n852), .B2(new_n788), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n837), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n707), .A2(new_n769), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT120), .Z(new_n858));
  INV_X1    g672(.A(new_n541), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n248), .A2(new_n858), .A3(new_n859), .A4(new_n666), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n620), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n858), .A2(new_n859), .A3(new_n771), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT48), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n862), .A2(new_n863), .A3(new_n742), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n862), .B2(new_n742), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n538), .B(new_n861), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n617), .A2(new_n618), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n771), .A2(new_n859), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n715), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n441), .A3(new_n669), .A4(new_n707), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT50), .Z(new_n872));
  NAND2_X1  g686(.A1(new_n862), .A2(new_n719), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n868), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n691), .A2(new_n435), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n608), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n780), .B2(new_n781), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n769), .A3(new_n870), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n878), .A2(KEYINPUT51), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n866), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n870), .A2(new_n491), .A3(new_n707), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n883), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n874), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n880), .B(new_n881), .C1(new_n882), .C2(new_n886), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n856), .A2(new_n887), .B1(G952), .B2(G953), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n666), .A2(new_n714), .A3(new_n669), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT49), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n875), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n770), .B1(new_n875), .B2(new_n890), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n889), .A2(new_n732), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n888), .A2(new_n893), .ZN(G75));
  NAND2_X1  g708(.A1(new_n852), .A2(new_n788), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n838), .A2(new_n844), .A3(new_n849), .A4(new_n850), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(G210), .A3(G902), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n445), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n898), .B2(new_n899), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n190), .A2(G952), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(G51));
  XOR2_X1   g720(.A(new_n760), .B(KEYINPUT57), .Z(new_n907));
  AND3_X1   g721(.A1(new_n895), .A2(new_n854), .A3(new_n896), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n854), .B1(new_n895), .B2(new_n896), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n433), .ZN(new_n911));
  OR3_X1    g725(.A1(new_n853), .A2(new_n188), .A3(new_n759), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n905), .B1(new_n911), .B2(new_n912), .ZN(G54));
  INV_X1    g727(.A(KEYINPUT58), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT121), .B1(new_n914), .B2(new_n545), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n914), .A2(new_n545), .A3(KEYINPUT121), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n897), .A2(G902), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n584), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n905), .ZN(G60));
  INV_X1    g735(.A(new_n613), .ZN(new_n922));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT59), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n922), .B1(new_n856), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n922), .B(new_n924), .C1(new_n908), .C2(new_n909), .ZN(new_n926));
  INV_X1    g740(.A(new_n905), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n925), .A2(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT60), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n827), .A2(new_n818), .A3(KEYINPUT116), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT116), .B1(new_n827), .B2(new_n818), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT53), .B1(new_n935), .B2(new_n822), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n849), .A2(new_n838), .A3(new_n844), .A4(new_n850), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n240), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n897), .A2(new_n635), .A3(new_n932), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n927), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT61), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n905), .B1(new_n938), .B2(new_n939), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n946), .B(new_n941), .C1(new_n943), .C2(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(G66));
  AOI21_X1  g762(.A(new_n190), .B1(new_n542), .B2(G224), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n790), .A2(new_n841), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n949), .B1(new_n950), .B2(new_n190), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n900), .B1(G898), .B2(new_n190), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n951), .B(new_n952), .Z(G69));
  MUX2_X1   g767(.A(new_n200), .B(new_n576), .S(KEYINPUT19), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n324), .B(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n768), .A2(new_n742), .A3(new_n811), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n777), .A2(new_n957), .A3(new_n786), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n744), .A2(new_n753), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT124), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n808), .A2(new_n813), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n961), .A2(new_n683), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n744), .A2(new_n963), .A3(new_n753), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n958), .A2(new_n960), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n956), .B1(new_n965), .B2(new_n190), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(G227), .B2(new_n190), .ZN(new_n967));
  OAI21_X1  g781(.A(G900), .B1(new_n955), .B2(G227), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(G953), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n777), .A2(new_n786), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n961), .A2(new_n673), .A3(new_n683), .ZN(new_n971));
  XOR2_X1   g785(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n657), .A2(new_n441), .A3(new_n668), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n974), .B(new_n686), .C1(new_n620), .C2(new_n794), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n962), .B(new_n673), .C1(KEYINPUT123), .C2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n970), .A2(new_n973), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n190), .A3(new_n956), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n967), .A2(new_n969), .A3(new_n979), .ZN(G72));
  NAND2_X1  g794(.A1(G472), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT63), .Z(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT125), .Z(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n965), .B2(new_n950), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n314), .A3(new_n325), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n978), .B2(new_n950), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n905), .B1(new_n986), .B2(new_n659), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT126), .B1(new_n325), .B2(new_n326), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(new_n345), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n836), .A2(new_n990), .A3(new_n982), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n988), .B1(new_n993), .B2(new_n994), .ZN(G57));
endmodule


