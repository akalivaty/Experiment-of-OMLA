//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n632, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  XNOR2_X1  g002(.A(KEYINPUT66), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT67), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n457));
  OAI21_X1  g032(.A(KEYINPUT70), .B1(new_n457), .B2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT70), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n457), .A2(G2104), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n463), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n458), .A2(new_n461), .A3(new_n465), .A4(new_n462), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT71), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n460), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT72), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT72), .ZN(new_n474));
  INV_X1    g049(.A(new_n472), .ZN(new_n475));
  AOI211_X1 g050(.A(new_n474), .B(new_n475), .C1(new_n466), .C2(new_n469), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(new_n462), .A3(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT68), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n480), .A2(KEYINPUT68), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(KEYINPUT69), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n477), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NAND4_X1  g064(.A1(new_n458), .A2(new_n461), .A3(G2105), .A4(new_n462), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n465), .A2(G112), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND4_X1   g069(.A1(new_n465), .A2(new_n458), .A3(new_n461), .A4(new_n462), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(G136), .B2(new_n495), .ZN(G162));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  AND4_X1   g074(.A1(G2105), .A2(new_n458), .A3(new_n461), .A4(new_n462), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G126), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n458), .A2(new_n461), .A3(new_n462), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n478), .A2(new_n462), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n502), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n501), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n504), .A2(KEYINPUT4), .B1(new_n506), .B2(new_n507), .ZN(new_n512));
  INV_X1    g087(.A(new_n497), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(G114), .B2(new_n465), .ZN(new_n514));
  INV_X1    g089(.A(G126), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n490), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT73), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G62), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(KEYINPUT74), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n526), .A3(G62), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n520), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n522), .ZN(new_n536));
  NOR2_X1   g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n536), .A2(new_n537), .B1(new_n531), .B2(new_n532), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n535), .A2(G50), .B1(G88), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n540), .B1(new_n528), .B2(new_n529), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n530), .A2(new_n541), .ZN(G303));
  INV_X1    g117(.A(G303), .ZN(G166));
  NAND2_X1  g118(.A1(new_n535), .A2(G51), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n539), .A2(G89), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT76), .Z(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(G168));
  INV_X1    g127(.A(G52), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n534), .A2(new_n553), .B1(new_n554), .B2(new_n538), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n520), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(G171));
  AND2_X1   g133(.A1(new_n523), .A2(G56), .ZN(new_n559));
  AND2_X1   g134(.A1(G68), .A2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n535), .A2(G43), .B1(G81), .B2(new_n539), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G53), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n534), .A2(KEYINPUT9), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n534), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(new_n523), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(G91), .B2(new_n539), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  AND2_X1   g160(.A1(new_n539), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n587));
  INV_X1    g162(.A(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n534), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n521), .B2(new_n522), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n533), .A2(G86), .A3(new_n523), .ZN(new_n597));
  OAI211_X1 g172(.A(G48), .B(G543), .C1(new_n531), .C2(new_n532), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G305));
  XNOR2_X1  g174(.A(KEYINPUT80), .B(G47), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n534), .A2(new_n600), .B1(new_n601), .B2(new_n538), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n520), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(G301), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n539), .A2(G92), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT10), .Z(new_n610));
  NAND2_X1  g185(.A1(new_n535), .A2(KEYINPUT81), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n534), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n579), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n611), .A2(new_n614), .B1(G651), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(KEYINPUT82), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(KEYINPUT82), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n608), .B1(new_n622), .B2(new_n607), .ZN(G321));
  XNOR2_X1  g198(.A(G321), .B(KEYINPUT83), .ZN(G284));
  NAND2_X1  g199(.A1(G299), .A2(new_n607), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(new_n628), .B2(G860), .ZN(G148));
  NOR2_X1   g204(.A1(new_n567), .A2(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n628), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT84), .Z(G323));
  XNOR2_X1  g208(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n634));
  XNOR2_X1  g209(.A(G323), .B(new_n634), .ZN(G282));
  NAND2_X1  g210(.A1(new_n506), .A2(new_n471), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  INV_X1    g215(.A(G111), .ZN(new_n641));
  AOI22_X1  g216(.A1(new_n640), .A2(KEYINPUT86), .B1(new_n641), .B2(G2105), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(KEYINPUT86), .B2(new_n640), .ZN(new_n643));
  INV_X1    g218(.A(G123), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n490), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(G135), .B2(new_n495), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(G2096), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(G2096), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n639), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT87), .ZN(G156));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT88), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT18), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n667), .A2(new_n668), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n675), .B(new_n679), .Z(G227));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n683), .B2(new_n689), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1981), .B(G1986), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  NAND2_X1  g274(.A1(G166), .A2(G16), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G16), .B2(G22), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  MUX2_X1   g279(.A(G6), .B(G305), .S(G16), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT92), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT32), .B(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n590), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n703), .A2(new_n704), .A3(new_n708), .A4(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n720));
  INV_X1    g295(.A(G119), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n490), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G131), .B2(new_n495), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n718), .B1(new_n723), .B2(new_n717), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT90), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G24), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n605), .B(KEYINPUT91), .Z(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G16), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G1986), .Z(new_n731));
  NAND4_X1  g306(.A1(new_n715), .A2(new_n716), .A3(new_n727), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT36), .ZN(new_n733));
  NOR2_X1   g308(.A1(G5), .A2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT99), .Z(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G171), .B2(G16), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G1961), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT100), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n709), .A2(G19), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT93), .ZN(new_n740));
  INV_X1    g315(.A(new_n567), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT94), .B(G1341), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT26), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n747), .A2(new_n748), .B1(new_n471), .B2(G105), .ZN(new_n749));
  INV_X1    g324(.A(G129), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n490), .B2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G141), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n467), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT97), .ZN(new_n754));
  OR3_X1    g329(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n751), .B2(new_n753), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G32), .B(new_n757), .S(G29), .Z(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n744), .B(new_n761), .C1(new_n742), .C2(new_n743), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n717), .A2(G33), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT25), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n495), .A2(G139), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n506), .A2(G127), .ZN(new_n767));
  INV_X1    g342(.A(G115), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n460), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n765), .B(new_n766), .C1(G2105), .C2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n763), .B1(new_n770), .B2(new_n717), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2072), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n709), .A2(G20), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT23), .Z(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G299), .B2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n709), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n709), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n717), .A2(G27), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G164), .B2(new_n717), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT101), .B(G2078), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G28), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT30), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n787), .B2(KEYINPUT30), .ZN(new_n789));
  OR2_X1    g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  NAND2_X1  g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n788), .A2(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n792), .B1(new_n647), .B2(new_n717), .C1(G1961), .C2(new_n736), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n780), .B2(G1966), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n778), .A2(new_n782), .A3(new_n786), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n758), .A2(new_n760), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n717), .B1(KEYINPUT24), .B2(G34), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(KEYINPUT24), .B2(G34), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n488), .B2(G29), .ZN(new_n799));
  INV_X1    g374(.A(G2084), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n762), .A2(new_n795), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n709), .A2(G4), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n622), .B2(new_n709), .ZN(new_n804));
  INV_X1    g379(.A(G1348), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G29), .A2(G35), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G162), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT29), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(G2090), .Z(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n717), .A2(G26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(G104), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n815));
  INV_X1    g390(.A(G140), .ZN(new_n816));
  INV_X1    g391(.A(G128), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n815), .B1(new_n467), .B2(new_n816), .C1(new_n817), .C2(new_n490), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT95), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(G29), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2067), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n802), .A2(new_n806), .A3(new_n810), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT102), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n733), .A2(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  INV_X1    g400(.A(G55), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n534), .A2(new_n826), .B1(new_n827), .B2(new_n538), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n520), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT103), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(KEYINPUT103), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n741), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n567), .A2(KEYINPUT103), .A3(new_n831), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n622), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n840));
  AOI21_X1  g415(.A(G860), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT104), .Z(new_n843));
  INV_X1    g418(.A(new_n831), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(G145));
  XNOR2_X1  g422(.A(new_n819), .B(new_n770), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n500), .A2(G130), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n465), .A2(G118), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G142), .B2(new_n495), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n637), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n848), .B(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n512), .A2(new_n516), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n757), .B(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(new_n723), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n855), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n488), .B(new_n647), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G162), .ZN(new_n861));
  AOI21_X1  g436(.A(G37), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n859), .A2(KEYINPUT105), .A3(new_n861), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n857), .B(new_n723), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n855), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n861), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n862), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT106), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g446(.A(KEYINPUT106), .B(new_n862), .C1(new_n863), .C2(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(G395));
  NAND2_X1  g450(.A1(new_n844), .A2(new_n607), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n590), .B(KEYINPUT110), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G303), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n605), .B(G305), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n631), .B(new_n836), .ZN(new_n882));
  INV_X1    g457(.A(G299), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n619), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT108), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(G299), .A2(new_n610), .A3(new_n618), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n884), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n894), .A2(new_n890), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n889), .B1(new_n896), .B2(new_n882), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n881), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n876), .B1(new_n898), .B2(new_n607), .ZN(G295));
  OAI21_X1  g474(.A(new_n876), .B1(new_n898), .B2(new_n607), .ZN(G331));
  XNOR2_X1  g475(.A(G168), .B(G171), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n836), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n836), .A2(new_n901), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n888), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n894), .A2(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n888), .A2(KEYINPUT41), .ZN(new_n908));
  OAI211_X1 g483(.A(KEYINPUT111), .B(new_n904), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n880), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n909), .B(new_n910), .C1(KEYINPUT111), .C2(new_n904), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n905), .B1(new_n891), .B2(new_n895), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n880), .A3(new_n904), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n913), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n880), .B1(new_n914), .B2(new_n904), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n911), .A2(KEYINPUT43), .A3(new_n913), .A4(new_n915), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  MUX2_X1   g498(.A(new_n920), .B(new_n923), .S(KEYINPUT44), .Z(G397));
  INV_X1    g499(.A(G2067), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n819), .B(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G1996), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n757), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n723), .B(new_n726), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(G290), .A2(G1986), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G290), .A2(G1986), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n512), .B2(new_n516), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n483), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n940));
  OAI21_X1  g515(.A(G40), .B1(new_n940), .B2(new_n484), .ZN(new_n941));
  NOR4_X1   g516(.A1(new_n473), .A2(new_n939), .A3(new_n476), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n935), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G8), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n510), .B1(new_n501), .B2(new_n509), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n512), .A2(new_n516), .A3(KEYINPUT73), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n936), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT50), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n473), .A2(new_n476), .A3(new_n941), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n951), .B(new_n936), .C1(new_n512), .C2(new_n516), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n949), .A2(new_n950), .A3(new_n800), .A4(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1966), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n464), .B1(new_n495), .B2(G137), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n467), .A2(KEYINPUT71), .A3(new_n468), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n472), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n474), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n470), .A2(KEYINPUT72), .A3(new_n472), .ZN(new_n959));
  INV_X1    g534(.A(G40), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n485), .B2(new_n486), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n961), .A4(new_n939), .ZN(new_n962));
  AOI211_X1 g537(.A(new_n938), .B(G1384), .C1(new_n511), .C2(new_n517), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n945), .B1(new_n953), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n965), .A2(G168), .ZN(new_n966));
  INV_X1    g541(.A(new_n937), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n958), .A2(new_n959), .A3(new_n961), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n590), .A2(G1976), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(G8), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n590), .B2(G1976), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G86), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n598), .B1(new_n538), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(G61), .B1(new_n536), .B2(new_n537), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n520), .B1(new_n978), .B2(new_n594), .ZN(new_n979));
  OAI21_X1  g554(.A(G1981), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1981), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n596), .A2(new_n597), .A3(new_n981), .A4(new_n598), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n980), .A2(KEYINPUT49), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT49), .B1(new_n980), .B2(new_n982), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n968), .A2(G8), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n968), .A2(KEYINPUT115), .A3(new_n985), .A4(G8), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n966), .A2(new_n975), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(G8), .B1(new_n530), .B2(new_n541), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT55), .B(G8), .C1(new_n530), .C2(new_n541), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT112), .B(G1971), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT45), .B(new_n936), .C1(new_n512), .C2(new_n516), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n958), .A2(new_n959), .A3(new_n961), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT45), .B1(new_n518), .B2(new_n936), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND4_X1   g577(.A1(new_n958), .A2(new_n959), .A3(new_n961), .A4(new_n952), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n949), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT113), .B(G2090), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1002), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n996), .B1(new_n1007), .B2(G8), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT63), .B1(new_n991), .B2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g584(.A(G1976), .B(G288), .C1(new_n988), .C2(new_n989), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n982), .B(KEYINPUT116), .Z(new_n1011));
  OAI211_X1 g586(.A(G8), .B(new_n968), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n518), .A2(new_n951), .A3(new_n936), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n937), .A2(KEYINPUT50), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n950), .A2(new_n1005), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1002), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n996), .B1(new_n1016), .B2(G8), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(KEYINPUT63), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1002), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n958), .A2(new_n959), .A3(new_n961), .A4(new_n952), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n951), .B1(new_n518), .B2(new_n936), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n1006), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n996), .B(G8), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT114), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1007), .A2(new_n1025), .A3(G8), .A4(new_n996), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1018), .A2(new_n966), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n990), .A2(new_n973), .A3(new_n974), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1009), .B(new_n1012), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1032));
  INV_X1    g607(.A(G2078), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1961), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(KEYINPUT53), .ZN(new_n1037));
  AOI211_X1 g612(.A(new_n960), .B(new_n1037), .C1(new_n483), .C2(G2105), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n939), .A2(new_n999), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT123), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT123), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n473), .B2(new_n476), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1030), .B1(new_n1034), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n948), .A2(new_n938), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(new_n950), .A3(new_n1033), .A4(new_n999), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1031), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1049), .A2(KEYINPUT124), .A3(new_n1036), .A4(new_n1043), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1045), .A2(new_n1050), .A3(G171), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n518), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1037), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n950), .A2(new_n1052), .A3(new_n939), .A4(new_n1053), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1036), .A2(new_n1054), .A3(KEYINPUT121), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT121), .B1(new_n1036), .B2(new_n1054), .ZN(new_n1056));
  OAI211_X1 g631(.A(G301), .B(new_n1049), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(KEYINPUT54), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n953), .A2(new_n964), .A3(G168), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n945), .B1(KEYINPUT120), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1060), .A2(KEYINPUT120), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n965), .A2(G286), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1063), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1059), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1028), .A2(new_n1017), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1058), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1961), .B1(new_n1003), .B2(new_n949), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n962), .A2(new_n963), .A3(new_n1037), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1036), .A2(new_n1054), .A3(KEYINPUT121), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1049), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G171), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1049), .A2(new_n1036), .A3(new_n1043), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(G171), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT54), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1071), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT56), .B(G2072), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1046), .A2(new_n950), .A3(new_n999), .A4(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n958), .A2(new_n959), .A3(new_n961), .A4(new_n1014), .ZN(new_n1088));
  AOI211_X1 g663(.A(KEYINPUT50), .B(G1384), .C1(new_n511), .C2(new_n517), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n776), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n577), .B2(new_n582), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1087), .A2(new_n1090), .A3(KEYINPUT118), .A4(new_n1095), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(KEYINPUT61), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1087), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1085), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n741), .A2(KEYINPUT117), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1000), .A2(new_n1001), .A3(G1996), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT58), .B(G1341), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n950), .B2(new_n967), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1107), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT59), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n1107), .C1(new_n1108), .C2(new_n1110), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1105), .A2(new_n1106), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1004), .A2(new_n805), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n950), .A2(new_n925), .A3(new_n967), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1116), .B(new_n1117), .C1(new_n622), .C2(KEYINPUT60), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n622), .A2(KEYINPUT60), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1116), .A2(new_n622), .A3(KEYINPUT60), .A4(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1095), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(new_n1106), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(new_n1102), .A3(KEYINPUT119), .A4(new_n1098), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1104), .A2(new_n1115), .A3(new_n1122), .A4(new_n1125), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1116), .A2(new_n1117), .B1(new_n621), .B2(new_n620), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1100), .B1(new_n1127), .B2(new_n1123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1029), .B1(new_n1084), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(G301), .B1(new_n1077), .B2(new_n1049), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1131), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1064), .A2(new_n1133), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(KEYINPUT125), .A3(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n1069), .A3(new_n1070), .A4(new_n1131), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1067), .A2(new_n1065), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1066), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT62), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1068), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1135), .A2(new_n1138), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n944), .B1(new_n1130), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n942), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n931), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n933), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(KEYINPUT48), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(KEYINPUT48), .B2(new_n1149), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n942), .A2(new_n927), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT46), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n926), .A2(new_n756), .A3(new_n755), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1147), .B2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT47), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n723), .A2(new_n726), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n929), .A2(new_n1157), .B1(G2067), .B2(new_n819), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n942), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1151), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT127), .B1(new_n1146), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n965), .A2(G168), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1008), .A2(new_n1028), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1012), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n1131), .B2(new_n1081), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1169), .A2(new_n1171), .A3(new_n1068), .A4(new_n1058), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1167), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1143), .B(new_n1144), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT125), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n943), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1160), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1161), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g756(.A(G319), .ZN(new_n1183));
  OR4_X1    g757(.A1(new_n1183), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1184));
  AOI21_X1  g758(.A(new_n1184), .B1(new_n916), .B2(new_n919), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n1185), .A2(new_n873), .ZN(G225));
  INV_X1    g760(.A(G225), .ZN(G308));
endmodule


