//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT2), .A2(G113), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT65), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT2), .A3(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT2), .A2(G113), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n196), .A2(KEYINPUT66), .A3(G119), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT66), .B1(new_n196), .B2(G119), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G116), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n196), .A2(KEYINPUT66), .A3(G119), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n197), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n193), .B1(new_n189), .B2(new_n191), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n212));
  OR2_X1    g026(.A1(KEYINPUT78), .A2(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT78), .A2(G107), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n210), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n202), .A2(new_n209), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT86), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n225));
  AOI21_X1  g039(.A(G107), .B1(new_n211), .B2(KEYINPUT3), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(new_n212), .ZN(new_n227));
  OAI21_X1  g041(.A(G101), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT79), .A2(G101), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT79), .A2(G101), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n215), .A2(new_n220), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(KEYINPUT4), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n223), .A2(new_n224), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n210), .B1(G104), .B2(G107), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n213), .A2(new_n214), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G104), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT83), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n207), .A2(KEYINPUT5), .ZN(new_n241));
  INV_X1    g055(.A(G113), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(new_n197), .B2(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n241), .A2(new_n244), .B1(new_n208), .B2(new_n207), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n232), .A2(KEYINPUT83), .A3(new_n237), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n234), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n224), .B1(new_n223), .B2(new_n233), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT87), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n222), .B(G101), .C1(new_n225), .C2(new_n227), .ZN(new_n251));
  INV_X1    g065(.A(new_n209), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n207), .A2(new_n208), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n232), .A2(KEYINPUT4), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(new_n221), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT86), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT87), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n258), .A3(new_n247), .A4(new_n234), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G122), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n250), .A2(KEYINPUT6), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n234), .A2(new_n247), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT88), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n257), .A4(new_n260), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n257), .A2(new_n247), .A3(new_n234), .A4(new_n260), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT88), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n263), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n250), .A2(new_n259), .A3(new_n261), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n262), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT89), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  OR2_X1    g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(G146), .ZN(new_n276));
  INV_X1    g090(.A(G146), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G143), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n273), .B(new_n274), .C1(new_n276), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(G146), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT0), .A4(G128), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G125), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n272), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G128), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(KEYINPUT1), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n287), .A2(new_n280), .A3(new_n281), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n280), .A2(new_n281), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(KEYINPUT64), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT64), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G128), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT1), .B1(new_n275), .B2(G146), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n288), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n284), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n285), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n279), .A2(new_n282), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(KEYINPUT89), .A3(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT90), .B(G224), .Z(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(G953), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n301), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n271), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n304), .A2(KEYINPUT7), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n285), .A2(new_n308), .A3(new_n300), .A4(new_n297), .ZN(new_n309));
  XOR2_X1   g123(.A(new_n309), .B(KEYINPUT93), .Z(new_n310));
  AND2_X1   g124(.A1(new_n232), .A2(new_n237), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n241), .A2(KEYINPUT91), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n244), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n241), .A2(KEYINPUT91), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n209), .B(new_n311), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT92), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n245), .B2(new_n311), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n241), .A2(new_n244), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT92), .B(new_n238), .C1(new_n318), .C2(new_n252), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n260), .B(KEYINPUT8), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n308), .B1(new_n298), .B2(new_n300), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n310), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n266), .A2(new_n268), .ZN(new_n325));
  AOI21_X1  g139(.A(G902), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G210), .B1(G237), .B2(G902), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n307), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n307), .B2(new_n326), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n187), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT9), .B(G234), .ZN(new_n331));
  OAI21_X1  g145(.A(G221), .B1(new_n331), .B2(G902), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT11), .ZN(new_n333));
  INV_X1    g147(.A(G134), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(G137), .ZN(new_n335));
  INV_X1    g149(.A(G137), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT11), .A3(G134), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(G137), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G131), .ZN(new_n340));
  AOI21_X1  g154(.A(G131), .B1(new_n334), .B2(G137), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(new_n341), .A3(new_n337), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n246), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT83), .B1(new_n232), .B2(new_n237), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n296), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n299), .B1(new_n222), .B2(new_n221), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n346), .A2(new_n348), .B1(new_n233), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n294), .A2(KEYINPUT80), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n280), .A2(new_n352), .A3(KEYINPUT1), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(G128), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n289), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n287), .A2(new_n280), .A3(new_n281), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(new_n311), .A3(KEYINPUT81), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n288), .B1(new_n354), .B2(new_n289), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(new_n238), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT10), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n350), .B1(new_n362), .B2(KEYINPUT82), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT81), .B1(new_n357), .B2(new_n311), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n360), .A2(new_n238), .A3(new_n359), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n347), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n343), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n362), .A2(KEYINPUT82), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n335), .A2(new_n337), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n372), .A2(new_n341), .B1(new_n339), .B2(G131), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n370), .A2(new_n371), .A3(new_n373), .A4(new_n350), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT71), .B(G953), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G227), .ZN(new_n377));
  XOR2_X1   g191(.A(G110), .B(G140), .Z(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT12), .B1(new_n343), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT64), .B(G128), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT1), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(G143), .B2(new_n277), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n289), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n356), .ZN(new_n388));
  OAI22_X1  g202(.A1(new_n364), .A2(new_n365), .B1(new_n388), .B2(new_n311), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n383), .B1(new_n389), .B2(new_n343), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n358), .A2(new_n361), .B1(new_n296), .B2(new_n238), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n391), .A2(new_n373), .A3(new_n382), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT85), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n382), .B1(new_n391), .B2(new_n373), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n343), .A3(new_n383), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n379), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n397), .A3(new_n374), .A4(new_n398), .ZN(new_n399));
  AOI211_X1 g213(.A(G469), .B(G902), .C1(new_n380), .C2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n374), .B1(new_n392), .B2(new_n390), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n379), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n369), .A2(new_n374), .A3(new_n398), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(G469), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(G469), .A2(G902), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n332), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT20), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT70), .B(G237), .Z(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(G214), .A3(new_n376), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n275), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n409), .A2(G143), .A3(G214), .A4(new_n376), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G131), .ZN(new_n414));
  INV_X1    g228(.A(G131), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G140), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G125), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT16), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n284), .A2(G140), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT76), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n418), .B2(G125), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n284), .A2(KEYINPUT76), .A3(G140), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n421), .B1(new_n426), .B2(new_n420), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G146), .ZN(new_n428));
  INV_X1    g242(.A(new_n426), .ZN(new_n429));
  XNOR2_X1  g243(.A(G125), .B(G140), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n431));
  AOI22_X1  g245(.A1(new_n429), .A2(KEYINPUT19), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT95), .A3(new_n277), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n430), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n434), .B(new_n277), .C1(new_n435), .C2(new_n426), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT95), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n417), .A2(new_n428), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n413), .A2(KEYINPUT18), .A3(G131), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n430), .A2(new_n277), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n426), .B2(new_n277), .ZN(new_n443));
  NAND2_X1  g257(.A1(KEYINPUT18), .A2(G131), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n411), .A2(new_n412), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G113), .B(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n211), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n277), .B(new_n421), .C1(new_n426), .C2(new_n420), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n428), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n415), .B1(new_n411), .B2(new_n412), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(KEYINPUT17), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n414), .A2(new_n456), .A3(new_n416), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n449), .A3(new_n446), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(G475), .A2(G902), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n408), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  AOI211_X1 g277(.A(KEYINPUT20), .B(new_n463), .C1(new_n451), .C2(new_n459), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n446), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n450), .ZN(new_n466));
  AOI21_X1  g280(.A(G902), .B1(new_n466), .B2(new_n459), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT96), .B(G475), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI22_X1  g283(.A1(new_n462), .A2(new_n464), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G217), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n331), .A2(new_n471), .A3(G953), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT97), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT78), .B(G107), .Z(new_n475));
  XNOR2_X1  g289(.A(G116), .B(G122), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G116), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n196), .A2(G122), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n236), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n474), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n290), .A2(new_n292), .A3(G143), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n485));
  OAI221_X1 g299(.A(new_n484), .B1(new_n286), .B2(G143), .C1(new_n334), .C2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n334), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n484), .B1(new_n286), .B2(G143), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n475), .A2(new_n476), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n236), .A2(new_n481), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT97), .A3(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n483), .A2(new_n486), .A3(new_n489), .A4(new_n492), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n481), .A2(KEYINPUT14), .ZN(new_n494));
  INV_X1    g308(.A(new_n480), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n216), .B1(new_n495), .B2(KEYINPUT14), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n482), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT99), .B(G134), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n488), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n498), .B(new_n484), .C1(new_n286), .C2(G143), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT100), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n503), .B1(new_n493), .B2(new_n502), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n473), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G902), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n493), .A2(new_n502), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT100), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n472), .A3(new_n504), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G478), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n512), .B(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n470), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G952), .ZN(new_n517));
  AOI211_X1 g331(.A(G953), .B(new_n517), .C1(G234), .C2(G237), .ZN(new_n518));
  AOI211_X1 g332(.A(new_n508), .B(new_n376), .C1(G234), .C2(G237), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT21), .B(G898), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n330), .A2(new_n407), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n471), .B1(G234), .B2(new_n508), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n376), .A2(G221), .A3(G234), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT22), .B(G137), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT23), .B1(new_n286), .B2(G119), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n286), .A2(G119), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n290), .A2(new_n292), .A3(G119), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n530), .B1(new_n384), .B2(G119), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT24), .B(G110), .Z(new_n536));
  AOI22_X1  g350(.A1(new_n534), .A2(G110), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n442), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n427), .B2(G146), .ZN(new_n539));
  OAI22_X1  g353(.A1(new_n534), .A2(G110), .B1(new_n535), .B2(new_n536), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n453), .A2(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n528), .B1(new_n541), .B2(KEYINPUT77), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT77), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(G110), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n535), .A2(new_n536), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n452), .B2(new_n428), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n539), .A2(new_n540), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n541), .A2(KEYINPUT77), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n542), .B1(new_n551), .B2(new_n528), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT25), .B1(new_n552), .B2(new_n508), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n453), .A2(new_n537), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n539), .A2(new_n540), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n554), .A2(KEYINPUT77), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT77), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n528), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n542), .ZN(new_n559));
  AND4_X1   g373(.A1(KEYINPUT25), .A2(new_n558), .A3(new_n508), .A4(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n525), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n525), .A2(G902), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n552), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n409), .A2(G210), .A3(new_n376), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT27), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT27), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n409), .A2(new_n569), .A3(G210), .A4(new_n376), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT26), .B(G101), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT67), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n373), .B2(new_n299), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n335), .A2(new_n341), .A3(new_n337), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n336), .A2(G134), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n415), .B1(new_n580), .B2(new_n338), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT68), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT68), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n342), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n585), .A3(new_n388), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n283), .A2(new_n343), .A3(KEYINPUT67), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n578), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT69), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n202), .A2(new_n589), .A3(new_n209), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n202), .B2(new_n209), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n576), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n578), .A2(new_n586), .A3(new_n587), .A4(KEYINPUT30), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n202), .A2(new_n209), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n583), .A2(new_n342), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n596), .A2(new_n296), .B1(new_n373), .B2(new_n299), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT30), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n566), .B1(new_n593), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n597), .A2(new_n595), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n578), .A2(new_n586), .A3(new_n587), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT69), .B1(new_n252), .B2(new_n253), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n202), .A2(new_n589), .A3(new_n209), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n602), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT28), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n283), .A2(new_n343), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n604), .A2(new_n586), .A3(new_n609), .A4(new_n605), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT73), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT28), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT73), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n608), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n601), .B1(new_n616), .B2(new_n576), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n592), .A2(new_n587), .A3(new_n586), .A4(new_n578), .ZN(new_n618));
  INV_X1    g432(.A(new_n576), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n600), .A2(new_n618), .A3(new_n566), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT72), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT72), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n593), .A2(new_n622), .A3(new_n566), .A4(new_n600), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n617), .A2(KEYINPUT74), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT74), .B1(new_n617), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n565), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT32), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT32), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n629), .B(new_n565), .C1(new_n625), .C2(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n603), .A2(new_n606), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n618), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT28), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n615), .A2(KEYINPUT75), .A3(new_n613), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT75), .B1(new_n615), .B2(new_n613), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT29), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n637), .A2(new_n638), .A3(new_n576), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n600), .A2(new_n618), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n619), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n616), .B2(new_n619), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n508), .B1(new_n642), .B2(KEYINPUT29), .ZN(new_n643));
  OAI21_X1  g457(.A(G472), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n564), .B1(new_n631), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n524), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(new_n231), .Z(G3));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n307), .A2(new_n648), .A3(new_n326), .A4(new_n327), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n187), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n328), .A2(new_n329), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n651), .B2(KEYINPUT101), .ZN(new_n652));
  INV_X1    g466(.A(new_n459), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n449), .B1(new_n440), .B2(new_n446), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n461), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT20), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n460), .A2(new_n408), .A3(new_n461), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n466), .A2(new_n459), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n508), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n656), .A2(new_n657), .B1(new_n659), .B2(new_n468), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n512), .A2(new_n513), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n512), .A2(KEYINPUT103), .A3(new_n513), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT33), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n665), .A2(KEYINPUT33), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n505), .A2(new_n473), .A3(new_n506), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n472), .B1(new_n510), .B2(new_n504), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n666), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n507), .A2(new_n511), .A3(new_n665), .A4(KEYINPUT33), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n513), .A2(G902), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n663), .A2(new_n664), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n660), .A2(new_n674), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n652), .A2(new_n522), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n508), .B1(new_n625), .B2(new_n626), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n617), .A2(new_n624), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT74), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n617), .A2(new_n624), .A3(KEYINPUT74), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n677), .A2(G472), .B1(new_n682), .B2(new_n565), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n561), .A2(new_n563), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n684), .B(new_n332), .C1(new_n400), .C2(new_n406), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n676), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT104), .Z(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT34), .B(G104), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G6));
  NAND2_X1  g504(.A1(new_n660), .A2(new_n515), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n652), .A2(new_n522), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n683), .A3(new_n686), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT35), .B(G107), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  INV_X1    g510(.A(new_n683), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n697), .A2(new_n330), .A3(new_n407), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  INV_X1    g513(.A(new_n525), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n552), .A2(KEYINPUT25), .A3(new_n508), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n558), .A2(new_n508), .A3(new_n559), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT25), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n700), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n528), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(KEYINPUT36), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n541), .B(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n708), .A2(G902), .A3(new_n525), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n699), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n709), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n561), .A2(KEYINPUT105), .A3(new_n711), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n522), .A2(new_n516), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n698), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT37), .B(G110), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G12));
  AOI21_X1  g530(.A(new_n629), .B1(new_n682), .B2(new_n565), .ZN(new_n717));
  INV_X1    g531(.A(new_n630), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n644), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n710), .A2(new_n712), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n407), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(G900), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n519), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n518), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n691), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n652), .A2(new_n719), .A3(new_n721), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G128), .ZN(G30));
  INV_X1    g541(.A(new_n262), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n267), .A2(KEYINPUT88), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n267), .A2(KEYINPUT88), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT6), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n250), .A2(new_n259), .A3(new_n261), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n326), .B1(new_n733), .B2(new_n305), .ZN(new_n734));
  INV_X1    g548(.A(new_n327), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n307), .A2(new_n326), .A3(new_n327), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT38), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n701), .A2(new_n704), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n709), .B1(new_n740), .B2(new_n525), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n470), .A2(new_n515), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n739), .A2(new_n187), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n332), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n374), .A2(new_n398), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n745), .A2(new_n369), .B1(new_n401), .B2(new_n379), .ZN(new_n746));
  OAI21_X1  g560(.A(G469), .B1(new_n746), .B2(G902), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n380), .A2(new_n399), .ZN(new_n748));
  INV_X1    g562(.A(G469), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n508), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n744), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n724), .B(KEYINPUT39), .Z(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n743), .B1(KEYINPUT40), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n640), .A2(new_n619), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n508), .B1(new_n633), .B2(new_n619), .ZN(new_n757));
  OAI21_X1  g571(.A(G472), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n717), .B2(new_n718), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n758), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n628), .B2(new_n630), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT106), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n754), .B(new_n765), .C1(KEYINPUT40), .C2(new_n753), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G143), .ZN(G45));
  NOR3_X1   g581(.A1(new_n660), .A2(new_n674), .A3(new_n724), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n652), .A2(new_n719), .A3(new_n721), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G146), .ZN(G48));
  NAND2_X1  g584(.A1(new_n719), .A2(new_n684), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n749), .A2(KEYINPUT107), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n398), .B1(new_n369), .B2(new_n374), .ZN(new_n773));
  INV_X1    g587(.A(new_n397), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n396), .B1(new_n394), .B2(new_n395), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n773), .B1(new_n776), .B2(new_n745), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n772), .B1(new_n777), .B2(G902), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n748), .B(new_n508), .C1(KEYINPUT107), .C2(new_n749), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n778), .A2(new_n779), .A3(new_n332), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n676), .ZN(new_n783));
  XNOR2_X1  g597(.A(KEYINPUT41), .B(G113), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G15));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n693), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G116), .ZN(G18));
  NAND4_X1  g601(.A1(new_n652), .A2(new_n719), .A3(new_n713), .A4(new_n780), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G119), .ZN(G21));
  INV_X1    g603(.A(new_n565), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n637), .A2(new_n576), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n601), .B1(new_n621), .B2(new_n623), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n793), .B(new_n564), .C1(new_n677), .C2(G472), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n332), .A2(new_n778), .A3(new_n779), .A4(new_n522), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n652), .A2(new_n794), .A3(new_n795), .A4(new_n742), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G122), .ZN(G24));
  AOI211_X1 g611(.A(new_n793), .B(new_n741), .C1(new_n677), .C2(G472), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n652), .A2(new_n768), .A3(new_n798), .A4(new_n780), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT108), .B(G125), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(G27));
  NAND3_X1  g615(.A1(new_n736), .A2(new_n187), .A3(new_n737), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n407), .ZN(new_n803));
  INV_X1    g617(.A(new_n724), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n675), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n645), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n809));
  NAND2_X1  g623(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n645), .A2(new_n807), .A3(new_n803), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n415), .ZN(G33));
  NAND4_X1  g627(.A1(new_n803), .A2(new_n719), .A3(new_n684), .A4(new_n725), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n645), .A2(KEYINPUT110), .A3(new_n725), .A4(new_n803), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G134), .ZN(G36));
  OR2_X1    g633(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(G469), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT46), .B1(new_n822), .B2(new_n405), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n400), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(KEYINPUT46), .A3(new_n405), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n744), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n752), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT43), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT111), .ZN(new_n829));
  XOR2_X1   g643(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n830));
  INV_X1    g644(.A(new_n674), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n660), .ZN(new_n832));
  MUX2_X1   g646(.A(new_n829), .B(new_n830), .S(new_n832), .Z(new_n833));
  INV_X1    g647(.A(new_n741), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n697), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT44), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT44), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n838), .A3(new_n697), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n802), .B(KEYINPUT112), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n827), .B1(new_n843), .B2(KEYINPUT113), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G137), .ZN(G39));
  XNOR2_X1  g662(.A(new_n826), .B(KEYINPUT47), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n719), .A2(new_n684), .A3(new_n805), .A4(new_n802), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G140), .ZN(G42));
  AND2_X1   g666(.A1(new_n778), .A2(new_n779), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(KEYINPUT49), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(KEYINPUT49), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n684), .A2(new_n187), .A3(new_n332), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n855), .A2(new_n856), .A3(new_n832), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n765), .ZN(new_n859));
  INV_X1    g673(.A(new_n739), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n726), .A2(new_n769), .A3(new_n799), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n736), .A2(KEYINPUT101), .A3(new_n737), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n649), .A2(new_n187), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n742), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n834), .A2(new_n724), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n751), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n763), .A2(KEYINPUT106), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n760), .B(new_n762), .C1(new_n628), .C2(new_n630), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n870), .B1(new_n765), .B2(new_n869), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n863), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT115), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n862), .B1(new_n880), .B2(new_n873), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n751), .A2(new_n651), .A3(new_n187), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n793), .B1(new_n677), .B2(G472), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n834), .A3(new_n768), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n803), .A2(new_n798), .A3(KEYINPUT114), .A4(new_n768), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n516), .A2(new_n710), .A3(new_n712), .A4(new_n804), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n631), .B2(new_n644), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n888), .A2(new_n889), .B1(new_n803), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n818), .A2(new_n892), .A3(new_n809), .A4(new_n811), .ZN(new_n893));
  INV_X1    g707(.A(new_n330), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n831), .A2(new_n470), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n521), .B1(new_n895), .B2(new_n691), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n686), .A2(new_n894), .A3(new_n896), .A4(new_n683), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n788), .A2(new_n796), .A3(new_n897), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n698), .A2(new_n713), .B1(new_n645), .B2(new_n524), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n783), .A3(new_n786), .A4(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n883), .A2(KEYINPUT53), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT117), .ZN(new_n903));
  OAI211_X1 g717(.A(KEYINPUT116), .B(new_n877), .C1(new_n881), .C2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n904), .A2(new_n901), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n877), .B1(new_n876), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT116), .B1(new_n881), .B2(new_n903), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n902), .B1(new_n910), .B2(KEYINPUT53), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n905), .A2(KEYINPUT53), .A3(new_n909), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n915), .B(KEYINPUT53), .C1(new_n883), .C2(new_n901), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n881), .A2(KEYINPUT52), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n877), .B(new_n862), .C1(new_n880), .C2(new_n873), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n901), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT53), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT118), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n913), .B(new_n914), .C1(new_n916), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n912), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n833), .A2(new_n518), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(new_n794), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n739), .A2(new_n781), .A3(new_n187), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT50), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT119), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n781), .A2(new_n802), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n859), .A2(new_n684), .A3(new_n518), .A4(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n660), .A3(new_n674), .ZN(new_n935));
  INV_X1    g749(.A(new_n798), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n925), .A2(new_n932), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n849), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n332), .B2(new_n854), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n926), .A2(new_n841), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT51), .B1(new_n931), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n930), .A3(KEYINPUT51), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n937), .A2(new_n771), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT48), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n934), .A2(new_n675), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n652), .A2(new_n780), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI211_X1 g763(.A(new_n517), .B(G953), .C1(new_n926), .C2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n944), .A2(new_n946), .A3(new_n947), .A4(new_n950), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n923), .A2(new_n943), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(G952), .A2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n861), .B1(new_n952), .B2(new_n953), .ZN(G75));
  NOR2_X1   g768(.A1(new_n376), .A2(G952), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n733), .A2(new_n305), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n307), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT55), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n913), .B1(new_n916), .B2(new_n921), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(G902), .ZN(new_n960));
  AOI211_X1 g774(.A(KEYINPUT56), .B(new_n958), .C1(new_n960), .C2(G210), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(G210), .A3(G902), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT56), .B1(new_n962), .B2(KEYINPUT120), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(KEYINPUT120), .B2(new_n962), .ZN(new_n964));
  AOI211_X1 g778(.A(new_n955), .B(new_n961), .C1(new_n958), .C2(new_n964), .ZN(G51));
  NAND2_X1  g779(.A1(new_n959), .A2(KEYINPUT54), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(KEYINPUT121), .A3(new_n922), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT121), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n959), .A2(new_n968), .A3(KEYINPUT54), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n405), .B(KEYINPUT57), .Z(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n748), .ZN(new_n972));
  INV_X1    g786(.A(new_n822), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n960), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n955), .B1(new_n972), .B2(new_n974), .ZN(G54));
  NAND3_X1  g789(.A1(new_n960), .A2(KEYINPUT58), .A3(G475), .ZN(new_n976));
  INV_X1    g790(.A(new_n460), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n978), .A2(new_n979), .A3(new_n955), .ZN(G60));
  NAND2_X1  g794(.A1(G478), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT59), .Z(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n670), .B2(new_n671), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n967), .A2(new_n969), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n955), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n984), .A2(KEYINPUT122), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(KEYINPUT122), .B1(new_n984), .B2(new_n985), .ZN(new_n987));
  INV_X1    g801(.A(new_n982), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n672), .B1(new_n923), .B2(new_n988), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(G63));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT60), .Z(new_n992));
  AND2_X1   g806(.A1(new_n959), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n708), .B(KEYINPUT123), .Z(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n995), .B(new_n985), .C1(new_n552), .C2(new_n993), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT61), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G66));
  OAI21_X1  g812(.A(G953), .B1(new_n302), .B2(new_n520), .ZN(new_n999));
  INV_X1    g813(.A(new_n900), .ZN(new_n1000));
  INV_X1    g814(.A(new_n376), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n733), .B1(G898), .B2(new_n376), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(G69));
  AOI21_X1  g818(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n827), .A2(new_n771), .A3(new_n866), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1006), .A2(new_n862), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n847), .A2(new_n851), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1008), .A2(new_n1001), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n594), .A2(new_n599), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(new_n432), .Z(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(new_n722), .B2(new_n376), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT126), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1011), .B(KEYINPUT124), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n766), .A2(new_n863), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT62), .Z(new_n1017));
  AOI211_X1 g831(.A(new_n802), .B(new_n753), .C1(new_n895), .C2(new_n691), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n645), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT125), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1017), .A2(new_n847), .A3(new_n851), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1015), .B1(new_n1021), .B2(new_n376), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n376), .B1(G227), .B2(G900), .ZN(new_n1023));
  OR3_X1    g837(.A1(new_n1013), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1023), .B1(new_n1013), .B2(new_n1022), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(G72));
  XNOR2_X1  g840(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1029), .B1(new_n1008), .B2(new_n900), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n955), .B1(new_n1030), .B2(new_n641), .ZN(new_n1031));
  INV_X1    g845(.A(new_n641), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n911), .A2(new_n1032), .A3(new_n755), .A4(new_n1029), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1029), .B1(new_n1021), .B2(new_n900), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n756), .ZN(new_n1035));
  AND3_X1   g849(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(G57));
endmodule


