//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT1), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n224), .A2(new_n209), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n218), .C1(new_n219), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n219), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT64), .Z(new_n228));
  NOR2_X1   g0028(.A1(new_n226), .A2(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  XNOR2_X1  g0045(.A(KEYINPUT8), .B(G58), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n207), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G150), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n207), .A2(new_n249), .ZN(new_n250));
  OAI22_X1  g0050(.A1(new_n246), .A2(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n251), .B1(G20), .B2(new_n203), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n216), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G13), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n257), .A2(new_n207), .A3(G1), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n254), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n206), .A2(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G50), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n257), .A2(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n261), .B1(G50), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT9), .ZN(new_n266));
  OR3_X1    g0066(.A1(new_n256), .A2(KEYINPUT9), .A3(new_n264), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(KEYINPUT67), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G222), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G77), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(G223), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n271), .B1(new_n272), .B2(new_n269), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(new_n277), .A3(G274), .ZN(new_n283));
  INV_X1    g0083(.A(G226), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G200), .ZN(new_n289));
  OR3_X1    g0089(.A1(new_n288), .A2(KEYINPUT69), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n268), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT69), .B1(new_n288), .B2(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(G190), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT68), .B(KEYINPUT10), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT67), .B1(new_n266), .B2(new_n267), .ZN(new_n296));
  OR3_X1    g0096(.A1(new_n291), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n266), .A2(new_n267), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n293), .C1(new_n289), .C2(new_n288), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G20), .A2(G77), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT15), .B(G87), .Z(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n302), .B1(new_n250), .B2(new_n246), .C1(new_n304), .C2(new_n247), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT66), .ZN(new_n307));
  NOR4_X1   g0107(.A1(new_n307), .A2(new_n257), .A3(new_n207), .A4(G1), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n305), .A2(new_n254), .B1(new_n272), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n254), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(G77), .A3(new_n260), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G238), .ZN(new_n314));
  INV_X1    g0114(.A(G107), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n273), .A2(new_n314), .B1(new_n315), .B2(new_n269), .ZN(new_n316));
  INV_X1    g0116(.A(new_n269), .ZN(new_n317));
  INV_X1    g0117(.A(G232), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n317), .A2(new_n318), .A3(G1698), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n278), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n283), .ZN(new_n321));
  INV_X1    g0121(.A(new_n286), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(G244), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n313), .B1(G190), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n289), .B2(new_n325), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n313), .B(new_n329), .C1(G179), .C2(new_n324), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n265), .B1(new_n288), .B2(G169), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n279), .A2(G179), .A3(new_n287), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n301), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT72), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G33), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n338), .A2(new_n340), .A3(G226), .A4(new_n270), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT70), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n269), .A2(KEYINPUT70), .A3(G226), .A4(new_n270), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n338), .A2(new_n340), .A3(G232), .A4(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n277), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n277), .A2(G238), .A3(new_n285), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT71), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n283), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n352), .B1(new_n283), .B2(new_n351), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT13), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n283), .A2(new_n351), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT71), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n283), .A2(new_n351), .A3(new_n352), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT13), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n348), .B1(new_n343), .B2(new_n344), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(new_n361), .C1(new_n362), .C2(new_n277), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT14), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(G169), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n356), .A2(new_n363), .A3(G179), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n365), .B1(new_n364), .B2(G169), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n337), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(G169), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n372), .A2(KEYINPUT72), .A3(new_n367), .A4(new_n366), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G68), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G20), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n376), .B1(new_n247), .B2(new_n272), .C1(new_n202), .C2(new_n250), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n254), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT11), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n311), .A2(G68), .A3(new_n260), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n262), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n382), .A2(KEYINPUT12), .A3(new_n376), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n309), .A2(new_n375), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(KEYINPUT12), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n374), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G190), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n386), .B1(new_n389), .B2(new_n364), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n289), .B1(new_n356), .B2(new_n363), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G159), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n250), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G58), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n375), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n398), .A2(new_n201), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n396), .B1(new_n399), .B2(G20), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n339), .A2(KEYINPUT73), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT73), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT3), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n403), .A3(G33), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n338), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n207), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n405), .B2(new_n207), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT16), .B(new_n400), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n406), .A2(G20), .ZN(new_n412));
  AOI21_X1  g0212(.A(G33), .B1(new_n401), .B2(new_n403), .ZN(new_n413));
  INV_X1    g0213(.A(new_n340), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n406), .B1(new_n269), .B2(G20), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n375), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n400), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n411), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n410), .A2(new_n419), .A3(new_n254), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n246), .B1(new_n206), .B2(G20), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n259), .B1(new_n258), .B2(new_n246), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT74), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT74), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n420), .A2(new_n425), .A3(new_n422), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G223), .A2(G1698), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n284), .B2(G1698), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(new_n404), .A3(new_n338), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n278), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT75), .B1(new_n286), .B2(new_n318), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT75), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n277), .A2(new_n285), .A3(new_n434), .A4(G232), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n321), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G169), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n432), .A2(new_n436), .A3(G179), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n424), .A2(new_n426), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n424), .A2(KEYINPUT18), .A3(new_n426), .A4(new_n440), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(KEYINPUT76), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n437), .A2(new_n389), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n289), .B1(new_n432), .B2(new_n436), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(new_n420), .A3(new_n422), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT17), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT76), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n441), .A2(new_n451), .A3(new_n442), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n336), .A2(new_n394), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT77), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(G41), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n280), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n281), .A2(G1), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G264), .A3(new_n277), .ZN(new_n461));
  INV_X1    g0261(.A(G294), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n249), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n338), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(G33), .ZN(new_n466));
  MUX2_X1   g0266(.A(G250), .B(G257), .S(G1698), .Z(new_n467));
  AOI21_X1  g0267(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n461), .B1(new_n468), .B2(new_n277), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n277), .A2(G274), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(G169), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT84), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n467), .A2(new_n404), .A3(new_n338), .ZN(new_n476));
  INV_X1    g0276(.A(new_n463), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n277), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n461), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(KEYINPUT84), .B(new_n461), .C1(new_n468), .C2(new_n277), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n472), .ZN(new_n482));
  INV_X1    g0282(.A(G179), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n474), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT23), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n207), .B2(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n315), .A2(KEYINPUT23), .A3(G20), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n249), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n207), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n269), .A2(new_n207), .A3(G87), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G87), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n404), .A2(new_n207), .A3(new_n338), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n485), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n493), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n494), .ZN(new_n502));
  AND4_X1   g0302(.A1(new_n485), .A2(new_n501), .A3(new_n502), .A4(new_n499), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n254), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n259), .B1(G1), .B2(new_n249), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT25), .ZN(new_n507));
  AOI21_X1  g0307(.A(G107), .B1(new_n507), .B2(KEYINPUT83), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT83), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n258), .A2(new_n508), .B1(new_n509), .B2(KEYINPUT25), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n258), .A2(new_n509), .A3(KEYINPUT25), .A4(new_n315), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n506), .A2(G107), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n484), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n514), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n289), .ZN(new_n517));
  OR3_X1    g0317(.A1(new_n469), .A2(G190), .A3(new_n473), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT85), .B1(new_n482), .B2(new_n289), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT86), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT86), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n516), .C1(new_n519), .C2(new_n520), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n515), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G97), .A2(G107), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(new_n497), .B1(new_n347), .B2(new_n207), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G97), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n527), .A2(new_n528), .B1(new_n247), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n404), .A2(new_n207), .A3(G68), .A4(new_n338), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT79), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT79), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n254), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n309), .A2(new_n304), .ZN(new_n537));
  MUX2_X1   g0337(.A(G238), .B(G244), .S(G1698), .Z(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(new_n404), .A3(new_n338), .ZN(new_n539));
  INV_X1    g0339(.A(new_n491), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n277), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n471), .A2(new_n459), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n206), .A2(G45), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n543), .A2(G250), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n277), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(G200), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n506), .A2(G87), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n536), .A2(new_n537), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT80), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n255), .B1(new_n532), .B2(KEYINPUT79), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(new_n535), .B1(new_n309), .B2(new_n304), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n553), .A2(KEYINPUT80), .A3(new_n547), .A4(new_n548), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n541), .A2(new_n546), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G190), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n328), .B1(new_n541), .B2(new_n546), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n471), .A2(new_n459), .B1(new_n544), .B2(new_n277), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n491), .B1(new_n466), .B2(new_n538), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n483), .B(new_n559), .C1(new_n560), .C2(new_n277), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n536), .A2(new_n537), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n505), .A2(new_n304), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G270), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n460), .A2(new_n277), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n472), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(G264), .A2(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n404), .A2(new_n338), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT81), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n317), .A2(G303), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n404), .A2(G257), .A3(new_n270), .A4(new_n338), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n404), .A2(KEYINPUT81), .A3(new_n338), .A4(new_n570), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n573), .A2(new_n574), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n569), .B1(new_n577), .B2(new_n278), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n490), .B1(new_n206), .B2(G33), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n255), .B(new_n579), .C1(new_n306), .C2(new_n308), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n263), .A2(new_n307), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n490), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n253), .A2(new_n216), .B1(G20), .B2(new_n490), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G283), .ZN(new_n586));
  INV_X1    g0386(.A(G97), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n586), .B(new_n207), .C1(G33), .C2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n585), .A2(KEYINPUT20), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT20), .B1(new_n585), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(G169), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT82), .B1(new_n578), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n577), .A2(new_n278), .ZN(new_n595));
  INV_X1    g0395(.A(new_n569), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(G190), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n584), .A2(new_n591), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n598), .C1(new_n289), .C2(new_n578), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  OAI211_X1 g0400(.A(KEYINPUT82), .B(new_n600), .C1(new_n578), .C2(new_n592), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n578), .B(G179), .C1(new_n591), .C2(new_n584), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n594), .A2(new_n599), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n460), .A2(G257), .A3(new_n277), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n472), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n338), .A2(new_n340), .A3(G250), .A4(G1698), .ZN(new_n606));
  AND2_X1   g0406(.A1(KEYINPUT4), .A2(G244), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n338), .A2(new_n340), .A3(new_n607), .A4(new_n270), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n608), .A3(new_n586), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT4), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n404), .A2(G244), .A3(new_n270), .A4(new_n338), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n605), .B1(new_n612), .B2(new_n277), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n315), .B1(new_n415), .B2(new_n416), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT6), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n615), .A2(new_n587), .A3(G107), .ZN(new_n616));
  XNOR2_X1  g0416(.A(G97), .B(G107), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n618), .A2(new_n207), .B1(new_n272), .B2(new_n250), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n254), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n263), .A2(G97), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n506), .B2(G97), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n328), .A2(new_n613), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT78), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n472), .A2(new_n604), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n611), .A2(new_n610), .ZN(new_n626));
  INV_X1    g0426(.A(new_n609), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n625), .B1(new_n628), .B2(new_n278), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n624), .B1(new_n629), .B2(new_n483), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n483), .B(new_n605), .C1(new_n612), .C2(new_n277), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(KEYINPUT78), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n623), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(G190), .B(new_n605), .C1(new_n612), .C2(new_n277), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n634), .A2(new_n620), .A3(new_n622), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n613), .A2(G200), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n566), .A2(new_n603), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n454), .A2(new_n525), .A3(new_n639), .ZN(G372));
  INV_X1    g0440(.A(KEYINPUT87), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n392), .A2(new_n330), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n388), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n386), .B1(new_n370), .B2(new_n373), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT87), .B1(new_n645), .B2(new_n642), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n646), .A3(new_n450), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n420), .A2(new_n422), .B1(new_n439), .B2(new_n438), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n301), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT88), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(new_n335), .ZN(new_n653));
  INV_X1    g0453(.A(new_n301), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n647), .B2(new_n649), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT88), .B1(new_n655), .B2(new_n334), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n629), .A2(new_n624), .A3(new_n483), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n631), .A2(KEYINPUT78), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n623), .B1(new_n635), .B2(new_n636), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n553), .A2(new_n547), .A3(new_n548), .A4(new_n556), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n565), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n594), .A2(new_n602), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n484), .A2(new_n514), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n601), .ZN(new_n667));
  INV_X1    g0467(.A(new_n524), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n482), .A2(new_n289), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT85), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n518), .A3(new_n517), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n523), .B1(new_n672), .B2(new_n516), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n664), .B(new_n667), .C1(new_n668), .C2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n565), .A2(new_n660), .A3(new_n662), .A4(new_n623), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n565), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n676));
  INV_X1    g0476(.A(new_n633), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n557), .A3(new_n565), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(KEYINPUT26), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n454), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n657), .A2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n522), .A2(new_n524), .ZN(new_n683));
  OR3_X1    g0483(.A1(new_n382), .A2(KEYINPUT27), .A3(G20), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT27), .B1(new_n382), .B2(G20), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n684), .A2(G213), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G343), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT89), .Z(new_n688));
  OAI211_X1 g0488(.A(new_n683), .B(new_n666), .C1(new_n516), .C2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n515), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n594), .A2(new_n601), .A3(new_n602), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n688), .A2(new_n598), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n603), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n690), .A2(new_n666), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n693), .A2(new_n688), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n525), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n210), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n526), .A2(new_n497), .A3(new_n490), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n706), .A2(new_n707), .A3(new_n206), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n215), .B2(new_n706), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  NAND4_X1  g0510(.A1(new_n683), .A2(new_n639), .A3(new_n666), .A4(new_n688), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n629), .A2(new_n480), .A3(new_n481), .A4(new_n555), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n578), .A2(G179), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n480), .A2(new_n481), .A3(new_n555), .ZN(new_n716));
  AOI211_X1 g0516(.A(new_n483), .B(new_n569), .C1(new_n577), .C2(new_n278), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT30), .A4(new_n629), .ZN(new_n718));
  INV_X1    g0518(.A(new_n578), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n555), .A2(G179), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n482), .A3(new_n613), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n715), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT31), .B1(new_n722), .B2(new_n690), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n715), .A2(new_n721), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT90), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT90), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n715), .A2(new_n726), .A3(new_n721), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(new_n718), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n688), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n723), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n711), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT91), .B1(new_n732), .B2(G330), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT91), .ZN(new_n734));
  INV_X1    g0534(.A(G330), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n734), .B(new_n735), .C1(new_n711), .C2(new_n731), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n566), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT26), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n739), .A3(new_n677), .ZN(new_n740));
  INV_X1    g0540(.A(new_n565), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT92), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n665), .A2(new_n743), .A3(new_n666), .A4(new_n601), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT92), .B1(new_n693), .B2(new_n515), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(new_n664), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n668), .A2(new_n673), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n740), .B(new_n742), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(KEYINPUT29), .A3(new_n688), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n661), .B(new_n663), .C1(new_n693), .C2(new_n515), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n524), .B2(new_n522), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n678), .A2(KEYINPUT26), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n663), .A2(new_n677), .A3(new_n739), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n565), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n688), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n737), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n710), .B1(new_n760), .B2(G1), .ZN(G364));
  NOR2_X1   g0561(.A1(new_n257), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n206), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n706), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n698), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G330), .B2(new_n696), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n705), .A2(new_n317), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G355), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G116), .B2(new_n210), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n705), .A2(new_n466), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n281), .B2(new_n215), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n241), .A2(new_n281), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n216), .B1(G20), .B2(new_n328), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT93), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(KEYINPUT93), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n765), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n207), .A2(G179), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(G190), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n497), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n207), .A2(new_n483), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n389), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n786), .A2(new_n389), .A3(G200), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n792), .A2(new_n202), .B1(new_n793), .B2(new_n315), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n790), .A2(G190), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n788), .B(new_n794), .C1(G68), .C2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n789), .A2(G190), .A3(new_n289), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT94), .Z(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G58), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G190), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n786), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n395), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT32), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n789), .A2(new_n801), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n317), .B(new_n805), .C1(G77), .C2(new_n807), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n389), .A2(G179), .A3(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n207), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n587), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n804), .B2(new_n803), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n796), .A2(new_n800), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT33), .B(G317), .ZN(new_n814));
  INV_X1    g0614(.A(new_n797), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n795), .A2(new_n814), .B1(new_n815), .B2(G322), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT95), .Z(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n317), .B1(new_n806), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n802), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(G329), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n793), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G303), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n810), .A2(new_n462), .B1(new_n787), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n823), .B(new_n825), .C1(G326), .C2(new_n791), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n817), .A2(new_n821), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n813), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n785), .B1(new_n828), .B2(new_n779), .ZN(new_n829));
  INV_X1    g0629(.A(new_n782), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n696), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n767), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  NAND2_X1  g0633(.A1(new_n331), .A2(new_n688), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n751), .B2(new_n754), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT96), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n680), .A2(KEYINPUT96), .A3(new_n835), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n690), .A2(new_n330), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n690), .A2(new_n313), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n327), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n330), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n755), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n765), .B1(new_n848), .B2(new_n737), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n737), .B2(new_n848), .ZN(new_n850));
  INV_X1    g0650(.A(new_n765), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n779), .A2(new_n780), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(new_n852), .B2(new_n272), .ZN(new_n853));
  INV_X1    g0653(.A(new_n779), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G116), .A2(new_n807), .B1(new_n820), .B2(G311), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n855), .B(new_n317), .C1(new_n462), .C2(new_n797), .ZN(new_n856));
  INV_X1    g0656(.A(new_n787), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n791), .A2(G303), .B1(new_n857), .B2(G107), .ZN(new_n858));
  INV_X1    g0658(.A(new_n795), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n822), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n793), .A2(new_n497), .ZN(new_n861));
  NOR4_X1   g0661(.A1(new_n856), .A2(new_n860), .A3(new_n811), .A4(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n791), .A2(G137), .B1(new_n807), .B2(G159), .ZN(new_n863));
  INV_X1    g0663(.A(G143), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n248), .B2(new_n859), .C1(new_n798), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT34), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n202), .A2(new_n787), .B1(new_n793), .B2(new_n375), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n466), .B1(new_n868), .B2(new_n802), .ZN(new_n869));
  INV_X1    g0669(.A(new_n810), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n867), .B(new_n869), .C1(G58), .C2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n862), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n846), .A2(new_n842), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n853), .B1(new_n854), .B2(new_n872), .C1(new_n873), .C2(new_n781), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n850), .A2(new_n874), .ZN(G384));
  INV_X1    g0675(.A(new_n618), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n876), .A2(KEYINPUT35), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(KEYINPUT35), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(G116), .A3(new_n217), .A4(new_n878), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  OR3_X1    g0680(.A1(new_n214), .A2(new_n272), .A3(new_n398), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n202), .A2(G68), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n206), .B(G13), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n410), .A2(new_n254), .ZN(new_n887));
  INV_X1    g0687(.A(new_n409), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(G68), .A3(new_n407), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT16), .B1(new_n889), .B2(new_n400), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n422), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n686), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n452), .A2(new_n450), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(new_n445), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n449), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n426), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n425), .B1(new_n420), .B2(new_n422), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n899), .B2(new_n440), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n686), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n891), .A2(new_n440), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n892), .A3(new_n449), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n900), .A2(new_n901), .B1(KEYINPUT37), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n886), .B1(new_n894), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n892), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n443), .A2(KEYINPUT76), .A3(new_n444), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n452), .A2(new_n450), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n904), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n688), .A2(new_n386), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n388), .B2(new_n393), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n645), .A2(new_n392), .A3(new_n913), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n873), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n722), .A2(new_n730), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n723), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n666), .B1(new_n668), .B2(new_n673), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n603), .A2(new_n638), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n738), .A3(new_n688), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n885), .B1(new_n912), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n917), .A2(new_n924), .ZN(new_n927));
  INV_X1    g0727(.A(new_n449), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT97), .B1(new_n928), .B2(new_n648), .ZN(new_n929));
  INV_X1    g0729(.A(new_n648), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT97), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n449), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n901), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .B1(new_n901), .B2(new_n900), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n901), .B1(new_n450), .B2(new_n649), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n886), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n911), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n927), .A2(KEYINPUT40), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n454), .A2(new_n923), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(G330), .A3(new_n942), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n454), .A2(new_n749), .A3(new_n757), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n657), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n937), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n388), .A2(new_n690), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT96), .B1(new_n680), .B2(new_n835), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n837), .B(new_n834), .C1(new_n674), .C2(new_n679), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n841), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n905), .A2(new_n911), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n915), .A2(new_n916), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n649), .A2(new_n686), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n946), .B(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n943), .A2(new_n962), .A3(KEYINPUT98), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n206), .B2(new_n762), .C1(new_n962), .C2(new_n943), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT98), .B1(new_n943), .B2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n884), .B1(new_n964), .B2(new_n965), .ZN(G367));
  OAI21_X1  g0766(.A(new_n783), .B1(new_n210), .B2(new_n304), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n772), .A2(new_n237), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n765), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(G137), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n787), .A2(new_n397), .B1(new_n802), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT104), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n792), .A2(new_n864), .B1(new_n375), .B2(new_n810), .ZN(new_n973));
  INV_X1    g0773(.A(new_n793), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(G77), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n859), .B2(new_n395), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n269), .B1(new_n806), .B2(new_n202), .C1(new_n248), .C2(new_n797), .ZN(new_n977));
  NOR4_X1   g0777(.A1(new_n972), .A2(new_n973), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(G317), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n405), .B1(new_n822), .B2(new_n806), .C1(new_n979), .C2(new_n802), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n787), .A2(new_n490), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT46), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(G303), .C2(new_n799), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n859), .A2(new_n462), .B1(new_n315), .B2(new_n810), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n792), .A2(new_n818), .B1(new_n793), .B2(new_n587), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n978), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT47), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n854), .B1(new_n987), .B2(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n969), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n688), .B1(new_n553), .B2(new_n548), .ZN(new_n991));
  MUX2_X1   g0791(.A(new_n663), .B(new_n741), .S(new_n991), .Z(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT99), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n990), .B1(new_n994), .B2(new_n830), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT105), .Z(new_n996));
  INV_X1    g0796(.A(KEYINPUT103), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n689), .A2(new_n691), .A3(new_n701), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n525), .A2(new_n702), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n998), .A2(new_n697), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n697), .B1(new_n998), .B2(new_n999), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT102), .B1(new_n759), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1001), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n697), .A3(new_n999), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT102), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1006), .A2(new_n1007), .A3(new_n737), .A4(new_n758), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT45), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n920), .A2(new_n701), .B1(new_n666), .B2(new_n690), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n620), .A2(new_n622), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n661), .B1(new_n1012), .B2(new_n688), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n677), .A2(new_n690), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1010), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n1015), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1011), .A2(KEYINPUT44), .A3(new_n1016), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT44), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n703), .B2(new_n1015), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n1019), .A2(new_n699), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n699), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n997), .B1(new_n1009), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1028), .A2(new_n1003), .A3(new_n1008), .A4(KEYINPUT103), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n760), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n706), .B(KEYINPUT41), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n764), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n525), .A2(new_n702), .A3(new_n1015), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT42), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n666), .B1(new_n636), .B2(new_n635), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n688), .B1(new_n1037), .B2(new_n677), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1035), .A2(KEYINPUT42), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT100), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT100), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n993), .B(KEYINPUT43), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1041), .A2(new_n1046), .A3(new_n1042), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT101), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1045), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n699), .B2(new_n1016), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n699), .A2(new_n1016), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n1045), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n996), .B1(new_n1034), .B2(new_n1055), .ZN(G387));
  NAND2_X1  g0856(.A1(new_n759), .A2(new_n1002), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT110), .Z(new_n1058));
  XNOR2_X1  g0858(.A(new_n706), .B(KEYINPUT109), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n1009), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1006), .A2(new_n764), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n797), .A2(new_n202), .B1(new_n802), .B2(new_n248), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G68), .B2(new_n807), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n870), .A2(new_n303), .B1(new_n857), .B2(G77), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n246), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G159), .A2(new_n791), .B1(new_n795), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n405), .B1(G97), .B2(new_n974), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n795), .A2(G311), .B1(new_n807), .B2(G303), .ZN(new_n1069));
  INV_X1    g0869(.A(G322), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n792), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G317), .B2(new_n799), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1072), .A2(KEYINPUT48), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n810), .A2(new_n822), .B1(new_n787), .B2(new_n462), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT108), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1072), .A2(KEYINPUT48), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(KEYINPUT49), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n466), .B1(G326), .B2(new_n820), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n490), .C2(new_n793), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT49), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1068), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n779), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n246), .A2(G50), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT50), .ZN(new_n1085));
  AOI211_X1 g0885(.A(G45), .B(new_n707), .C1(G68), .C2(G77), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n772), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n234), .B2(new_n281), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n768), .A2(new_n707), .B1(new_n315), .B2(new_n705), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(KEYINPUT106), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n783), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT106), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n765), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT107), .Z(new_n1094));
  OAI211_X1 g0894(.A(new_n1083), .B(new_n1094), .C1(new_n692), .C2(new_n830), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1061), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1060), .A2(new_n1096), .ZN(G393));
  INV_X1    g0897(.A(new_n1059), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1009), .B2(new_n1026), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1030), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1015), .A2(new_n830), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT111), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n784), .B1(G97), .B2(new_n705), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n771), .A2(new_n244), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n851), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n859), .A2(new_n202), .B1(new_n787), .B2(new_n375), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n466), .B1(new_n864), .B2(new_n802), .C1(new_n246), .C2(new_n806), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n810), .A2(new_n272), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n861), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n792), .A2(new_n248), .B1(new_n395), .B2(new_n797), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT51), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n792), .A2(new_n979), .B1(new_n818), .B2(new_n797), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT52), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n859), .A2(new_n824), .B1(new_n793), .B2(new_n315), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n317), .B1(new_n802), .B2(new_n1070), .C1(new_n462), .C2(new_n806), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n810), .A2(new_n490), .B1(new_n787), .B2(new_n822), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1109), .A2(new_n1111), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1102), .B(new_n1105), .C1(new_n854), .C2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1026), .B2(new_n763), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1100), .A2(new_n1120), .ZN(G390));
  AOI21_X1  g0921(.A(new_n851), .B1(new_n852), .B2(new_n246), .ZN(new_n1122));
  INV_X1    g0922(.A(G128), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n792), .A2(new_n1123), .B1(new_n395), .B2(new_n810), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G137), .B2(new_n795), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n269), .B1(new_n793), .B2(new_n202), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT113), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1125), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n857), .B2(G150), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1131), .A2(new_n787), .A3(new_n248), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n815), .A2(G132), .B1(new_n807), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(G125), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n802), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n1130), .A2(new_n1133), .A3(new_n1134), .A4(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n791), .A2(G283), .B1(new_n807), .B2(G97), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n315), .B2(new_n859), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT115), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n317), .B1(new_n802), .B2(new_n462), .C1(new_n797), .C2(new_n490), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n793), .A2(new_n375), .ZN(new_n1145));
  NOR4_X1   g0945(.A1(new_n1144), .A2(new_n788), .A3(new_n1108), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1140), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(KEYINPUT116), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(KEYINPUT116), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n779), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT39), .B1(new_n911), .B2(new_n936), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n912), .B2(KEYINPUT39), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1122), .B1(new_n1148), .B2(new_n1150), .C1(new_n1152), .C2(new_n781), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n748), .A2(new_n688), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n841), .B1(new_n1154), .B2(new_n846), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n957), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n949), .B1(new_n911), .B2(new_n936), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n873), .B(new_n957), .C1(new_n733), .C2(new_n736), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n949), .B1(new_n954), .B2(new_n957), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(new_n1159), .C1(new_n1152), .C2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n842), .B1(new_n838), .B2(new_n839), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1162), .A2(new_n956), .B1(new_n388), .B2(new_n690), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n948), .A2(new_n950), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1163), .A2(new_n1164), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n923), .A2(G330), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n917), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1161), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1158), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1167), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT112), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n923), .A2(new_n1172), .A3(G330), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n873), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1172), .B1(new_n923), .B2(G330), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n956), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1155), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(new_n1159), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n873), .B1(new_n733), .B2(new_n736), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1167), .B1(new_n1179), .B2(new_n956), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1180), .B2(new_n1162), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1166), .A2(new_n453), .A3(new_n394), .A4(new_n336), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n944), .B(new_n1182), .C1(new_n653), .C2(new_n656), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1171), .A2(new_n1161), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n1059), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1181), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1169), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1153), .B1(new_n763), .B2(new_n1169), .C1(new_n1185), .C2(new_n1188), .ZN(G378));
  NOR2_X1   g0989(.A1(new_n256), .A2(new_n264), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n686), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n301), .B2(new_n335), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n334), .B(new_n1192), .C1(new_n297), .C2(new_n300), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  OR3_X1    g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n956), .B1(new_n840), .B2(new_n841), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n959), .B1(new_n1201), .B2(new_n955), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1200), .B1(new_n1202), .B2(new_n951), .ZN(new_n1203));
  AND4_X1   g1003(.A1(new_n951), .A2(new_n958), .A3(new_n960), .A4(new_n1200), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n926), .A2(G330), .A3(new_n938), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n926), .A2(G330), .A3(new_n938), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1200), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n961), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1202), .A2(new_n951), .A3(new_n1200), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1207), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n764), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT119), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n851), .B1(new_n852), .B2(new_n202), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n797), .A2(new_n1123), .B1(new_n806), .B2(new_n970), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n795), .A2(G132), .B1(new_n857), .B2(new_n1136), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1138), .B2(new_n792), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(G150), .C2(new_n870), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n974), .A2(G159), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G33), .B(G41), .C1(new_n820), .C2(G124), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n791), .A2(G116), .B1(new_n974), .B2(G58), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n587), .B2(new_n859), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n815), .A2(G107), .B1(new_n820), .B2(G283), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n304), .B2(new_n806), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n405), .A2(new_n280), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n810), .A2(new_n375), .B1(new_n787), .B2(new_n272), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1226), .A2(new_n1228), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  XOR2_X1   g1032(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1233));
  OR2_X1    g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1229), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1236));
  AND4_X1   g1036(.A1(new_n1224), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1214), .B1(new_n854), .B2(new_n1237), .C1(new_n1200), .C2(new_n781), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT118), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1212), .A2(new_n1213), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1205), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1209), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n763), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1239), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT119), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1240), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1183), .B1(new_n1169), .B2(new_n1186), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(KEYINPUT57), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1184), .A2(new_n1183), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1249), .B(new_n1059), .C1(new_n1250), .C2(KEYINPUT57), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1246), .A2(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n956), .A2(new_n780), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n859), .A2(new_n1135), .B1(new_n787), .B2(new_n395), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G50), .B2(new_n870), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n799), .A2(G137), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n806), .A2(new_n248), .B1(new_n802), .B2(new_n1123), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(new_n405), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n791), .A2(G132), .B1(new_n974), .B2(G58), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1255), .A2(new_n1256), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n792), .A2(new_n462), .B1(new_n787), .B2(new_n587), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G116), .B2(new_n795), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n870), .A2(new_n303), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n797), .A2(new_n822), .B1(new_n802), .B2(new_n824), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n269), .B(new_n1264), .C1(G107), .C2(new_n807), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n975), .A3(new_n1263), .A4(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n854), .B1(new_n1260), .B2(new_n1266), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n851), .B(new_n1267), .C1(new_n375), .C2(new_n852), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1181), .A2(new_n764), .B1(new_n1253), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1186), .A2(new_n1033), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1183), .A2(new_n1181), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(G381));
  XOR2_X1   g1072(.A(G375), .B(KEYINPUT120), .Z(new_n1273));
  NAND3_X1  g1073(.A1(new_n1060), .A2(new_n832), .A3(new_n1096), .ZN(new_n1274));
  NOR4_X1   g1074(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1153), .B1(new_n1169), .B2(new_n763), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1185), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1277), .B2(new_n1187), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  OR3_X1    g1079(.A1(new_n1273), .A2(G387), .A3(new_n1279), .ZN(G407));
  INV_X1    g1080(.A(G343), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(G213), .ZN(new_n1282));
  OR3_X1    g1082(.A1(new_n1273), .A2(G378), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G407), .A2(new_n1283), .A3(G213), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT121), .Z(G409));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1100), .A2(new_n1120), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(G387), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1274), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n832), .B1(new_n1060), .B2(new_n1096), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(G387), .A2(new_n1287), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1032), .B1(new_n1030), .B2(new_n760), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1052), .B(new_n1054), .C1(new_n1293), .C2(new_n764), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G390), .B1(new_n1294), .B2(new_n996), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n1288), .A2(new_n1291), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(new_n1287), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(G390), .A2(new_n1294), .A3(new_n996), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1291), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1297), .A2(new_n1286), .A3(new_n1298), .A4(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1246), .A2(new_n1251), .A3(G378), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1212), .A2(new_n1239), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1247), .A2(new_n1248), .A3(new_n1033), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1278), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1282), .ZN(new_n1307));
  OR2_X1    g1107(.A1(new_n1180), .A2(new_n1162), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1182), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n652), .B1(new_n651), .B2(new_n335), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n655), .A2(KEYINPUT88), .A3(new_n334), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n945), .B(new_n1309), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1308), .A2(KEYINPUT60), .A3(new_n1312), .A4(new_n1178), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1183), .B2(new_n1181), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1059), .B(new_n1313), .C1(new_n1316), .C2(new_n1271), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1317), .A2(G384), .A3(new_n1269), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G384), .B1(new_n1317), .B2(new_n1269), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1281), .A2(G213), .A3(G2897), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1320), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(KEYINPUT124), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT124), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1324), .B(new_n1320), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1321), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1307), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT126), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1306), .A2(new_n1282), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT62), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1306), .A2(new_n1333), .A3(new_n1282), .A4(new_n1330), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1329), .A2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1326), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(KEYINPUT126), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1301), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT63), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1337), .B(new_n1301), .C1(new_n1340), .C2(new_n1331), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1331), .A2(new_n1340), .ZN(new_n1342));
  OR2_X1    g1142(.A1(new_n1342), .A2(KEYINPUT123), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(KEYINPUT123), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1341), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT127), .B1(new_n1339), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1301), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1332), .B(new_n1334), .C1(new_n1337), .C2(KEYINPUT126), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1337), .A2(KEYINPUT126), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1347), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT127), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1350), .B(new_n1351), .C1(new_n1352), .C2(new_n1341), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1346), .A2(new_n1353), .ZN(G405));
  XNOR2_X1  g1154(.A(G375), .B(G378), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1301), .B(new_n1355), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1356), .B(new_n1330), .ZN(G402));
endmodule


