//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  XNOR2_X1  g000(.A(G143), .B(G146), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n187), .A2(new_n189), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT66), .A2(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT66), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n191), .A2(new_n192), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(new_n187), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT11), .A2(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT64), .A2(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT11), .A2(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT11), .A2(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n199), .A2(new_n208), .A3(new_n201), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n206), .B1(G134), .B2(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n196), .A2(new_n207), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT70), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT2), .A2(G113), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT69), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G119), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n222), .A3(G116), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT2), .A2(G113), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n219), .A2(G116), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n218), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n218), .A2(new_n224), .B1(new_n223), .B2(new_n225), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n207), .A2(new_n211), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(new_n196), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G146), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n194), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT0), .B(G128), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n187), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n202), .A2(new_n206), .A3(new_n205), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n206), .B1(new_n202), .B2(new_n205), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n213), .A2(new_n229), .A3(new_n232), .A4(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n202), .A2(new_n205), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n238), .B1(new_n247), .B2(new_n207), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(KEYINPUT70), .B2(new_n212), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(KEYINPUT72), .A3(new_n229), .A4(new_n232), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n253), .B(KEYINPUT27), .Z(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT65), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n212), .B1(new_n248), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT67), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n247), .A2(new_n207), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n261), .A3(new_n239), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n212), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n260), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n213), .A2(KEYINPUT30), .A3(new_n232), .A4(new_n242), .ZN(new_n273));
  INV_X1    g087(.A(new_n229), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT71), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n274), .ZN(new_n278));
  AOI211_X1 g092(.A(new_n277), .B(new_n278), .C1(new_n265), .C2(new_n271), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n259), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT31), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n269), .A2(new_n274), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n251), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT28), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n274), .A2(new_n248), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT28), .B1(new_n285), .B2(new_n212), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n256), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n242), .A2(KEYINPUT65), .B1(new_n196), .B2(new_n230), .ZN(new_n290));
  AOI211_X1 g104(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n290), .C2(new_n268), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n270), .B1(new_n269), .B2(new_n260), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n275), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n277), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n272), .A2(KEYINPUT71), .A3(new_n275), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n259), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n281), .A2(new_n289), .A3(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G472), .A2(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n300), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(new_n302), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT74), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n296), .A2(new_n251), .A3(new_n256), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n256), .B1(new_n284), .B2(new_n287), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n249), .A2(new_n232), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n274), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n251), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n286), .B1(new_n314), .B2(KEYINPUT28), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(KEYINPUT73), .A3(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n245), .A2(new_n250), .B1(new_n312), .B2(new_n274), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n287), .B(new_n316), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G902), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G472), .B1(new_n311), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n299), .A2(new_n327), .A3(new_n305), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n303), .A2(new_n307), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT9), .B(G234), .ZN(new_n330));
  OAI21_X1  g144(.A(G221), .B1(new_n330), .B2(G902), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G140), .ZN(new_n333));
  INV_X1    g147(.A(G227), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G953), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n267), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(KEYINPUT12), .ZN(new_n341));
  INV_X1    g155(.A(G104), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G107), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G107), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n343), .A2(new_n344), .ZN(new_n349));
  OAI21_X1  g163(.A(G101), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n346), .A3(G104), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(new_n343), .ZN(new_n353));
  INV_X1    g167(.A(G101), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT3), .B1(new_n342), .B2(G107), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n347), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n353), .A2(new_n354), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n188), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n190), .B1(new_n187), .B2(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n350), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n196), .B1(new_n359), .B2(new_n350), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n339), .B(new_n341), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n350), .A2(new_n359), .ZN(new_n365));
  INV_X1    g179(.A(new_n196), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n350), .A2(new_n359), .A3(new_n361), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n340), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n338), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT12), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT80), .B1(new_n367), .B2(new_n368), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n372), .B2(new_n267), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n352), .B(new_n343), .C1(new_n355), .C2(new_n356), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT78), .B1(new_n347), .B2(KEYINPUT3), .ZN(new_n376));
  OAI21_X1  g190(.A(G101), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT4), .A3(new_n359), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(G101), .C1(new_n375), .C2(new_n376), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n239), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n368), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n196), .A2(new_n350), .A3(new_n359), .A4(KEYINPUT10), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n381), .A2(new_n338), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n337), .B1(new_n374), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n385), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(new_n336), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n267), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT82), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n390), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT82), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n370), .A2(new_n373), .A3(new_n387), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n393), .B(new_n394), .C1(new_n395), .C2(new_n337), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(G469), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G469), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(new_n324), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n374), .A2(new_n388), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n390), .A2(new_n385), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n336), .ZN(new_n402));
  AOI21_X1  g216(.A(G902), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n399), .B1(new_n403), .B2(new_n398), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n332), .B1(new_n397), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G475), .ZN(new_n406));
  INV_X1    g220(.A(G140), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G125), .ZN(new_n408));
  INV_X1    g222(.A(G125), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G140), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n410), .A3(KEYINPUT16), .ZN(new_n411));
  OR3_X1    g225(.A1(new_n409), .A2(KEYINPUT16), .A3(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n193), .ZN(new_n414));
  AOI21_X1  g228(.A(G146), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n252), .A2(G214), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n233), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n252), .A2(G143), .A3(G214), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n206), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT17), .ZN(new_n421));
  INV_X1    g235(.A(new_n419), .ZN(new_n422));
  AOI21_X1  g236(.A(G143), .B1(new_n252), .B2(G214), .ZN(new_n423));
  OAI21_X1  g237(.A(G131), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(new_n206), .A3(new_n419), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n416), .B(new_n421), .C1(new_n426), .C2(KEYINPUT17), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n408), .A2(new_n410), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n408), .A2(new_n410), .A3(KEYINPUT89), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(G146), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n408), .A2(new_n410), .A3(new_n193), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n422), .A2(new_n423), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT18), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n435), .B1(new_n436), .B2(new_n206), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT18), .B(G131), .C1(new_n422), .C2(new_n423), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n427), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G113), .B(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT92), .B(G104), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n441), .B(new_n442), .Z(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n427), .A2(new_n443), .A3(new_n439), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n406), .B1(new_n447), .B2(new_n324), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n430), .A2(KEYINPUT19), .A3(new_n431), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n428), .A2(KEYINPUT19), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n193), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n414), .A2(KEYINPUT75), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n413), .B2(new_n193), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n422), .A2(new_n423), .A3(G131), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT90), .B1(new_n456), .B2(new_n420), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n424), .A2(new_n425), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n439), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT91), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT91), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n439), .C1(new_n455), .C2(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n444), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n446), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT93), .ZN(new_n467));
  NOR2_X1   g281(.A1(G475), .A2(G902), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT93), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n446), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT20), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n466), .A2(new_n475), .A3(new_n468), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n448), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G116), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n346), .B1(new_n479), .B2(KEYINPUT14), .ZN(new_n480));
  XNOR2_X1  g294(.A(G116), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n191), .A2(G143), .A3(new_n192), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT95), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n188), .A2(G143), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n484), .B1(new_n483), .B2(new_n486), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n208), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n488), .A2(new_n208), .A3(new_n489), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n482), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n481), .B(new_n346), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n485), .A2(KEYINPUT13), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n485), .A2(KEYINPUT13), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n483), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(G134), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n497), .B2(G134), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n490), .B(new_n494), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G217), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n330), .A2(new_n503), .A3(G953), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n493), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n493), .B2(new_n502), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT96), .ZN(new_n510));
  INV_X1    g324(.A(G478), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n509), .A2(new_n510), .A3(new_n324), .A4(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n508), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n515), .A2(new_n510), .A3(new_n324), .A4(new_n506), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n512), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G953), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n519), .A2(G952), .ZN(new_n520));
  INV_X1    g334(.A(G234), .ZN(new_n521));
  INV_X1    g335(.A(G237), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI211_X1 g338(.A(new_n324), .B(new_n519), .C1(G234), .C2(G237), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT21), .B(G898), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n405), .A2(new_n477), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n223), .A2(KEYINPUT5), .A3(new_n225), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT69), .B(G119), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT5), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(G116), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(G113), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n534), .A2(new_n226), .A3(new_n359), .A4(new_n350), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n377), .A2(KEYINPUT4), .A3(new_n359), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n380), .B1(new_n227), .B2(new_n228), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(G110), .B(G122), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n535), .B(new_n539), .C1(new_n536), .C2(new_n537), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(KEYINPUT6), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n538), .A2(new_n544), .A3(new_n540), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n366), .A2(new_n409), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT83), .B1(new_n239), .B2(new_n409), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT83), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n238), .A2(new_n548), .A3(G125), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G224), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(G953), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n550), .B(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n543), .A2(new_n545), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n546), .A2(new_n547), .A3(new_n549), .A4(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n239), .A2(new_n409), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n196), .A2(G125), .ZN(new_n559));
  OAI22_X1  g373(.A1(new_n558), .A2(new_n559), .B1(new_n555), .B2(new_n552), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n539), .B(KEYINPUT8), .Z(new_n562));
  NAND2_X1  g376(.A1(new_n534), .A2(new_n226), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n365), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n564), .B2(new_n535), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n566), .B2(new_n542), .ZN(new_n567));
  OAI21_X1  g381(.A(G210), .B1(G237), .B2(G902), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n554), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT87), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT87), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n568), .B(KEYINPUT85), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n554), .A2(new_n567), .A3(KEYINPUT84), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT84), .B1(new_n554), .B2(new_n567), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT86), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT86), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n581), .B(new_n575), .C1(new_n577), .C2(new_n578), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n574), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G214), .B1(G237), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n529), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n519), .A2(G221), .A3(G234), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n191), .A2(new_n192), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n591), .A2(G119), .B1(new_n531), .B2(G128), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT24), .B(G110), .Z(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n220), .A2(new_n222), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT23), .B1(new_n595), .B2(new_n188), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n191), .A2(new_n192), .ZN(new_n597));
  OAI22_X1  g411(.A1(new_n219), .A2(new_n597), .B1(new_n595), .B2(new_n188), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n598), .B2(KEYINPUT23), .ZN(new_n599));
  INV_X1    g413(.A(G110), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n594), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n452), .A2(new_n454), .A3(new_n433), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n599), .A2(new_n600), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n592), .A2(new_n593), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(new_n414), .B2(new_n415), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n590), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  OAI221_X1 g422(.A(new_n605), .B1(new_n415), .B2(new_n414), .C1(new_n599), .C2(new_n600), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n609), .B(new_n589), .C1(new_n601), .C2(new_n602), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n324), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT25), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n608), .A2(KEYINPUT25), .A3(new_n324), .A4(new_n610), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n503), .B1(G234), .B2(new_n324), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n608), .A2(new_n610), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n616), .A2(G902), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT76), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n617), .A2(KEYINPUT77), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT77), .B1(new_n617), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n329), .A2(new_n586), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  INV_X1    g440(.A(new_n624), .ZN(new_n627));
  INV_X1    g441(.A(new_n405), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G472), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n299), .A2(new_n324), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n299), .B2(new_n324), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n568), .B1(new_n554), .B2(new_n567), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n570), .B2(KEYINPUT98), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n569), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n585), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n527), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n515), .A2(new_n506), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n643), .A2(KEYINPUT33), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n493), .A2(new_n502), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n504), .B1(new_n646), .B2(KEYINPUT100), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT99), .B1(new_n504), .B2(KEYINPUT100), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n493), .B2(new_n502), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT33), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n644), .A2(G478), .A3(new_n324), .A4(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n511), .B1(new_n643), .B2(G902), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n476), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n471), .B2(new_n473), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n653), .B1(new_n655), .B2(new_n448), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n642), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n635), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT101), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  NAND4_X1  g475(.A1(new_n467), .A2(new_n468), .A3(new_n470), .A4(new_n472), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n448), .B1(new_n474), .B2(new_n662), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n641), .A2(new_n663), .A3(new_n518), .A4(new_n640), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n635), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT102), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT35), .B(G107), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  INV_X1    g482(.A(new_n616), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n613), .B2(new_n614), .ZN(new_n670));
  OR4_X1    g484(.A1(KEYINPUT36), .A2(new_n603), .A3(new_n607), .A4(new_n590), .ZN(new_n671));
  OAI22_X1  g485(.A1(new_n603), .A2(new_n607), .B1(KEYINPUT36), .B2(new_n590), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n671), .A2(new_n620), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n586), .A2(new_n634), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  NAND3_X1  g492(.A1(new_n405), .A2(new_n640), .A3(new_n675), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n525), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n523), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n663), .A2(new_n518), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n329), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n188), .ZN(G30));
  XNOR2_X1  g500(.A(new_n682), .B(KEYINPUT39), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n628), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT40), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n518), .B1(new_n655), .B2(new_n448), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n691), .A2(new_n585), .A3(new_n675), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n583), .B(new_n694), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n689), .A2(new_n690), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n307), .A2(new_n328), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n294), .A2(new_n295), .B1(new_n245), .B2(new_n250), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n256), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n324), .B1(new_n314), .B2(new_n257), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n303), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n693), .A2(new_n695), .A3(new_n696), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  OAI211_X1 g519(.A(new_n653), .B(new_n682), .C1(new_n655), .C2(new_n448), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n679), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n329), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n193), .ZN(G48));
  OR2_X1    g523(.A1(new_n403), .A2(new_n398), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n403), .A2(new_n398), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n331), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n329), .A2(new_n657), .A3(new_n624), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND4_X1  g530(.A1(new_n329), .A2(new_n624), .A3(new_n664), .A4(new_n713), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  INV_X1    g532(.A(new_n640), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n712), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n477), .A2(new_n528), .A3(new_n675), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n329), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  OAI211_X1 g537(.A(new_n281), .B(new_n298), .C1(new_n257), .C2(new_n315), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n300), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n299), .A2(new_n324), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT105), .B(G472), .Z(new_n728));
  AOI22_X1  g542(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n710), .A2(new_n641), .A3(new_n331), .A4(new_n711), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n719), .A2(new_n692), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n617), .A2(new_n621), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n724), .A2(KEYINPUT104), .A3(new_n300), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n729), .A2(new_n731), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NOR3_X1   g550(.A1(new_n719), .A2(new_n706), .A3(new_n712), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n729), .A3(new_n675), .A4(new_n734), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT106), .B(G125), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G27));
  AND3_X1   g554(.A1(new_n571), .A2(new_n584), .A3(new_n573), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n386), .A2(new_n391), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n332), .B1(new_n404), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n582), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n554), .A2(new_n567), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT84), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n576), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n581), .B1(new_n749), .B2(new_n575), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n741), .B(new_n744), .C1(new_n745), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n706), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n297), .B1(new_n296), .B2(new_n259), .ZN(new_n753));
  AOI211_X1 g567(.A(KEYINPUT31), .B(new_n258), .C1(new_n294), .C2(new_n295), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n304), .B1(new_n755), .B2(new_n289), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n326), .B1(new_n756), .B2(KEYINPUT32), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n624), .B(new_n752), .C1(new_n697), .C2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  AOI21_X1  g573(.A(G902), .B1(new_n317), .B2(new_n322), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n309), .B1(new_n698), .B2(new_n256), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(KEYINPUT29), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n302), .A2(new_n301), .B1(new_n762), .B2(G472), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n732), .B1(new_n763), .B2(new_n306), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n751), .A2(new_n759), .A3(new_n706), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n758), .A2(new_n759), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n206), .ZN(G33));
  NOR2_X1   g581(.A1(new_n751), .A2(new_n683), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n329), .A2(new_n624), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(new_n448), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n471), .A2(new_n473), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(new_n654), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT107), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT43), .A3(new_n653), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n776));
  INV_X1    g590(.A(new_n653), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n776), .B1(new_n773), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n634), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n780), .A3(new_n675), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n741), .B1(new_n745), .B2(new_n750), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n742), .A2(KEYINPUT45), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(G469), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT45), .B1(new_n392), .B2(new_n396), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n399), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT46), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n711), .B1(new_n790), .B2(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n331), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n688), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n781), .A2(new_n782), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n783), .A2(new_n785), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT108), .B(G137), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(G39));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n793), .B(new_n799), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n329), .A2(new_n624), .A3(new_n706), .A4(new_n784), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  NOR3_X1   g617(.A1(new_n695), .A2(new_n584), .A3(new_n712), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n729), .A2(new_n734), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n733), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n806), .A3(new_n524), .A4(new_n779), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n806), .A2(new_n524), .A3(new_n779), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n710), .A2(new_n711), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n331), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n810), .B(new_n785), .C1(new_n800), .C2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n785), .A2(new_n524), .A3(new_n713), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n775), .B2(new_n778), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n675), .A3(new_n805), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n703), .A2(new_n627), .A3(new_n814), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(KEYINPUT116), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(KEYINPUT116), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n477), .A3(new_n777), .A4(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n809), .A2(new_n813), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n821), .A2(new_n822), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n773), .A2(new_n818), .A3(new_n653), .A4(new_n819), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n810), .A2(new_n720), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n815), .A2(new_n829), .A3(KEYINPUT48), .A4(new_n764), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n815), .A2(new_n764), .ZN(new_n831));
  XNOR2_X1  g645(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n828), .A2(new_n520), .A3(new_n830), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n825), .A2(new_n826), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n329), .B1(new_n684), .B2(new_n707), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n744), .A2(new_n674), .A3(new_n682), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n719), .A3(new_n692), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n697), .B2(new_n702), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n738), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT111), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n838), .A2(new_n841), .A3(new_n738), .A4(KEYINPUT52), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(new_n845), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n514), .A2(new_n517), .A3(KEYINPUT109), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT109), .B1(new_n514), .B2(new_n517), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n477), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n527), .B1(new_n854), .B2(new_n656), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n583), .A2(new_n585), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n629), .A2(new_n634), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n625), .A2(new_n676), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n853), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n674), .B1(new_n523), .B2(new_n681), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n663), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n861), .A2(new_n784), .A3(new_n628), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n329), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n752), .A2(new_n729), .A3(new_n734), .A4(new_n675), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n769), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT110), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n769), .A2(new_n863), .A3(new_n864), .A4(KEYINPUT110), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n850), .B(new_n858), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n714), .A2(new_n717), .A3(new_n722), .A4(new_n735), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT114), .B1(new_n870), .B2(new_n766), .ZN(new_n871));
  OR3_X1    g685(.A1(new_n870), .A2(new_n766), .A3(KEYINPUT114), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n849), .A2(new_n869), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n870), .A2(new_n766), .A3(new_n858), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n844), .A2(new_n846), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n867), .A2(new_n868), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n877), .A2(KEYINPUT113), .A3(new_n850), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT113), .B1(new_n877), .B2(new_n850), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n837), .B(new_n873), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n880), .A2(KEYINPUT115), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n849), .A2(new_n876), .A3(new_n874), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n877), .A2(new_n850), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n882), .A2(KEYINPUT53), .B1(KEYINPUT112), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n877), .A2(new_n850), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT112), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT54), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n880), .A2(KEYINPUT115), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n881), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n836), .A2(new_n890), .B1(G952), .B2(G953), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n733), .A2(new_n584), .A3(new_n331), .A4(new_n653), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(KEYINPUT49), .B2(new_n811), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n774), .B(new_n893), .C1(KEYINPUT49), .C2(new_n811), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n894), .A2(new_n703), .A3(new_n695), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n895), .ZN(G75));
  NAND2_X1  g710(.A1(new_n877), .A2(new_n850), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT113), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n877), .A2(KEYINPUT113), .A3(new_n850), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n324), .B1(new_n901), .B2(new_n873), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT56), .B1(new_n902), .B2(G210), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n543), .A2(new_n545), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT119), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n553), .B(KEYINPUT55), .Z(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n902), .B2(new_n575), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n519), .A2(G952), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(G51));
  XNOR2_X1  g727(.A(new_n399), .B(KEYINPUT57), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n837), .B1(new_n901), .B2(new_n873), .ZN(new_n915));
  INV_X1    g729(.A(new_n880), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT121), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n400), .A2(new_n402), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(new_n914), .C1(new_n915), .C2(new_n916), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n789), .B(KEYINPUT122), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n902), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n912), .B1(new_n922), .B2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n467), .A2(new_n470), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n926), .A2(new_n928), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n912), .ZN(G60));
  AND2_X1   g745(.A1(new_n644), .A2(new_n650), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT59), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n932), .B1(new_n890), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n912), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n915), .A2(new_n916), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n932), .A2(new_n934), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n935), .A2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(new_n901), .A2(new_n873), .ZN(new_n941));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT60), .Z(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n618), .B(KEYINPUT123), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n941), .A2(new_n671), .A3(new_n672), .A4(new_n943), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n936), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n936), .A4(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G66));
  OAI21_X1  g766(.A(G953), .B1(new_n526), .B2(new_n551), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n870), .A2(new_n858), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(G953), .ZN(new_n955));
  INV_X1    g769(.A(new_n905), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(G898), .B2(new_n519), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G69));
  NAND2_X1  g772(.A1(new_n272), .A2(new_n273), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n449), .A2(new_n450), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n959), .B(new_n960), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n796), .A2(new_n802), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n719), .A2(new_n692), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n794), .A2(new_n964), .A3(new_n764), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n838), .A2(new_n769), .A3(new_n738), .ZN(new_n966));
  OR3_X1    g780(.A1(new_n965), .A2(new_n766), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n519), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n680), .A2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n968), .A2(new_n972), .A3(new_n969), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n962), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(G953), .B1(new_n334), .B2(new_n680), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT125), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n704), .A2(new_n738), .A3(new_n838), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n784), .B1(new_n656), .B2(new_n854), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n329), .A2(new_n980), .A3(new_n624), .A4(new_n689), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT124), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n983), .A2(new_n963), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n961), .B1(new_n984), .B2(new_n519), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n974), .A2(new_n976), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n976), .B1(new_n974), .B2(new_n985), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(G72));
  NOR2_X1   g802(.A1(new_n884), .A2(new_n887), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n308), .A2(new_n991), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n989), .A2(new_n699), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n954), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n991), .B1(new_n984), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n995), .A2(new_n699), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n963), .A2(new_n994), .A3(new_n967), .ZN(new_n997));
  INV_X1    g811(.A(new_n991), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n256), .B(new_n698), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n936), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(KEYINPUT127), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n999), .A2(new_n1002), .A3(new_n936), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n993), .B(new_n996), .C1(new_n1001), .C2(new_n1003), .ZN(G57));
endmodule


