

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728;

  INV_X2 U372 ( .A(G953), .ZN(n722) );
  XOR2_X1 U373 ( .A(G146), .B(G125), .Z(n426) );
  INV_X1 U374 ( .A(n470), .ZN(n669) );
  NOR2_X1 U375 ( .A1(n511), .A2(n639), .ZN(n656) );
  NAND2_X2 U376 ( .A1(n460), .A2(n459), .ZN(n504) );
  XNOR2_X2 U377 ( .A(n539), .B(n538), .ZN(n614) );
  NOR2_X2 U378 ( .A1(G953), .A2(G237), .ZN(n431) );
  NOR2_X1 U379 ( .A1(n715), .A2(KEYINPUT81), .ZN(n580) );
  XNOR2_X1 U380 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X2 U381 ( .A(n712), .B(n365), .ZN(n395) );
  XNOR2_X2 U382 ( .A(n466), .B(KEYINPUT19), .ZN(n520) );
  AND2_X2 U383 ( .A1(n520), .A2(n519), .ZN(n521) );
  INV_X1 U384 ( .A(KEYINPUT70), .ZN(n407) );
  OR2_X2 U385 ( .A1(n619), .A2(G902), .ZN(n356) );
  XNOR2_X1 U386 ( .A(n374), .B(n373), .ZN(n375) );
  NOR2_X1 U387 ( .A1(n471), .A2(n465), .ZN(n496) );
  XNOR2_X1 U388 ( .A(n452), .B(n359), .ZN(n385) );
  XNOR2_X1 U389 ( .A(n513), .B(KEYINPUT33), .ZN(n683) );
  XNOR2_X1 U390 ( .A(n398), .B(KEYINPUT96), .ZN(n399) );
  XNOR2_X1 U391 ( .A(G113), .B(G143), .ZN(n428) );
  XNOR2_X1 U392 ( .A(G107), .B(G104), .ZN(n366) );
  XNOR2_X1 U393 ( .A(n355), .B(n354), .ZN(n476) );
  INV_X1 U394 ( .A(KEYINPUT30), .ZN(n354) );
  XNOR2_X1 U395 ( .A(n419), .B(KEYINPUT25), .ZN(n420) );
  XNOR2_X1 U396 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U397 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U398 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U399 ( .A(n491), .B(KEYINPUT40), .ZN(n726) );
  AND2_X1 U400 ( .A1(n353), .A2(n639), .ZN(n491) );
  AND2_X1 U401 ( .A1(n594), .A2(n611), .ZN(G63) );
  XOR2_X1 U402 ( .A(n609), .B(n608), .Z(n352) );
  AND2_X1 U403 ( .A1(n593), .A2(G953), .ZN(n697) );
  INV_X1 U404 ( .A(n697), .ZN(n611) );
  NAND2_X1 U405 ( .A1(n353), .A2(n511), .ZN(n646) );
  XNOR2_X2 U406 ( .A(n490), .B(KEYINPUT39), .ZN(n353) );
  NAND2_X1 U407 ( .A1(n470), .A2(n494), .ZN(n355) );
  XNOR2_X2 U408 ( .A(n356), .B(n396), .ZN(n470) );
  XNOR2_X2 U409 ( .A(n357), .B(G143), .ZN(n452) );
  XNOR2_X2 U410 ( .A(G128), .B(KEYINPUT79), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U412 ( .A(n592), .B(n591), .ZN(n594) );
  BUF_X1 U413 ( .A(n616), .Z(n693) );
  BUF_X1 U414 ( .A(n470), .Z(n558) );
  XNOR2_X2 U415 ( .A(n553), .B(KEYINPUT106), .ZN(n728) );
  NOR2_X2 U416 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X2 U417 ( .A1(n599), .A2(n697), .ZN(n600) );
  XNOR2_X1 U418 ( .A(n509), .B(KEYINPUT38), .ZN(n651) );
  AND2_X1 U419 ( .A1(G210), .A2(n457), .ZN(n358) );
  INV_X1 U420 ( .A(KEYINPUT73), .ZN(n373) );
  XNOR2_X1 U421 ( .A(n369), .B(n368), .ZN(n370) );
  NOR2_X1 U422 ( .A1(n637), .A2(n652), .ZN(n459) );
  XNOR2_X1 U423 ( .A(n376), .B(n375), .ZN(n379) );
  NOR2_X1 U424 ( .A1(n652), .A2(n651), .ZN(n658) );
  XNOR2_X1 U425 ( .A(n498), .B(n497), .ZN(n727) );
  NOR2_X1 U426 ( .A1(n478), .A2(n477), .ZN(n635) );
  XNOR2_X1 U427 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n503) );
  XNOR2_X1 U428 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n359) );
  INV_X1 U429 ( .A(G137), .ZN(n360) );
  XNOR2_X1 U430 ( .A(n360), .B(G134), .ZN(n362) );
  XNOR2_X1 U431 ( .A(G131), .B(KEYINPUT68), .ZN(n361) );
  XNOR2_X1 U432 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n385), .B(n363), .ZN(n712) );
  INV_X1 U434 ( .A(KEYINPUT66), .ZN(n364) );
  XNOR2_X1 U435 ( .A(n364), .B(G101), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n380), .B(G146), .ZN(n365) );
  XNOR2_X1 U437 ( .A(n366), .B(G110), .ZN(n376) );
  NAND2_X1 U438 ( .A1(G227), .A2(n722), .ZN(n367) );
  XNOR2_X1 U439 ( .A(n376), .B(n367), .ZN(n369) );
  XNOR2_X1 U440 ( .A(G140), .B(KEYINPUT95), .ZN(n368) );
  XNOR2_X1 U441 ( .A(n395), .B(n370), .ZN(n609) );
  NOR2_X1 U442 ( .A1(n609), .A2(G902), .ZN(n371) );
  XNOR2_X2 U443 ( .A(n371), .B(G469), .ZN(n471) );
  INV_X1 U444 ( .A(KEYINPUT1), .ZN(n372) );
  XNOR2_X2 U445 ( .A(n471), .B(n372), .ZN(n662) );
  XNOR2_X1 U446 ( .A(n662), .B(KEYINPUT91), .ZN(n531) );
  XNOR2_X1 U447 ( .A(G122), .B(KEYINPUT16), .ZN(n374) );
  XNOR2_X1 U448 ( .A(G116), .B(G113), .ZN(n378) );
  XNOR2_X1 U449 ( .A(KEYINPUT3), .B(G119), .ZN(n377) );
  XNOR2_X1 U450 ( .A(n378), .B(n377), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n379), .B(n393), .ZN(n698) );
  XNOR2_X1 U452 ( .A(n380), .B(n426), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n698), .B(n381), .ZN(n388) );
  XOR2_X1 U454 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n383) );
  NAND2_X1 U455 ( .A1(G224), .A2(n722), .ZN(n382) );
  XNOR2_X1 U456 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U457 ( .A(n384), .B(KEYINPUT75), .Z(n386) );
  XNOR2_X1 U458 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U459 ( .A(n388), .B(n387), .ZN(n601) );
  XNOR2_X1 U460 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n389) );
  XNOR2_X2 U461 ( .A(n389), .B(G902), .ZN(n590) );
  NAND2_X1 U462 ( .A1(n601), .A2(n590), .ZN(n390) );
  OR2_X1 U463 ( .A1(G237), .A2(G902), .ZN(n457) );
  XNOR2_X2 U464 ( .A(n390), .B(n358), .ZN(n509) );
  INV_X1 U465 ( .A(n509), .ZN(n478) );
  NAND2_X1 U466 ( .A1(n431), .A2(G210), .ZN(n391) );
  XNOR2_X1 U467 ( .A(n391), .B(KEYINPUT5), .ZN(n392) );
  XNOR2_X1 U468 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U469 ( .A(n395), .B(n394), .ZN(n619) );
  XNOR2_X1 U470 ( .A(G472), .B(KEYINPUT72), .ZN(n396) );
  XNOR2_X2 U471 ( .A(n669), .B(KEYINPUT6), .ZN(n547) );
  NAND2_X1 U472 ( .A1(n590), .A2(G234), .ZN(n397) );
  XNOR2_X1 U473 ( .A(KEYINPUT20), .B(n397), .ZN(n418) );
  NAND2_X1 U474 ( .A1(n418), .A2(G221), .ZN(n398) );
  XOR2_X1 U475 ( .A(KEYINPUT21), .B(n399), .Z(n666) );
  NAND2_X1 U476 ( .A1(G234), .A2(G237), .ZN(n400) );
  XNOR2_X1 U477 ( .A(n400), .B(KEYINPUT14), .ZN(n403) );
  NAND2_X1 U478 ( .A1(G902), .A2(n403), .ZN(n515) );
  NOR2_X1 U479 ( .A1(G900), .A2(n515), .ZN(n401) );
  NAND2_X1 U480 ( .A1(G953), .A2(n401), .ZN(n402) );
  XNOR2_X1 U481 ( .A(KEYINPUT107), .B(n402), .ZN(n405) );
  NAND2_X1 U482 ( .A1(G952), .A2(n403), .ZN(n404) );
  XNOR2_X1 U483 ( .A(KEYINPUT94), .B(n404), .ZN(n680) );
  NOR2_X1 U484 ( .A1(G953), .A2(n680), .ZN(n514) );
  NOR2_X1 U485 ( .A1(n405), .A2(n514), .ZN(n406) );
  XOR2_X1 U486 ( .A(n406), .B(KEYINPUT80), .Z(n472) );
  NAND2_X1 U487 ( .A1(n666), .A2(n472), .ZN(n408) );
  XNOR2_X1 U488 ( .A(n408), .B(n407), .ZN(n423) );
  XOR2_X1 U489 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n411) );
  NAND2_X1 U490 ( .A1(G234), .A2(n722), .ZN(n409) );
  XOR2_X1 U491 ( .A(KEYINPUT8), .B(n409), .Z(n449) );
  NAND2_X1 U492 ( .A1(G221), .A2(n449), .ZN(n410) );
  XNOR2_X1 U493 ( .A(n411), .B(n410), .ZN(n417) );
  XOR2_X1 U494 ( .A(G110), .B(G137), .Z(n413) );
  XNOR2_X1 U495 ( .A(G119), .B(G128), .ZN(n412) );
  XNOR2_X1 U496 ( .A(n413), .B(n412), .ZN(n415) );
  XNOR2_X1 U497 ( .A(KEYINPUT10), .B(G140), .ZN(n427) );
  XOR2_X1 U498 ( .A(n427), .B(n426), .Z(n414) );
  XNOR2_X1 U499 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U500 ( .A(n417), .B(n416), .ZN(n695) );
  NOR2_X1 U501 ( .A1(n695), .A2(G902), .ZN(n421) );
  NAND2_X1 U502 ( .A1(G217), .A2(n418), .ZN(n419) );
  XNOR2_X2 U503 ( .A(n421), .B(n420), .ZN(n665) );
  INV_X1 U504 ( .A(n665), .ZN(n422) );
  AND2_X1 U505 ( .A1(n423), .A2(n422), .ZN(n463) );
  NAND2_X1 U506 ( .A1(n547), .A2(n463), .ZN(n424) );
  XNOR2_X1 U507 ( .A(n424), .B(KEYINPUT108), .ZN(n425) );
  INV_X1 U508 ( .A(n425), .ZN(n460) );
  XNOR2_X1 U509 ( .A(n427), .B(n426), .ZN(n711) );
  XOR2_X1 U510 ( .A(KEYINPUT11), .B(G131), .Z(n429) );
  XNOR2_X1 U511 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U512 ( .A(n711), .B(n430), .ZN(n438) );
  XOR2_X1 U513 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n433) );
  NAND2_X1 U514 ( .A1(G214), .A2(n431), .ZN(n432) );
  XNOR2_X1 U515 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U516 ( .A(n434), .B(KEYINPUT99), .Z(n436) );
  XNOR2_X1 U517 ( .A(G122), .B(G104), .ZN(n435) );
  XNOR2_X1 U518 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U519 ( .A(n438), .B(n437), .ZN(n596) );
  NOR2_X1 U520 ( .A1(G902), .A2(n596), .ZN(n442) );
  XOR2_X1 U521 ( .A(KEYINPUT13), .B(KEYINPUT101), .Z(n440) );
  XNOR2_X1 U522 ( .A(KEYINPUT100), .B(G475), .ZN(n439) );
  XNOR2_X1 U523 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U524 ( .A(n442), .B(n441), .ZN(n492) );
  INV_X1 U525 ( .A(n492), .ZN(n468) );
  XOR2_X1 U526 ( .A(G107), .B(G122), .Z(n444) );
  XNOR2_X1 U527 ( .A(G116), .B(G134), .ZN(n443) );
  XNOR2_X1 U528 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U529 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n446) );
  XNOR2_X1 U530 ( .A(KEYINPUT102), .B(KEYINPUT9), .ZN(n445) );
  XNOR2_X1 U531 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U532 ( .A(n448), .B(n447), .Z(n451) );
  NAND2_X1 U533 ( .A1(G217), .A2(n449), .ZN(n450) );
  XNOR2_X1 U534 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U535 ( .A(n453), .B(n452), .ZN(n591) );
  INV_X1 U536 ( .A(G902), .ZN(n454) );
  NAND2_X1 U537 ( .A1(n591), .A2(n454), .ZN(n455) );
  XNOR2_X1 U538 ( .A(n455), .B(G478), .ZN(n493) );
  NOR2_X1 U539 ( .A1(n468), .A2(n493), .ZN(n456) );
  XNOR2_X1 U540 ( .A(n456), .B(KEYINPUT104), .ZN(n639) );
  INV_X1 U541 ( .A(n639), .ZN(n637) );
  NAND2_X1 U542 ( .A1(n457), .A2(G214), .ZN(n458) );
  XOR2_X1 U543 ( .A(KEYINPUT93), .B(n458), .Z(n494) );
  NOR2_X1 U544 ( .A1(n478), .A2(n504), .ZN(n461) );
  XOR2_X1 U545 ( .A(KEYINPUT36), .B(n461), .Z(n462) );
  NOR2_X1 U546 ( .A1(n531), .A2(n462), .ZN(n644) );
  NAND2_X1 U547 ( .A1(n558), .A2(n463), .ZN(n464) );
  XNOR2_X1 U548 ( .A(n464), .B(KEYINPUT28), .ZN(n465) );
  NAND2_X1 U549 ( .A1(n509), .A2(n494), .ZN(n466) );
  NAND2_X1 U550 ( .A1(n496), .A2(n520), .ZN(n636) );
  NAND2_X1 U551 ( .A1(n636), .A2(KEYINPUT47), .ZN(n467) );
  XNOR2_X1 U552 ( .A(n467), .B(KEYINPUT84), .ZN(n482) );
  NAND2_X1 U553 ( .A1(n493), .A2(n468), .ZN(n632) );
  XNOR2_X1 U554 ( .A(KEYINPUT105), .B(n632), .ZN(n511) );
  NAND2_X1 U555 ( .A1(KEYINPUT47), .A2(n656), .ZN(n469) );
  XNOR2_X1 U556 ( .A(KEYINPUT85), .B(n469), .ZN(n479) );
  INV_X1 U557 ( .A(n471), .ZN(n557) );
  AND2_X1 U558 ( .A1(n557), .A2(n472), .ZN(n474) );
  NAND2_X1 U559 ( .A1(n666), .A2(n665), .ZN(n473) );
  XNOR2_X2 U560 ( .A(n473), .B(KEYINPUT67), .ZN(n663) );
  AND2_X1 U561 ( .A1(n474), .A2(n663), .ZN(n475) );
  NAND2_X1 U562 ( .A1(n476), .A2(n475), .ZN(n489) );
  NAND2_X1 U563 ( .A1(n493), .A2(n492), .ZN(n525) );
  OR2_X1 U564 ( .A1(n489), .A2(n525), .ZN(n477) );
  NOR2_X1 U565 ( .A1(n479), .A2(n635), .ZN(n480) );
  XNOR2_X1 U566 ( .A(n480), .B(KEYINPUT82), .ZN(n481) );
  AND2_X1 U567 ( .A1(n482), .A2(n481), .ZN(n487) );
  XNOR2_X1 U568 ( .A(n656), .B(KEYINPUT86), .ZN(n562) );
  INV_X1 U569 ( .A(n562), .ZN(n484) );
  NOR2_X1 U570 ( .A1(n636), .A2(KEYINPUT47), .ZN(n483) );
  NAND2_X1 U571 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U572 ( .A(KEYINPUT74), .B(n485), .ZN(n486) );
  NAND2_X1 U573 ( .A1(n487), .A2(n486), .ZN(n488) );
  NOR2_X1 U574 ( .A1(n644), .A2(n488), .ZN(n501) );
  OR2_X2 U575 ( .A1(n489), .A2(n651), .ZN(n490) );
  NOR2_X1 U576 ( .A1(n493), .A2(n492), .ZN(n654) );
  INV_X1 U577 ( .A(n494), .ZN(n652) );
  NAND2_X1 U578 ( .A1(n654), .A2(n658), .ZN(n495) );
  XNOR2_X1 U579 ( .A(n495), .B(KEYINPUT41), .ZN(n682) );
  NAND2_X1 U580 ( .A1(n682), .A2(n496), .ZN(n498) );
  NOR2_X1 U581 ( .A1(n726), .A2(n727), .ZN(n499) );
  XNOR2_X1 U582 ( .A(n499), .B(KEYINPUT46), .ZN(n500) );
  AND2_X2 U583 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U584 ( .A(n503), .B(n502), .ZN(n510) );
  XOR2_X1 U585 ( .A(KEYINPUT109), .B(n504), .Z(n505) );
  NOR2_X1 U586 ( .A1(n662), .A2(n505), .ZN(n507) );
  NOR2_X1 U587 ( .A1(n509), .A2(n508), .ZN(n648) );
  NOR2_X2 U588 ( .A1(n510), .A2(n648), .ZN(n582) );
  NAND2_X1 U589 ( .A1(n582), .A2(n646), .ZN(n715) );
  NAND2_X1 U590 ( .A1(n662), .A2(n663), .ZN(n554) );
  INV_X1 U591 ( .A(n554), .ZN(n512) );
  NAND2_X1 U592 ( .A1(n512), .A2(n547), .ZN(n513) );
  INV_X1 U593 ( .A(n514), .ZN(n518) );
  INV_X1 U594 ( .A(n515), .ZN(n516) );
  NOR2_X1 U595 ( .A1(G898), .A2(n722), .ZN(n700) );
  NAND2_X1 U596 ( .A1(n516), .A2(n700), .ZN(n517) );
  NAND2_X1 U597 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X2 U598 ( .A(n521), .B(KEYINPUT0), .ZN(n561) );
  NAND2_X1 U599 ( .A1(n683), .A2(n561), .ZN(n524) );
  XNOR2_X1 U600 ( .A(KEYINPUT76), .B(KEYINPUT34), .ZN(n522) );
  XNOR2_X1 U601 ( .A(n522), .B(KEYINPUT71), .ZN(n523) );
  XNOR2_X1 U602 ( .A(n524), .B(n523), .ZN(n527) );
  INV_X1 U603 ( .A(n525), .ZN(n526) );
  NAND2_X1 U604 ( .A1(n527), .A2(n526), .ZN(n529) );
  INV_X1 U605 ( .A(KEYINPUT35), .ZN(n528) );
  XNOR2_X1 U606 ( .A(n529), .B(n528), .ZN(n615) );
  OR2_X1 U607 ( .A1(n547), .A2(n665), .ZN(n530) );
  OR2_X1 U608 ( .A1(n531), .A2(n530), .ZN(n533) );
  INV_X1 U609 ( .A(KEYINPUT78), .ZN(n532) );
  XNOR2_X1 U610 ( .A(n533), .B(n532), .ZN(n536) );
  AND2_X1 U611 ( .A1(n666), .A2(n654), .ZN(n534) );
  NAND2_X1 U612 ( .A1(n561), .A2(n534), .ZN(n535) );
  XNOR2_X1 U613 ( .A(n535), .B(KEYINPUT22), .ZN(n548) );
  INV_X1 U614 ( .A(n548), .ZN(n540) );
  NAND2_X1 U615 ( .A1(n536), .A2(n540), .ZN(n539) );
  INV_X1 U616 ( .A(KEYINPUT77), .ZN(n537) );
  XNOR2_X1 U617 ( .A(n537), .B(KEYINPUT32), .ZN(n538) );
  INV_X1 U618 ( .A(n540), .ZN(n543) );
  INV_X1 U619 ( .A(n662), .ZN(n550) );
  NOR2_X1 U620 ( .A1(n558), .A2(n665), .ZN(n541) );
  NAND2_X1 U621 ( .A1(n550), .A2(n541), .ZN(n542) );
  NOR2_X1 U622 ( .A1(n543), .A2(n542), .ZN(n630) );
  NOR2_X1 U623 ( .A1(n630), .A2(KEYINPUT44), .ZN(n544) );
  NAND2_X1 U624 ( .A1(n614), .A2(n544), .ZN(n545) );
  NAND2_X1 U625 ( .A1(n545), .A2(KEYINPUT88), .ZN(n546) );
  NAND2_X1 U626 ( .A1(n615), .A2(n546), .ZN(n566) );
  NOR2_X1 U627 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U628 ( .A(n549), .B(KEYINPUT87), .ZN(n552) );
  NAND2_X1 U629 ( .A1(n550), .A2(n665), .ZN(n551) );
  NOR2_X1 U630 ( .A1(n554), .A2(n669), .ZN(n672) );
  NAND2_X1 U631 ( .A1(n672), .A2(n561), .ZN(n556) );
  XOR2_X1 U632 ( .A(KEYINPUT97), .B(KEYINPUT31), .Z(n555) );
  XNOR2_X1 U633 ( .A(n556), .B(n555), .ZN(n642) );
  NAND2_X1 U634 ( .A1(n557), .A2(n663), .ZN(n559) );
  NOR2_X1 U635 ( .A1(n559), .A2(n558), .ZN(n560) );
  AND2_X1 U636 ( .A1(n561), .A2(n560), .ZN(n626) );
  NOR2_X1 U637 ( .A1(n642), .A2(n626), .ZN(n563) );
  NOR2_X1 U638 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U639 ( .A1(n728), .A2(n564), .ZN(n565) );
  AND2_X1 U640 ( .A1(n566), .A2(n565), .ZN(n577) );
  INV_X1 U641 ( .A(n615), .ZN(n567) );
  NAND2_X1 U642 ( .A1(n567), .A2(KEYINPUT88), .ZN(n572) );
  INV_X1 U643 ( .A(n614), .ZN(n570) );
  INV_X1 U644 ( .A(n630), .ZN(n568) );
  NAND2_X1 U645 ( .A1(n568), .A2(KEYINPUT44), .ZN(n569) );
  NOR2_X1 U646 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U647 ( .A1(n572), .A2(n571), .ZN(n575) );
  INV_X1 U648 ( .A(KEYINPUT44), .ZN(n573) );
  NAND2_X1 U649 ( .A1(n573), .A2(KEYINPUT88), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U651 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U652 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n578) );
  XNOR2_X2 U653 ( .A(n579), .B(n578), .ZN(n702) );
  NAND2_X1 U654 ( .A1(n580), .A2(n702), .ZN(n581) );
  INV_X1 U655 ( .A(KEYINPUT2), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n581), .A2(n583), .ZN(n589) );
  INV_X1 U657 ( .A(n582), .ZN(n586) );
  XOR2_X1 U658 ( .A(n646), .B(KEYINPUT81), .Z(n584) );
  NAND2_X1 U659 ( .A1(n584), .A2(KEYINPUT2), .ZN(n585) );
  NOR2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n587), .A2(n702), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n650) );
  NOR2_X4 U663 ( .A1(n650), .A2(n590), .ZN(n616) );
  NAND2_X1 U664 ( .A1(n693), .A2(G478), .ZN(n592) );
  INV_X1 U665 ( .A(G952), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n616), .A2(G475), .ZN(n598) );
  XOR2_X1 U667 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n595) );
  XNOR2_X1 U668 ( .A(n600), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U669 ( .A1(n616), .A2(G210), .ZN(n605) );
  XOR2_X1 U670 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n603) );
  XNOR2_X1 U671 ( .A(n601), .B(KEYINPUT83), .ZN(n602) );
  XNOR2_X1 U672 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U673 ( .A(n605), .B(n604), .ZN(n606) );
  NOR2_X2 U674 ( .A1(n606), .A2(n697), .ZN(n607) );
  XNOR2_X1 U675 ( .A(n607), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U676 ( .A1(n616), .A2(G469), .ZN(n610) );
  XOR2_X1 U677 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n608) );
  XNOR2_X1 U678 ( .A(n610), .B(n352), .ZN(n612) );
  NAND2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U680 ( .A(n613), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U681 ( .A(n614), .B(G119), .ZN(G21) );
  XNOR2_X1 U682 ( .A(n615), .B(G122), .ZN(G24) );
  NAND2_X1 U683 ( .A1(n616), .A2(G472), .ZN(n621) );
  XNOR2_X1 U684 ( .A(KEYINPUT90), .B(KEYINPUT112), .ZN(n617) );
  XNOR2_X1 U685 ( .A(n617), .B(KEYINPUT62), .ZN(n618) );
  XNOR2_X1 U686 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U687 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X2 U688 ( .A1(n622), .A2(n697), .ZN(n624) );
  XNOR2_X1 U689 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n623) );
  XNOR2_X1 U690 ( .A(n624), .B(n623), .ZN(G57) );
  NAND2_X1 U691 ( .A1(n639), .A2(n626), .ZN(n625) );
  XNOR2_X1 U692 ( .A(n625), .B(G104), .ZN(G6) );
  XOR2_X1 U693 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n628) );
  INV_X1 U694 ( .A(n632), .ZN(n641) );
  NAND2_X1 U695 ( .A1(n626), .A2(n641), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U697 ( .A(G107), .B(n629), .ZN(G9) );
  XNOR2_X1 U698 ( .A(n630), .B(G110), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n631), .B(KEYINPUT113), .ZN(G12) );
  NOR2_X1 U700 ( .A1(n636), .A2(n632), .ZN(n634) );
  XNOR2_X1 U701 ( .A(G128), .B(KEYINPUT29), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(G30) );
  XOR2_X1 U703 ( .A(G143), .B(n635), .Z(G45) );
  NOR2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U705 ( .A(G146), .B(n638), .Z(G48) );
  NAND2_X1 U706 ( .A1(n639), .A2(n642), .ZN(n640) );
  XNOR2_X1 U707 ( .A(n640), .B(G113), .ZN(G15) );
  NAND2_X1 U708 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U709 ( .A(n643), .B(G116), .ZN(G18) );
  XNOR2_X1 U710 ( .A(n644), .B(G125), .ZN(n645) );
  XNOR2_X1 U711 ( .A(n645), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U712 ( .A(G134), .B(KEYINPUT114), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n647), .B(n646), .ZN(G36) );
  XNOR2_X1 U714 ( .A(G140), .B(n648), .ZN(n649) );
  XNOR2_X1 U715 ( .A(n649), .B(KEYINPUT115), .ZN(G42) );
  XOR2_X1 U716 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n692) );
  BUF_X1 U717 ( .A(n650), .Z(n688) );
  NAND2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U719 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U720 ( .A(n655), .B(KEYINPUT116), .ZN(n660) );
  INV_X1 U721 ( .A(n656), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U723 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U724 ( .A1(n683), .A2(n661), .ZN(n677) );
  NOR2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U726 ( .A(n664), .B(KEYINPUT50), .ZN(n671) );
  NOR2_X1 U727 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U728 ( .A(n667), .B(KEYINPUT49), .ZN(n668) );
  NAND2_X1 U729 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U730 ( .A1(n671), .A2(n670), .ZN(n673) );
  NOR2_X1 U731 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U732 ( .A(KEYINPUT51), .B(n674), .ZN(n675) );
  NAND2_X1 U733 ( .A1(n682), .A2(n675), .ZN(n676) );
  NAND2_X1 U734 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U735 ( .A(KEYINPUT52), .B(n678), .Z(n679) );
  NOR2_X1 U736 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U737 ( .A(KEYINPUT117), .B(n681), .Z(n686) );
  NAND2_X1 U738 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U739 ( .A(KEYINPUT118), .B(n684), .Z(n685) );
  NOR2_X1 U740 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U741 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U742 ( .A(n689), .B(KEYINPUT119), .ZN(n690) );
  NAND2_X1 U743 ( .A1(n690), .A2(n722), .ZN(n691) );
  XNOR2_X1 U744 ( .A(n692), .B(n691), .ZN(G75) );
  NAND2_X1 U745 ( .A1(n693), .A2(G217), .ZN(n694) );
  XNOR2_X1 U746 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U747 ( .A1(n697), .A2(n696), .ZN(G66) );
  XNOR2_X1 U748 ( .A(G101), .B(n698), .ZN(n699) );
  XNOR2_X1 U749 ( .A(n699), .B(KEYINPUT124), .ZN(n701) );
  NOR2_X1 U750 ( .A1(n701), .A2(n700), .ZN(n709) );
  NAND2_X1 U751 ( .A1(n702), .A2(n722), .ZN(n703) );
  XOR2_X1 U752 ( .A(KEYINPUT123), .B(n703), .Z(n707) );
  NAND2_X1 U753 ( .A1(G953), .A2(G224), .ZN(n704) );
  XNOR2_X1 U754 ( .A(KEYINPUT61), .B(n704), .ZN(n705) );
  NAND2_X1 U755 ( .A1(n705), .A2(G898), .ZN(n706) );
  NAND2_X1 U756 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U757 ( .A(n709), .B(n708), .ZN(G69) );
  INV_X1 U758 ( .A(KEYINPUT95), .ZN(n710) );
  XNOR2_X1 U759 ( .A(n711), .B(n710), .ZN(n713) );
  XNOR2_X1 U760 ( .A(n713), .B(n712), .ZN(n717) );
  INV_X1 U761 ( .A(n717), .ZN(n714) );
  XNOR2_X1 U762 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U763 ( .A1(n716), .A2(n722), .ZN(n725) );
  XNOR2_X1 U764 ( .A(n717), .B(KEYINPUT125), .ZN(n718) );
  XNOR2_X1 U765 ( .A(G227), .B(n718), .ZN(n719) );
  NAND2_X1 U766 ( .A1(G900), .A2(n719), .ZN(n720) );
  XOR2_X1 U767 ( .A(KEYINPUT126), .B(n720), .Z(n721) );
  NOR2_X1 U768 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U769 ( .A(KEYINPUT127), .B(n723), .ZN(n724) );
  NAND2_X1 U770 ( .A1(n725), .A2(n724), .ZN(G72) );
  XOR2_X1 U771 ( .A(n726), .B(G131), .Z(G33) );
  XOR2_X1 U772 ( .A(n727), .B(G137), .Z(G39) );
  XOR2_X1 U773 ( .A(G101), .B(n728), .Z(G3) );
endmodule

