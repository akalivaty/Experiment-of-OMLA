//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  OR4_X1    g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n460), .B2(new_n461), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(KEYINPUT68), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n468), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n475), .B2(G2105), .ZN(G160));
  AOI21_X1  g051(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n459), .B1(new_n470), .B2(new_n471), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n468), .A2(new_n472), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n491), .B2(new_n494), .ZN(G164));
  NOR2_X1   g070(.A1(KEYINPUT6), .A2(G651), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G88), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n502), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n499), .A2(new_n500), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n506), .A2(new_n510), .ZN(G166));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  INV_X1    g088(.A(G51), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n505), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n504), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G168));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n497), .B2(new_n498), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G52), .ZN(new_n525));
  INV_X1    g100(.A(new_n501), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT69), .B(G90), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n509), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(G171));
  NAND2_X1  g106(.A1(G68), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G56), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n518), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n501), .A2(G81), .B1(new_n524), .B2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n535), .A2(new_n536), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n543));
  XOR2_X1   g118(.A(new_n543), .B(KEYINPUT71), .Z(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(G78), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n554), .B(new_n555), .C1(new_n505), .C2(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n556), .B1(KEYINPUT72), .B2(KEYINPUT9), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n524), .B(new_n558), .C1(KEYINPUT72), .C2(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n501), .A2(G91), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n553), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n501), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n524), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  INV_X1    g144(.A(G61), .ZN(new_n570));
  INV_X1    g145(.A(G73), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n518), .A2(new_n570), .B1(new_n571), .B2(new_n523), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n501), .B2(G86), .ZN(new_n573));
  AND2_X1   g148(.A1(KEYINPUT6), .A2(G651), .ZN(new_n574));
  OAI211_X1 g149(.A(G48), .B(G543), .C1(new_n574), .C2(new_n496), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n504), .A2(KEYINPUT74), .A3(G48), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT75), .ZN(G305));
  NAND2_X1  g156(.A1(new_n501), .A2(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n505), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n509), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NOR2_X1   g164(.A1(G171), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT76), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n507), .A2(new_n504), .A3(G92), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(KEYINPUT10), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n593), .A2(new_n594), .B1(G54), .B2(new_n524), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n549), .B2(new_n550), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT77), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G321));
  NOR2_X1   g179(.A1(G286), .A2(new_n589), .ZN(new_n605));
  XNOR2_X1  g180(.A(G299), .B(KEYINPUT78), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n589), .ZN(G297));
  AOI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n589), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g189(.A1(new_n468), .A2(new_n472), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n464), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n479), .A2(G123), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT79), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n477), .A2(G135), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n459), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n620), .A2(new_n621), .A3(new_n628), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(G14), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n641), .ZN(G401));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n646), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT81), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n647), .A2(new_n648), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1971), .B(G1976), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT82), .ZN(new_n669));
  OR3_X1    g244(.A1(new_n661), .A2(new_n664), .A3(new_n667), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n677), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n681), .B1(new_n678), .B2(new_n682), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(G229));
  MUX2_X1   g260(.A(G6), .B(G305), .S(G16), .Z(new_n686));
  XOR2_X1   g261(.A(KEYINPUT32), .B(G1981), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT87), .B(G16), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(G22), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n693), .ZN(new_n695));
  INV_X1    g270(.A(G1971), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT33), .B(G1976), .Z(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  NAND4_X1  g278(.A1(new_n690), .A2(new_n691), .A3(new_n697), .A4(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n587), .A2(new_n692), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G24), .B2(new_n692), .ZN(new_n708));
  OAI21_X1  g283(.A(KEYINPUT89), .B1(new_n708), .B2(new_n674), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n479), .A2(G119), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT86), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n712));
  INV_X1    g287(.A(G107), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(G2105), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n477), .B2(G131), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT85), .B(G29), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G25), .B(new_n716), .S(new_n718), .Z(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n719), .B(new_n721), .ZN(new_n722));
  AOI211_X1 g297(.A(new_n709), .B(new_n722), .C1(new_n674), .C2(new_n708), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n705), .A2(new_n706), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n705), .A2(KEYINPUT36), .A3(new_n706), .A4(new_n723), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT24), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(G34), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(G34), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n717), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G160), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G2084), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n602), .A2(new_n698), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G4), .B2(new_n698), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n736), .B1(new_n739), .B2(G1348), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n734), .A2(new_n735), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n718), .A2(G35), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n718), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2090), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n745), .B2(new_n744), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n717), .A2(G27), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT96), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n494), .A2(new_n491), .ZN(new_n750));
  INV_X1    g325(.A(new_n489), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n749), .B1(new_n752), .B2(new_n718), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G1348), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n740), .A2(new_n747), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n692), .A2(G20), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT23), .Z(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G299), .B2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT99), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT98), .B(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n733), .A2(G32), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n479), .A2(G129), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n464), .A2(G105), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n477), .A2(G141), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OR3_X1    g347(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n765), .B1(new_n774), .B2(new_n733), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT27), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1996), .ZN(new_n777));
  NOR2_X1   g352(.A1(G171), .A2(new_n698), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G5), .B2(new_n698), .ZN(new_n779));
  INV_X1    g354(.A(G1961), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G11), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT30), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n784), .A2(G28), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n733), .B1(new_n784), .B2(G28), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n783), .B1(new_n785), .B2(new_n786), .C1(new_n627), .C2(new_n717), .ZN(new_n787));
  OR3_X1    g362(.A1(new_n781), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n693), .A2(G19), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n541), .B2(new_n693), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1341), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n698), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n698), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1966), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n717), .A2(G26), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT28), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n477), .A2(G140), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n479), .A2(G128), .ZN(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n733), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2067), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n788), .A2(new_n791), .A3(new_n794), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n758), .A2(new_n764), .A3(new_n777), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G29), .A2(G33), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT90), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n615), .A2(G127), .ZN(new_n809));
  INV_X1    g384(.A(G115), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n463), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT92), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n809), .B(KEYINPUT92), .C1(new_n810), .C2(new_n463), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n813), .A2(G2105), .A3(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT93), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT93), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT25), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n477), .A2(G139), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT91), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n816), .A2(new_n817), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n808), .B1(new_n823), .B2(new_n733), .ZN(new_n824));
  INV_X1    g399(.A(G2072), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT95), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n825), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT94), .Z(new_n829));
  NOR3_X1   g404(.A1(new_n806), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n726), .A2(new_n727), .A3(new_n830), .ZN(G150));
  INV_X1    g406(.A(G150), .ZN(G311));
  NAND2_X1  g407(.A1(new_n602), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(new_n509), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n501), .A2(G93), .B1(new_n524), .B2(G55), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n541), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n834), .B(new_n839), .Z(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n838), .A2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  XNOR2_X1  g422(.A(new_n802), .B(G164), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n477), .A2(G142), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n479), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n459), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n848), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n823), .B(new_n774), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n716), .B(KEYINPUT100), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n617), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n857), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(new_n854), .A3(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G160), .B(G162), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n627), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n861), .A2(new_n867), .A3(new_n862), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT40), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n862), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n865), .B1(new_n870), .B2(new_n860), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  AND4_X1   g447(.A1(KEYINPUT40), .A2(new_n871), .A3(new_n868), .A4(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n869), .A2(new_n873), .ZN(G395));
  XOR2_X1   g449(.A(new_n601), .B(G299), .Z(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT41), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n839), .B(new_n611), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n875), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n876), .A2(new_n882), .A3(new_n878), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(G305), .B(G290), .ZN(new_n885));
  XNOR2_X1  g460(.A(G166), .B(new_n700), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n883), .A2(new_n881), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n880), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G868), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n838), .A2(G868), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n589), .B1(new_n890), .B2(new_n892), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT102), .B1(new_n899), .B2(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(G295));
  NAND2_X1  g476(.A1(new_n894), .A2(new_n897), .ZN(G331));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n839), .B(G301), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(G168), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n875), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n904), .A2(G168), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(G168), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n876), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n887), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n906), .A2(new_n909), .A3(new_n887), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n903), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n910), .A2(new_n911), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n919), .A2(new_n872), .A3(new_n914), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  OAI211_X1 g496(.A(KEYINPUT44), .B(new_n918), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n922), .ZN(G397));
  NAND2_X1  g498(.A1(G303), .A2(G8), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT55), .ZN(new_n925));
  INV_X1    g500(.A(G2090), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT50), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n752), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n459), .B1(new_n473), .B2(new_n474), .ZN(new_n931));
  INV_X1    g506(.A(G40), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n931), .A2(new_n932), .A3(new_n466), .ZN(new_n933));
  AND4_X1   g508(.A1(new_n926), .A2(new_n929), .A3(new_n930), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n752), .A2(new_n928), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g512(.A(KEYINPUT105), .B(G1384), .Z(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n750), .B2(new_n751), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT110), .B1(new_n939), .B2(KEYINPUT45), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n941));
  NOR4_X1   g516(.A1(G164), .A2(new_n941), .A3(new_n936), .A4(new_n938), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n933), .B(new_n937), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n934), .B1(new_n943), .B2(new_n696), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n945));
  OAI21_X1  g520(.A(G8), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n929), .A2(new_n930), .A3(new_n933), .A4(new_n926), .ZN(new_n947));
  AOI21_X1  g522(.A(G1384), .B1(new_n750), .B2(new_n751), .ZN(new_n948));
  OAI211_X1 g523(.A(G40), .B(G160), .C1(new_n948), .C2(KEYINPUT45), .ZN(new_n949));
  INV_X1    g524(.A(new_n938), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n752), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n941), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n939), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n947), .B(new_n945), .C1(new_n954), .C2(G1971), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n925), .B1(new_n946), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n958), .A2(G2084), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n948), .A2(KEYINPUT45), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n937), .A2(new_n933), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1966), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n964), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n957), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n952), .A2(new_n953), .ZN(new_n968));
  INV_X1    g543(.A(new_n949), .ZN(new_n969));
  AOI21_X1  g544(.A(G1971), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT111), .B1(new_n970), .B2(new_n934), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n924), .B(KEYINPUT55), .Z(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(G8), .A3(new_n972), .A4(new_n955), .ZN(new_n973));
  INV_X1    g548(.A(G1976), .ZN(new_n974));
  NOR2_X1   g549(.A1(G288), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n977), .B(new_n978), .C1(new_n933), .C2(new_n948), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n948), .A2(G160), .A3(G40), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT112), .B1(new_n980), .B2(G8), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n976), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT113), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n475), .A2(G2105), .ZN(new_n984));
  INV_X1    g559(.A(new_n466), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(G40), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(G8), .B1(new_n986), .B2(new_n935), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n977), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n980), .A2(KEYINPUT112), .A3(G8), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n976), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n983), .A2(new_n992), .A3(KEYINPUT52), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n501), .A2(G86), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n570), .B1(new_n499), .B2(new_n500), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n571), .A2(new_n523), .ZN(new_n996));
  OAI21_X1  g571(.A(G651), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n579), .A2(new_n672), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n573), .A2(KEYINPUT114), .A3(new_n672), .A4(new_n579), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n580), .A2(G1981), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1002), .A2(KEYINPUT49), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT49), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n975), .B1(new_n988), .B2(new_n989), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(G288), .B2(new_n974), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n990), .A2(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n973), .A2(new_n993), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT116), .B1(new_n967), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT63), .ZN(new_n1012));
  OAI21_X1  g587(.A(G8), .B1(new_n970), .B2(new_n934), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n925), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n973), .A2(new_n1014), .A3(new_n993), .A4(new_n1009), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n964), .A2(G8), .A3(G168), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n971), .A2(G8), .A3(new_n955), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n965), .B1(new_n1018), .B2(new_n925), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n976), .B(new_n1008), .C1(new_n979), .C2(new_n981), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1005), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1002), .A2(KEYINPUT49), .A3(new_n1003), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n979), .A2(new_n981), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n982), .B2(KEYINPUT113), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1025), .B1(new_n992), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1019), .A2(new_n1028), .A3(new_n1029), .A4(new_n973), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1011), .A2(new_n1017), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n700), .A2(new_n974), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1002), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1024), .B1(new_n1034), .B2(KEYINPUT115), .ZN(new_n1036));
  INV_X1    g611(.A(new_n973), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1035), .A2(new_n1036), .B1(new_n1028), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1031), .A2(KEYINPUT117), .A3(new_n1038), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n1043));
  INV_X1    g618(.A(G1996), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n968), .A2(new_n1044), .A3(new_n969), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n980), .A2(KEYINPUT118), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n933), .A2(new_n1047), .A3(new_n948), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT58), .B(G1341), .Z(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1043), .B1(new_n1051), .B2(new_n541), .ZN(new_n1052));
  INV_X1    g627(.A(new_n541), .ZN(new_n1053));
  AOI211_X1 g628(.A(KEYINPUT59), .B(new_n1053), .C1(new_n1045), .C2(new_n1050), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n1056));
  AOI21_X1  g631(.A(G2067), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n958), .A2(new_n756), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n601), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1059), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n602), .B1(new_n1061), .B2(new_n1057), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1056), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NOR4_X1   g638(.A1(new_n1061), .A2(new_n1057), .A3(KEYINPUT60), .A4(new_n601), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1055), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT61), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n968), .A2(new_n969), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n553), .B2(new_n561), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1956), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n958), .A2(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1068), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1066), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT120), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n1066), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1068), .A2(new_n1074), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT119), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1072), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1068), .A2(new_n1085), .A3(new_n1074), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1068), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1068), .A2(new_n1072), .A3(KEYINPUT121), .A4(new_n1074), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(KEYINPUT61), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT122), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1066), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1091), .A4(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1065), .A2(new_n1081), .A3(new_n1093), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1062), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1088), .B1(new_n1087), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1015), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n959), .A2(new_n963), .A3(G168), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G8), .ZN(new_n1104));
  AOI21_X1  g679(.A(G168), .B1(new_n959), .B2(new_n963), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT51), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1107), .A3(G8), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n954), .A2(new_n754), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1111), .A2(new_n1112), .B1(new_n780), .B2(new_n958), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT123), .B1(new_n961), .B2(G2078), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n969), .A2(new_n1115), .A3(new_n754), .A4(new_n960), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(KEYINPUT53), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(G301), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1112), .B1(new_n943), .B2(G2078), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n958), .A2(new_n780), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1112), .B(G2078), .C1(new_n986), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n752), .A2(new_n950), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT106), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT45), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n939), .A2(KEYINPUT106), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n933), .A2(KEYINPUT124), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1122), .A2(new_n1127), .A3(new_n968), .A4(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1119), .A2(new_n1120), .A3(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1130), .A2(G171), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1110), .B1(new_n1118), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1102), .A2(new_n1109), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1110), .B1(new_n1130), .B2(G171), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1113), .A2(G301), .A3(new_n1117), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1135), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1101), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1106), .A2(new_n1143), .A3(new_n1108), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1118), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1145), .B2(new_n1015), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1109), .A2(KEYINPUT62), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1102), .A2(KEYINPUT126), .A3(new_n1118), .A4(new_n1144), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1041), .A2(new_n1042), .A3(new_n1141), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1125), .A2(new_n933), .A3(new_n1126), .ZN(new_n1151));
  INV_X1    g726(.A(G2067), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n801), .B(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT108), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1151), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n773), .B(G1996), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n716), .A2(new_n721), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n720), .B1(new_n711), .B2(new_n715), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n587), .A2(new_n674), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT107), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n674), .B2(new_n587), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1156), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT109), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1150), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n802), .A2(new_n1152), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1151), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1156), .A2(new_n1044), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT46), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT127), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1151), .B1(new_n774), .B2(new_n1153), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT47), .Z(new_n1180));
  NOR2_X1   g755(.A1(new_n1164), .A2(new_n1151), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT48), .Z(new_n1182));
  AOI211_X1 g757(.A(new_n1172), .B(new_n1180), .C1(new_n1162), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1169), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g759(.A1(new_n871), .A2(new_n868), .A3(new_n872), .ZN(new_n1186));
  OR3_X1    g760(.A1(G401), .A2(new_n457), .A3(G227), .ZN(new_n1187));
  NOR3_X1   g761(.A1(new_n683), .A2(new_n684), .A3(new_n1187), .ZN(new_n1188));
  OAI211_X1 g762(.A(new_n1186), .B(new_n1188), .C1(new_n915), .C2(new_n916), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


