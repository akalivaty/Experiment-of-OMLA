//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT64), .B1(new_n190), .B2(G143), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n192), .A3(G146), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n195), .A2(new_n197), .B1(G143), .B2(new_n190), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n188), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n194), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT0), .B(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n195), .A2(new_n197), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(new_n191), .ZN(new_n204));
  AND4_X1   g018(.A1(KEYINPUT0), .A2(new_n191), .A3(new_n193), .A4(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(G125), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n208));
  INV_X1    g022(.A(G224), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G953), .ZN(new_n210));
  INV_X1    g024(.A(G953), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT84), .A3(G224), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g027(.A(new_n213), .B(KEYINPUT83), .Z(new_n214));
  XNOR2_X1  g028(.A(new_n207), .B(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT76), .A2(G104), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT3), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT76), .A2(G104), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT3), .A2(G107), .ZN(new_n221));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G107), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(G101), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G107), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(G104), .B2(new_n218), .ZN(new_n227));
  OR2_X1    g041(.A1(KEYINPUT76), .A2(G104), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n222), .A2(new_n228), .A3(new_n216), .ZN(new_n229));
  INV_X1    g043(.A(G101), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n225), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT67), .B1(new_n233), .B2(G116), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n236), .A2(G119), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n242), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n238), .A3(new_n240), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n227), .A2(new_n229), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G101), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n232), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G107), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n228), .A2(new_n251), .A3(new_n216), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n230), .B1(G104), .B2(G107), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n231), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G113), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n239), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n241), .B2(new_n257), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(new_n245), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n250), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n250), .A2(new_n260), .A3(KEYINPUT82), .ZN(new_n264));
  XNOR2_X1  g078(.A(G110), .B(G122), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n250), .A2(new_n260), .A3(new_n265), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT6), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n265), .B1(new_n261), .B2(new_n262), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT6), .A3(new_n264), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n215), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G210), .B1(G237), .B2(G902), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n274), .B(KEYINPUT88), .Z(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(KEYINPUT87), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT86), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT7), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n201), .A2(new_n206), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n210), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n282), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n201), .A2(new_n206), .A3(new_n284), .A4(new_n280), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n268), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n265), .B(KEYINPUT8), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n258), .B1(new_n241), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(new_n245), .A3(new_n231), .A4(new_n254), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n291), .A2(KEYINPUT85), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n259), .A2(new_n245), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n231), .A2(new_n254), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n291), .A2(KEYINPUT85), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n288), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n278), .B1(new_n286), .B2(new_n296), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n273), .A2(new_n277), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n277), .ZN(new_n299));
  INV_X1    g113(.A(new_n215), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n271), .A2(KEYINPUT6), .A3(new_n264), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n271), .A2(new_n264), .B1(KEYINPUT6), .B2(new_n268), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n297), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n299), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n187), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G113), .B(G122), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(new_n223), .ZN(new_n308));
  NOR2_X1   g122(.A1(G237), .A2(G953), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n309), .A2(G143), .A3(G214), .ZN(new_n310));
  AOI21_X1  g124(.A(G143), .B1(new_n309), .B2(G214), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT18), .A2(G131), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G146), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n190), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n312), .A2(new_n313), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G237), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n211), .A3(G214), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n192), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n309), .A2(G143), .A3(G214), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT89), .ZN(new_n328));
  INV_X1    g142(.A(new_n313), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n328), .B1(new_n327), .B2(new_n329), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n322), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT16), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n316), .A2(KEYINPUT16), .A3(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G146), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT19), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n315), .B(new_n317), .C1(KEYINPUT90), .C2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n320), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G131), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n325), .B2(new_n326), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n310), .A2(new_n311), .A3(G131), .ZN(new_n343));
  OAI221_X1 g157(.A(new_n336), .B1(new_n340), .B2(G146), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n308), .B1(new_n333), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n319), .A2(new_n321), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n327), .B2(new_n329), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT89), .B1(new_n312), .B2(new_n313), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n330), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n334), .A2(new_n335), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n190), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT17), .B(G131), .C1(new_n310), .C2(new_n311), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n336), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n343), .A2(new_n342), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT17), .ZN(new_n355));
  AOI22_X1  g169(.A1(KEYINPUT92), .A2(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n351), .A2(new_n352), .A3(new_n357), .A4(new_n336), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n349), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n308), .B(KEYINPUT91), .Z(new_n360));
  AOI21_X1  g174(.A(new_n345), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(G475), .A2(G902), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT20), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n353), .A2(KEYINPUT92), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n354), .A2(new_n355), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n358), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n360), .A3(new_n333), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n333), .A2(new_n344), .ZN(new_n369));
  INV_X1    g183(.A(new_n308), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n362), .ZN(new_n374));
  INV_X1    g188(.A(new_n368), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n308), .B1(new_n367), .B2(new_n333), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n278), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n364), .A2(new_n374), .B1(new_n377), .B2(G475), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n211), .A2(G952), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(G234), .B2(G237), .ZN(new_n380));
  NAND2_X1  g194(.A1(G234), .A2(G237), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(G902), .A3(G953), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT94), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT21), .B(G898), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT93), .B1(new_n192), .B2(G128), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n188), .A3(G143), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n192), .A2(G128), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n192), .A2(KEYINPUT13), .A3(G128), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G134), .ZN(new_n396));
  INV_X1    g210(.A(G122), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G116), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n236), .A2(G122), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(G107), .ZN(new_n401));
  INV_X1    g215(.A(G134), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n390), .A2(new_n402), .A3(new_n391), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n396), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n251), .B1(new_n398), .B2(KEYINPUT14), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n405), .A2(new_n400), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n400), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n390), .A2(new_n402), .A3(new_n391), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n402), .B1(new_n390), .B2(new_n391), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n406), .B(new_n407), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT9), .B(G234), .ZN(new_n411));
  INV_X1    g225(.A(G217), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n411), .A2(new_n412), .A3(G953), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n404), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n404), .B2(new_n410), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n278), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G478), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT15), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n416), .B(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n378), .A2(new_n386), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n306), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT68), .B1(new_n204), .B2(new_n205), .ZN(new_n424));
  XNOR2_X1  g238(.A(G143), .B(G146), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT0), .A3(G128), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT68), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(new_n198), .C2(new_n202), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT11), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n402), .B2(G137), .ZN(new_n430));
  INV_X1    g244(.A(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT11), .A3(G134), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n402), .A2(G137), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G131), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n430), .A2(new_n432), .A3(new_n341), .A4(new_n433), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n424), .A2(new_n428), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n246), .ZN(new_n439));
  INV_X1    g253(.A(new_n433), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n402), .A2(G137), .ZN(new_n441));
  OAI21_X1  g255(.A(G131), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n200), .A2(new_n436), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT28), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT28), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n438), .A2(new_n446), .A3(new_n439), .A4(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT65), .B1(new_n204), .B2(new_n205), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT65), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n426), .B(new_n450), .C1(new_n198), .C2(new_n202), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n451), .A3(new_n437), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT66), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT66), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n454), .A3(new_n451), .A4(new_n437), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n455), .A3(new_n443), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n246), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n309), .A2(G210), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT27), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT26), .B(G101), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n461), .B(KEYINPUT69), .Z(new_n462));
  NAND3_X1  g276(.A1(new_n448), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n444), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n456), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n438), .A2(KEYINPUT30), .A3(new_n443), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n246), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n423), .B(new_n463), .C1(new_n470), .C2(new_n461), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n439), .B1(new_n438), .B2(new_n443), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n448), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n461), .A2(KEYINPUT29), .ZN(new_n475));
  OAI211_X1 g289(.A(KEYINPUT71), .B(new_n278), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT71), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n472), .B(new_n475), .C1(new_n445), .C2(new_n447), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(G902), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G472), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n462), .B1(new_n448), .B2(new_n457), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n466), .A2(new_n469), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n444), .A2(new_n461), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT31), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n200), .A2(new_n436), .A3(new_n442), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n452), .B2(KEYINPUT66), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT30), .B1(new_n488), .B2(new_n455), .ZN(new_n489));
  OAI211_X1 g303(.A(KEYINPUT31), .B(new_n485), .C1(new_n489), .C2(new_n468), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n483), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(G472), .A2(G902), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(KEYINPUT32), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n485), .B1(new_n489), .B2(new_n468), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT31), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n482), .B1(new_n498), .B2(new_n490), .ZN(new_n499));
  INV_X1    g313(.A(new_n493), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n481), .A2(new_n494), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n351), .A2(new_n336), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n233), .A2(G128), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n188), .A2(G119), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT24), .B(G110), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT23), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n233), .B2(G128), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n504), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n508), .B1(G110), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT22), .B(G137), .ZN(new_n515));
  NAND2_X1  g329(.A1(G221), .A2(G234), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT73), .B1(new_n516), .B2(G953), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT73), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n518), .A2(new_n211), .A3(G221), .A4(G234), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n515), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT72), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n318), .A2(G146), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n316), .A2(KEYINPUT16), .A3(G140), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n525), .B1(new_n527), .B2(G146), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n506), .A2(new_n507), .ZN(new_n529));
  INV_X1    g343(.A(G110), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n510), .A2(new_n511), .A3(new_n530), .A4(new_n504), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n524), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  AND4_X1   g347(.A1(new_n524), .A2(new_n532), .A3(new_n336), .A4(new_n321), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n514), .B(new_n523), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n336), .A3(new_n321), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT72), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n528), .A2(new_n524), .A3(new_n532), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n537), .A2(new_n538), .B1(new_n503), .B2(new_n513), .ZN(new_n539));
  INV_X1    g353(.A(new_n522), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n540), .A2(KEYINPUT74), .A3(new_n520), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT74), .B1(new_n540), .B2(new_n520), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n535), .B(new_n278), .C1(new_n539), .C2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n514), .B1(new_n533), .B2(new_n534), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n541), .A2(new_n542), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n549), .A2(KEYINPUT25), .A3(new_n278), .A4(new_n535), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n412), .B1(G234), .B2(new_n278), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n544), .A2(new_n553), .A3(new_n545), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n549), .A2(new_n535), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n552), .A2(G902), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G221), .B1(new_n411), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT79), .B(G469), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G110), .B(G140), .ZN(new_n564));
  INV_X1    g378(.A(G227), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(G953), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n564), .B(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n437), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n424), .A2(new_n428), .ZN(new_n569));
  AOI211_X1 g383(.A(KEYINPUT4), .B(new_n230), .C1(new_n227), .C2(new_n229), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n248), .B1(new_n247), .B2(G101), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n231), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT10), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n294), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n569), .A2(new_n572), .B1(new_n200), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n194), .B1(new_n199), .B2(new_n425), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n231), .A2(new_n576), .A3(new_n254), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT77), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n577), .A2(new_n578), .A3(new_n573), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n577), .B2(new_n573), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n568), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n577), .A2(new_n573), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT77), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n232), .A2(new_n424), .A3(new_n428), .A4(new_n249), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n200), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n578), .A3(new_n573), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n437), .ZN(new_n589));
  OAI211_X1 g403(.A(KEYINPUT80), .B(new_n567), .C1(new_n582), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n577), .B1(new_n255), .B2(new_n200), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n592), .B(new_n594), .C1(new_n595), .C2(new_n437), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n595), .A2(KEYINPUT78), .A3(new_n591), .A4(new_n437), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n575), .A2(new_n568), .A3(new_n581), .ZN(new_n600));
  INV_X1    g414(.A(new_n567), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n590), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n588), .A2(new_n437), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n601), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(KEYINPUT80), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n278), .B(new_n563), .C1(new_n603), .C2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n592), .B1(new_n595), .B2(new_n437), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n593), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n600), .A2(new_n597), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n588), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n567), .B1(new_n611), .B2(new_n568), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n610), .A2(new_n567), .B1(new_n612), .B2(new_n604), .ZN(new_n613));
  OAI21_X1  g427(.A(G469), .B1(new_n613), .B2(G902), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n561), .B1(new_n607), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n422), .A2(new_n502), .A3(new_n559), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G101), .ZN(G3));
  OAI21_X1  g431(.A(G472), .B1(new_n499), .B2(G902), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n492), .A2(new_n493), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n559), .A3(new_n615), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n276), .B1(new_n273), .B2(new_n297), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n303), .A2(new_n275), .A3(new_n304), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n187), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  OAI22_X1  g440(.A1(new_n414), .A2(new_n415), .B1(KEYINPUT95), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n404), .A2(new_n410), .ZN(new_n628));
  INV_X1    g442(.A(new_n413), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n404), .A2(new_n410), .A3(new_n413), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n632));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n627), .A2(new_n633), .A3(G478), .A4(new_n278), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n416), .A2(new_n417), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n373), .B1(new_n372), .B2(new_n362), .ZN(new_n638));
  AOI211_X1 g452(.A(KEYINPUT20), .B(new_n363), .C1(new_n368), .C2(new_n371), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n367), .A2(new_n333), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n370), .ZN(new_n641));
  AOI21_X1  g455(.A(G902), .B1(new_n641), .B2(new_n368), .ZN(new_n642));
  INV_X1    g456(.A(G475), .ZN(new_n643));
  OAI22_X1  g457(.A1(new_n638), .A2(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NOR4_X1   g459(.A1(new_n622), .A2(new_n385), .A3(new_n625), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT34), .B(G104), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n377), .A2(G475), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n649), .B(new_n419), .C1(new_n638), .C2(new_n639), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT96), .B1(new_n650), .B2(new_n385), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n378), .A2(new_n652), .A3(new_n386), .A4(new_n419), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n622), .A2(new_n655), .A3(new_n625), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT35), .B(G107), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  OAI21_X1  g472(.A(new_n547), .B1(new_n548), .B2(KEYINPUT36), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT36), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n539), .A2(new_n660), .A3(new_n543), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n659), .A2(new_n557), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n555), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n555), .A2(KEYINPUT97), .A3(new_n663), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n421), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n306), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n621), .A3(new_n615), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  NAND2_X1  g488(.A1(new_n502), .A2(new_n615), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n554), .A2(new_n552), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n665), .B(new_n662), .C1(new_n677), .C2(new_n551), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT97), .B1(new_n555), .B2(new_n663), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n380), .B1(new_n383), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n650), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n680), .A2(new_n684), .A3(new_n625), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n676), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT100), .B(G128), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G30));
  XOR2_X1   g502(.A(new_n682), .B(KEYINPUT39), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n615), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT40), .Z(new_n691));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n680), .A2(new_n187), .A3(new_n419), .A4(new_n644), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT38), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n298), .B2(new_n305), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n277), .B1(new_n273), .B2(new_n297), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n303), .A2(new_n299), .A3(new_n304), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT38), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n496), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n462), .B1(new_n473), .B2(new_n444), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n278), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G472), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n494), .A2(new_n501), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n695), .A2(new_n701), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n693), .A2(new_n694), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT102), .B(G143), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G45));
  NAND2_X1  g525(.A1(new_n364), .A2(new_n374), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n636), .B1(new_n712), .B2(new_n649), .ZN(new_n713));
  INV_X1    g527(.A(new_n682), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n680), .A2(new_n625), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n676), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  INV_X1    g532(.A(new_n559), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n498), .A2(new_n490), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n500), .B1(new_n720), .B2(new_n483), .ZN(new_n721));
  AOI22_X1  g535(.A1(KEYINPUT32), .A2(new_n721), .B1(new_n480), .B2(G472), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n722), .B2(new_n501), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n645), .A2(new_n385), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n605), .A2(KEYINPUT80), .B1(new_n612), .B2(new_n599), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n567), .B1(new_n582), .B2(new_n589), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT80), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(G902), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(G469), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n607), .B(new_n560), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n625), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n723), .A2(new_n724), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  NAND3_X1  g549(.A1(new_n723), .A2(new_n654), .A3(new_n732), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  AND2_X1   g551(.A1(new_n668), .A2(new_n502), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n607), .B1(new_n729), .B2(new_n730), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  INV_X1    g555(.A(new_n625), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n740), .A2(new_n741), .A3(new_n560), .A4(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT103), .B1(new_n731), .B2(new_n625), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n738), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  INV_X1    g560(.A(new_n731), .ZN(new_n747));
  INV_X1    g561(.A(new_n462), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n474), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n486), .B2(new_n491), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n493), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n618), .A2(new_n559), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n644), .A2(new_n419), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n385), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n747), .A2(new_n752), .A3(new_n742), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  OAI211_X1 g570(.A(new_n618), .B(new_n751), .C1(new_n678), .C2(new_n679), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n715), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n743), .A2(new_n758), .A3(new_n744), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  INV_X1    g574(.A(KEYINPUT32), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n499), .B2(new_n500), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n481), .A2(new_n494), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n559), .ZN(new_n764));
  INV_X1    g578(.A(new_n715), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n698), .A2(new_n699), .A3(new_n187), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n615), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT42), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n615), .A2(new_n766), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n715), .A2(KEYINPUT42), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n723), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n341), .ZN(G33));
  NAND4_X1  g587(.A1(new_n502), .A2(new_n559), .A3(new_n615), .A4(new_n766), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT104), .B1(new_n774), .B2(new_n684), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT104), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n723), .A2(new_n769), .A3(new_n776), .A4(new_n683), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  NAND2_X1  g593(.A1(new_n612), .A2(new_n604), .ZN(new_n780));
  INV_X1    g594(.A(new_n610), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n780), .B1(new_n781), .B2(new_n601), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n730), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n613), .A2(KEYINPUT45), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n784), .A2(new_n785), .B1(G469), .B2(G902), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n607), .B1(new_n786), .B2(KEYINPUT46), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT105), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n561), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n378), .A2(new_n637), .ZN(new_n794));
  AND2_X1   g608(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n795));
  NOR2_X1   g609(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n378), .B(new_n637), .C1(KEYINPUT106), .C2(KEYINPUT43), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n799), .B(new_n620), .C1(new_n679), .C2(new_n678), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n766), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n800), .B2(new_n801), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n793), .A2(new_n689), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  NOR2_X1   g620(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  OAI22_X1  g623(.A1(new_n792), .A2(new_n561), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n791), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT105), .B1(new_n786), .B2(KEYINPUT46), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n560), .B(new_n808), .C1(new_n813), .C2(new_n787), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n502), .A2(new_n803), .A3(new_n559), .A4(new_n715), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n810), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT108), .B(G140), .Z(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(G42));
  XOR2_X1   g632(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n616), .A2(new_n670), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n743), .A2(new_n744), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n738), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n502), .A2(new_n559), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n747), .A2(new_n654), .A3(new_n742), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n740), .A2(new_n560), .A3(new_n742), .A4(new_n724), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n644), .A2(new_n420), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n386), .B1(new_n828), .B2(new_n713), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n306), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n559), .A3(new_n615), .A4(new_n621), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n755), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n772), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n823), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n676), .B1(new_n685), .B2(new_n716), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n625), .A2(new_n753), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n664), .A2(new_n682), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n706), .A3(new_n615), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n836), .A2(new_n759), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n836), .A2(new_n759), .A3(KEYINPUT52), .A4(new_n839), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n835), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n644), .A2(new_n419), .A3(new_n682), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n766), .B(new_n845), .C1(new_n679), .C2(new_n678), .ZN(new_n846));
  OAI22_X1  g660(.A1(new_n675), .A2(new_n846), .B1(new_n767), .B2(new_n757), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n778), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT110), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT110), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n778), .A2(new_n851), .A3(new_n848), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n820), .B1(new_n844), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n842), .A2(new_n843), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n745), .A2(new_n616), .A3(new_n670), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n736), .A2(new_n733), .A3(new_n755), .A4(new_n831), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n857), .A3(new_n772), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  AOI211_X1 g673(.A(KEYINPUT110), .B(new_n847), .C1(new_n777), .C2(new_n775), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n851), .B1(new_n778), .B2(new_n848), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n859), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n854), .A2(new_n864), .A3(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n380), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n803), .A2(new_n731), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(new_n799), .ZN(new_n869));
  INV_X1    g683(.A(new_n757), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n706), .A2(new_n719), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n868), .A2(new_n378), .A3(new_n872), .A4(new_n636), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT51), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n187), .B1(new_n697), .B2(new_n700), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n867), .B1(new_n797), .B2(new_n798), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n747), .A4(new_n752), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT50), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT50), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n810), .A2(new_n814), .B1(new_n561), .B2(new_n740), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n876), .A2(new_n752), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n766), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n874), .B(new_n883), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n869), .A2(new_n559), .A3(new_n763), .ZN(new_n888));
  NOR2_X1   g702(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT119), .Z(new_n890));
  AOI22_X1  g704(.A1(new_n888), .A2(new_n890), .B1(KEYINPUT120), .B2(KEYINPUT48), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n868), .A2(new_n713), .A3(new_n872), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(G952), .A3(new_n211), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n822), .A2(new_n885), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT117), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n822), .A2(new_n885), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(KEYINPUT118), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n901), .B(new_n894), .C1(new_n896), .C2(new_n898), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n887), .B(new_n892), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n871), .A2(new_n873), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n881), .A2(KEYINPUT115), .A3(new_n882), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT115), .B1(new_n881), .B2(new_n882), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT116), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT116), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n909), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n908), .B(new_n910), .C1(new_n884), .C2(new_n886), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n903), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n853), .A2(new_n855), .A3(new_n858), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT111), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n863), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n914), .B2(new_n863), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n914), .A2(new_n819), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n866), .B(new_n913), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(G952), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n211), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n739), .B(KEYINPUT49), .Z(new_n925));
  INV_X1    g739(.A(new_n187), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n794), .A2(new_n561), .A3(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n925), .A2(new_n701), .A3(new_n872), .A4(new_n927), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT109), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n924), .A2(new_n929), .ZN(G75));
  NAND2_X1  g744(.A1(new_n922), .A2(G953), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT123), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n914), .A2(new_n819), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n844), .A2(KEYINPUT53), .A3(new_n853), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n278), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(new_n275), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n270), .A2(new_n215), .A3(new_n272), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(new_n303), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n932), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(G902), .B1(new_n854), .B2(new_n864), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT121), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n943), .B(G902), .C1(new_n854), .C2(new_n864), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n275), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n939), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n939), .A2(new_n946), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT56), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n940), .B1(new_n945), .B2(new_n949), .ZN(G51));
  INV_X1    g764(.A(new_n932), .ZN(new_n951));
  NAND2_X1  g765(.A1(G469), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT57), .Z(new_n953));
  AOI21_X1  g767(.A(new_n920), .B1(new_n933), .B2(new_n934), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n865), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n725), .A2(new_n728), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT124), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n942), .A2(new_n785), .A3(new_n784), .A4(new_n944), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(G54));
  AND2_X1   g774(.A1(KEYINPUT58), .A2(G475), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n942), .A2(new_n944), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n372), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n942), .A2(new_n361), .A3(new_n944), .A4(new_n961), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n951), .B1(new_n963), .B2(new_n964), .ZN(G60));
  NAND2_X1  g779(.A1(new_n627), .A2(new_n633), .ZN(new_n966));
  NAND2_X1  g780(.A1(G478), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT59), .Z(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n865), .B2(new_n954), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n932), .ZN(new_n971));
  INV_X1    g785(.A(new_n968), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n917), .A2(new_n918), .ZN(new_n973));
  INV_X1    g787(.A(new_n916), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n920), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n972), .B1(new_n975), .B2(new_n865), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n971), .B1(new_n976), .B2(new_n966), .ZN(G63));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  NAND2_X1  g792(.A1(G217), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT60), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n933), .B2(new_n934), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n659), .A2(new_n661), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n556), .B(KEYINPUT125), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n932), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n978), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n981), .A2(new_n985), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n932), .A4(new_n983), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(G66));
  OAI21_X1  g804(.A(G953), .B1(new_n384), .B2(new_n209), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n856), .A2(new_n857), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(G953), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n270), .B(new_n272), .C1(G898), .C2(new_n211), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT126), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n993), .B(new_n995), .ZN(G69));
  AND2_X1   g810(.A1(new_n836), .A2(new_n759), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n834), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n793), .A2(new_n689), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n764), .A2(new_n625), .A3(new_n753), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(new_n778), .A3(new_n805), .A4(new_n816), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1002), .A2(G953), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n466), .A2(new_n467), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT127), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(new_n340), .Z(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n681), .B2(new_n211), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n709), .A2(new_n997), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n803), .B1(new_n645), .B2(new_n650), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1011), .A2(new_n723), .A3(new_n615), .A4(new_n689), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n816), .A2(new_n805), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n709), .A2(new_n1014), .A3(new_n997), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1010), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1006), .B1(new_n1016), .B2(new_n211), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1008), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(G953), .B1(new_n565), .B2(new_n681), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(G72));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  INV_X1    g836(.A(new_n992), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1022), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n470), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n1025), .A2(new_n461), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1022), .B1(new_n1002), .B2(new_n1023), .ZN(new_n1028));
  OR2_X1    g842(.A1(new_n1025), .A2(new_n461), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n951), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n919), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1022), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1030), .A2(new_n1026), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1032), .B1(new_n1033), .B2(new_n1035), .ZN(G57));
endmodule


