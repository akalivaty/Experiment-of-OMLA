

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768;

  AND2_X1 U368 ( .A1(n645), .A2(n644), .ZN(n647) );
  XNOR2_X1 U369 ( .A(n756), .B(n348), .ZN(n347) );
  INV_X1 U370 ( .A(KEYINPUT73), .ZN(n348) );
  OR2_X1 U371 ( .A1(n583), .A2(n594), .ZN(n584) );
  NOR2_X1 U372 ( .A1(n566), .A2(n537), .ZN(n678) );
  XNOR2_X1 U373 ( .A(n507), .B(n428), .ZN(n753) );
  INV_X1 U374 ( .A(KEYINPUT3), .ZN(n387) );
  XNOR2_X2 U375 ( .A(n380), .B(n587), .ZN(n375) );
  AND2_X2 U376 ( .A1(n376), .A2(n657), .ZN(n403) );
  XNOR2_X2 U377 ( .A(n481), .B(KEYINPUT4), .ZN(n507) );
  NAND2_X1 U378 ( .A1(n368), .A2(n347), .ZN(n371) );
  OR2_X2 U379 ( .A1(n630), .A2(G902), .ZN(n438) );
  NOR2_X1 U380 ( .A1(G953), .A2(G237), .ZN(n490) );
  INV_X1 U381 ( .A(G953), .ZN(n463) );
  NOR2_X1 U382 ( .A1(n627), .A2(KEYINPUT67), .ZN(n376) );
  XNOR2_X1 U383 ( .A(n378), .B(n377), .ZN(n627) );
  AND2_X1 U384 ( .A1(n367), .A2(n365), .ZN(n361) );
  XOR2_X1 U385 ( .A(KEYINPUT109), .B(n534), .Z(n765) );
  XNOR2_X1 U386 ( .A(n611), .B(n610), .ZN(n619) );
  XNOR2_X1 U387 ( .A(KEYINPUT103), .B(n538), .ZN(n714) );
  XNOR2_X1 U388 ( .A(n384), .B(n532), .ZN(n536) );
  AND2_X1 U389 ( .A1(n400), .A2(n351), .ZN(n399) );
  NAND2_X1 U390 ( .A1(n373), .A2(KEYINPUT2), .ZN(n370) );
  NAND2_X1 U391 ( .A1(n648), .A2(n639), .ZN(n378) );
  INV_X1 U392 ( .A(KEYINPUT69), .ZN(n426) );
  INV_X1 U393 ( .A(G237), .ZN(n516) );
  XNOR2_X1 U394 ( .A(n396), .B(n411), .ZN(n395) );
  INV_X1 U395 ( .A(KEYINPUT46), .ZN(n411) );
  OR2_X1 U396 ( .A1(n767), .A2(n766), .ZN(n396) );
  XNOR2_X1 U397 ( .A(n385), .B(n435), .ZN(n505) );
  XNOR2_X1 U398 ( .A(G113), .B(G116), .ZN(n435) );
  XNOR2_X1 U399 ( .A(n387), .B(G119), .ZN(n385) );
  NAND2_X1 U400 ( .A1(n353), .A2(n539), .ZN(n392) );
  NAND2_X1 U401 ( .A1(n383), .A2(n544), .ZN(n621) );
  XNOR2_X1 U402 ( .A(n536), .B(n382), .ZN(n383) );
  INV_X1 U403 ( .A(KEYINPUT1), .ZN(n382) );
  INV_X1 U404 ( .A(n369), .ZN(n364) );
  NOR2_X1 U405 ( .A1(n379), .A2(n413), .ZN(n416) );
  XNOR2_X1 U406 ( .A(G478), .B(KEYINPUT102), .ZN(n484) );
  XNOR2_X1 U407 ( .A(n584), .B(n595), .ZN(n586) );
  INV_X1 U408 ( .A(n383), .ZN(n699) );
  XNOR2_X1 U409 ( .A(G902), .B(KEYINPUT87), .ZN(n453) );
  XOR2_X1 U410 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n430) );
  XNOR2_X1 U411 ( .A(n398), .B(n557), .ZN(n397) );
  NAND2_X1 U412 ( .A1(n556), .A2(n765), .ZN(n398) );
  AND2_X1 U413 ( .A1(n555), .A2(n423), .ZN(n556) );
  XNOR2_X1 U414 ( .A(G113), .B(G143), .ZN(n493) );
  XNOR2_X1 U415 ( .A(G134), .B(G137), .ZN(n427) );
  NOR2_X1 U416 ( .A1(n628), .A2(n629), .ZN(n368) );
  INV_X1 U417 ( .A(n629), .ZN(n373) );
  XNOR2_X1 U418 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n508) );
  NAND2_X1 U419 ( .A1(n366), .A2(KEYINPUT74), .ZN(n365) );
  INV_X1 U420 ( .A(KEYINPUT74), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n381), .B(KEYINPUT33), .ZN(n689) );
  NAND2_X1 U422 ( .A1(n414), .A2(n413), .ZN(n381) );
  XNOR2_X1 U423 ( .A(n621), .B(KEYINPUT105), .ZN(n414) );
  AND2_X1 U424 ( .A1(n535), .A2(n409), .ZN(n408) );
  INV_X1 U425 ( .A(G902), .ZN(n531) );
  OR2_X1 U426 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U427 ( .A(n529), .B(n386), .ZN(n748) );
  XNOR2_X1 U428 ( .A(n505), .B(n504), .ZN(n386) );
  XOR2_X1 U429 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n422) );
  XNOR2_X1 U430 ( .A(G119), .B(G110), .ZN(n448) );
  XNOR2_X1 U431 ( .A(G116), .B(G107), .ZN(n479) );
  XNOR2_X1 U432 ( .A(n753), .B(G146), .ZN(n393) );
  XNOR2_X1 U433 ( .A(n389), .B(n388), .ZN(n529) );
  XNOR2_X1 U434 ( .A(G101), .B(G107), .ZN(n388) );
  XNOR2_X1 U435 ( .A(n506), .B(KEYINPUT72), .ZN(n389) );
  XNOR2_X1 U436 ( .A(G110), .B(G104), .ZN(n506) );
  INV_X1 U437 ( .A(KEYINPUT34), .ZN(n587) );
  XNOR2_X1 U438 ( .A(KEYINPUT30), .B(KEYINPUT108), .ZN(n541) );
  NAND2_X1 U439 ( .A1(n659), .A2(G475), .ZN(n643) );
  BUF_X1 U440 ( .A(n659), .Z(n735) );
  AND2_X1 U441 ( .A1(n635), .A2(G953), .ZN(n739) );
  XNOR2_X1 U442 ( .A(n564), .B(KEYINPUT40), .ZN(n767) );
  INV_X1 U443 ( .A(n614), .ZN(n421) );
  AND2_X1 U444 ( .A1(n586), .A2(n390), .ZN(n623) );
  INV_X1 U445 ( .A(n703), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(KEYINPUT104), .ZN(n768) );
  NAND2_X1 U447 ( .A1(n349), .A2(n354), .ZN(n391) );
  AND2_X1 U448 ( .A1(n619), .A2(n612), .ZN(n349) );
  AND2_X1 U449 ( .A1(n620), .A2(KEYINPUT67), .ZN(n350) );
  AND2_X1 U450 ( .A1(n392), .A2(n768), .ZN(n351) );
  OR2_X1 U451 ( .A1(n679), .A2(n665), .ZN(n353) );
  AND2_X1 U452 ( .A1(n699), .A2(n626), .ZN(n354) );
  AND2_X1 U453 ( .A1(n740), .A2(n363), .ZN(n355) );
  AND2_X1 U454 ( .A1(n740), .A2(n756), .ZN(n356) );
  AND2_X1 U455 ( .A1(n615), .A2(n409), .ZN(n357) );
  AND2_X1 U456 ( .A1(n625), .A2(n615), .ZN(n358) );
  XOR2_X1 U457 ( .A(KEYINPUT81), .B(KEYINPUT45), .Z(n359) );
  XOR2_X1 U458 ( .A(n642), .B(n641), .Z(n360) );
  NOR2_X4 U459 ( .A1(n579), .A2(n578), .ZN(n756) );
  NAND2_X1 U460 ( .A1(n361), .A2(n362), .ZN(n688) );
  NOR2_X1 U461 ( .A1(n408), .A2(n357), .ZN(n407) );
  NAND2_X1 U462 ( .A1(n364), .A2(n355), .ZN(n362) );
  INV_X1 U463 ( .A(n740), .ZN(n366) );
  NAND2_X1 U464 ( .A1(n369), .A2(KEYINPUT74), .ZN(n367) );
  NAND2_X1 U465 ( .A1(n756), .A2(KEYINPUT2), .ZN(n369) );
  NAND2_X1 U466 ( .A1(n371), .A2(n370), .ZN(n372) );
  AND2_X2 U467 ( .A1(n372), .A2(n688), .ZN(n659) );
  XNOR2_X2 U468 ( .A(n374), .B(n589), .ZN(n657) );
  NAND2_X2 U469 ( .A1(n375), .A2(n588), .ZN(n374) );
  INV_X1 U470 ( .A(KEYINPUT83), .ZN(n377) );
  NAND2_X1 U471 ( .A1(n617), .A2(n613), .ZN(n379) );
  NOR2_X1 U472 ( .A1(n379), .A2(n419), .ZN(n418) );
  NAND2_X1 U473 ( .A1(n689), .A2(n586), .ZN(n380) );
  NAND2_X1 U474 ( .A1(n729), .A2(n531), .ZN(n384) );
  AND2_X1 U475 ( .A1(n586), .A2(n358), .ZN(n665) );
  XNOR2_X1 U476 ( .A(n393), .B(n437), .ZN(n630) );
  XNOR2_X1 U477 ( .A(n393), .B(n530), .ZN(n729) );
  XNOR2_X2 U478 ( .A(n394), .B(KEYINPUT48), .ZN(n579) );
  NAND2_X1 U479 ( .A1(n397), .A2(n395), .ZN(n394) );
  NAND2_X1 U480 ( .A1(n402), .A2(n399), .ZN(n412) );
  NAND2_X1 U481 ( .A1(n401), .A2(n350), .ZN(n400) );
  INV_X1 U482 ( .A(n657), .ZN(n401) );
  XNOR2_X1 U483 ( .A(n403), .B(KEYINPUT44), .ZN(n402) );
  NAND2_X1 U484 ( .A1(n407), .A2(n404), .ZN(n410) );
  NAND2_X1 U485 ( .A1(n406), .A2(n405), .ZN(n404) );
  NOR2_X1 U486 ( .A1(n615), .A2(n409), .ZN(n405) );
  INV_X1 U487 ( .A(n535), .ZN(n406) );
  INV_X1 U488 ( .A(KEYINPUT28), .ZN(n409) );
  NOR2_X2 U489 ( .A1(n568), .A2(n583), .ZN(n673) );
  NAND2_X1 U490 ( .A1(n410), .A2(n548), .ZN(n568) );
  XNOR2_X2 U491 ( .A(n412), .B(n359), .ZN(n740) );
  INV_X1 U492 ( .A(n612), .ZN(n413) );
  NAND2_X1 U493 ( .A1(n415), .A2(n421), .ZN(n420) );
  NAND2_X1 U494 ( .A1(n619), .A2(n416), .ZN(n415) );
  NAND2_X1 U495 ( .A1(n420), .A2(n417), .ZN(n648) );
  NAND2_X1 U496 ( .A1(n619), .A2(n418), .ZN(n417) );
  NAND2_X1 U497 ( .A1(n612), .A2(n614), .ZN(n419) );
  NAND2_X1 U498 ( .A1(n523), .A2(n708), .ZN(n524) );
  BUF_X1 U499 ( .A(n546), .Z(n576) );
  OR2_X1 U500 ( .A1(KEYINPUT47), .A2(n554), .ZN(n423) );
  XOR2_X1 U501 ( .A(n478), .B(n477), .Z(n424) );
  NAND2_X1 U502 ( .A1(n673), .A2(n539), .ZN(n554) );
  INV_X1 U503 ( .A(KEYINPUT70), .ZN(n557) );
  XNOR2_X1 U504 ( .A(n473), .B(n472), .ZN(n502) );
  BUF_X1 U505 ( .A(n753), .Z(n755) );
  XNOR2_X1 U506 ( .A(n485), .B(n484), .ZN(n566) );
  XNOR2_X1 U507 ( .A(n542), .B(n541), .ZN(n561) );
  XNOR2_X1 U508 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X2 U509 ( .A(G143), .B(KEYINPUT64), .ZN(n425) );
  XNOR2_X2 U510 ( .A(n425), .B(G128), .ZN(n481) );
  XNOR2_X1 U511 ( .A(n426), .B(G131), .ZN(n486) );
  XNOR2_X1 U512 ( .A(n486), .B(n427), .ZN(n428) );
  NAND2_X1 U513 ( .A1(n490), .A2(G210), .ZN(n429) );
  XNOR2_X1 U514 ( .A(n430), .B(n429), .ZN(n432) );
  INV_X1 U515 ( .A(KEYINPUT96), .ZN(n431) );
  XNOR2_X1 U516 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U517 ( .A(G101), .B(KEYINPUT94), .ZN(n433) );
  XNOR2_X1 U518 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U519 ( .A(n505), .B(n436), .ZN(n437) );
  XNOR2_X2 U520 ( .A(n438), .B(G472), .ZN(n540) );
  XNOR2_X1 U521 ( .A(n540), .B(KEYINPUT6), .ZN(n585) );
  NAND2_X1 U522 ( .A1(G234), .A2(n463), .ZN(n439) );
  XNOR2_X1 U523 ( .A(n422), .B(n439), .ZN(n476) );
  NAND2_X1 U524 ( .A1(n476), .A2(G221), .ZN(n444) );
  XNOR2_X1 U525 ( .A(G128), .B(G137), .ZN(n440) );
  XNOR2_X1 U526 ( .A(n440), .B(KEYINPUT80), .ZN(n442) );
  XNOR2_X1 U527 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n441) );
  XNOR2_X1 U528 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U529 ( .A(n444), .B(n443), .ZN(n451) );
  XNOR2_X1 U530 ( .A(G146), .B(G125), .ZN(n509) );
  INV_X1 U531 ( .A(KEYINPUT10), .ZN(n445) );
  XNOR2_X1 U532 ( .A(n445), .B(G140), .ZN(n446) );
  XNOR2_X1 U533 ( .A(n509), .B(n446), .ZN(n488) );
  INV_X1 U534 ( .A(n488), .ZN(n754) );
  XNOR2_X1 U535 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n447) );
  XNOR2_X1 U536 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U537 ( .A(n754), .B(n449), .ZN(n450) );
  XNOR2_X1 U538 ( .A(n451), .B(n450), .ZN(n660) );
  NAND2_X1 U539 ( .A1(n660), .A2(n531), .ZN(n457) );
  INV_X1 U540 ( .A(KEYINPUT15), .ZN(n452) );
  XNOR2_X1 U541 ( .A(n453), .B(n452), .ZN(n629) );
  NAND2_X1 U542 ( .A1(n629), .A2(G234), .ZN(n454) );
  XNOR2_X1 U543 ( .A(n454), .B(KEYINPUT20), .ZN(n458) );
  NAND2_X1 U544 ( .A1(n458), .A2(G217), .ZN(n455) );
  XNOR2_X1 U545 ( .A(n455), .B(KEYINPUT25), .ZN(n456) );
  XNOR2_X2 U546 ( .A(n457), .B(n456), .ZN(n613) );
  INV_X1 U547 ( .A(n613), .ZN(n626) );
  INV_X1 U548 ( .A(n458), .ZN(n460) );
  INV_X1 U549 ( .A(G221), .ZN(n459) );
  XNOR2_X1 U550 ( .A(n461), .B(KEYINPUT21), .ZN(n694) );
  INV_X1 U551 ( .A(n694), .ZN(n469) );
  NAND2_X1 U552 ( .A1(G234), .A2(G237), .ZN(n462) );
  XNOR2_X1 U553 ( .A(n462), .B(KEYINPUT14), .ZN(n693) );
  INV_X1 U554 ( .A(G952), .ZN(n635) );
  NAND2_X1 U555 ( .A1(n463), .A2(n635), .ZN(n465) );
  OR2_X1 U556 ( .A1(n463), .A2(G902), .ZN(n464) );
  AND2_X1 U557 ( .A1(n465), .A2(n464), .ZN(n466) );
  AND2_X1 U558 ( .A1(n693), .A2(n466), .ZN(n582) );
  NAND2_X1 U559 ( .A1(G953), .A2(G900), .ZN(n467) );
  NAND2_X1 U560 ( .A1(n582), .A2(n467), .ZN(n468) );
  XOR2_X1 U561 ( .A(KEYINPUT76), .B(n468), .Z(n543) );
  NAND2_X1 U562 ( .A1(n469), .A2(n543), .ZN(n470) );
  NOR2_X1 U563 ( .A1(n626), .A2(n470), .ZN(n471) );
  XNOR2_X1 U564 ( .A(n471), .B(KEYINPUT71), .ZN(n535) );
  NOR2_X1 U565 ( .A1(n585), .A2(n535), .ZN(n473) );
  INV_X1 U566 ( .A(KEYINPUT106), .ZN(n472) );
  XOR2_X1 U567 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n475) );
  XNOR2_X1 U568 ( .A(G134), .B(KEYINPUT7), .ZN(n474) );
  XNOR2_X1 U569 ( .A(n475), .B(n474), .ZN(n478) );
  NAND2_X1 U570 ( .A1(G217), .A2(n476), .ZN(n477) );
  XOR2_X1 U571 ( .A(KEYINPUT100), .B(G122), .Z(n480) );
  XNOR2_X1 U572 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U573 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U574 ( .A(n424), .B(n483), .ZN(n736) );
  NOR2_X1 U575 ( .A1(n736), .A2(G902), .ZN(n485) );
  XNOR2_X1 U576 ( .A(n486), .B(G104), .ZN(n487) );
  XNOR2_X1 U577 ( .A(n487), .B(G122), .ZN(n489) );
  XNOR2_X1 U578 ( .A(n489), .B(n488), .ZN(n498) );
  XOR2_X1 U579 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n492) );
  NAND2_X1 U580 ( .A1(G214), .A2(n490), .ZN(n491) );
  XNOR2_X1 U581 ( .A(n492), .B(n491), .ZN(n496) );
  XOR2_X1 U582 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n494) );
  XNOR2_X1 U583 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U584 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U585 ( .A(n498), .B(n497), .ZN(n642) );
  NAND2_X1 U586 ( .A1(n642), .A2(n531), .ZN(n500) );
  XNOR2_X1 U587 ( .A(KEYINPUT13), .B(G475), .ZN(n499) );
  XNOR2_X1 U588 ( .A(n500), .B(n499), .ZN(n565) );
  INV_X1 U589 ( .A(n565), .ZN(n537) );
  AND2_X1 U590 ( .A1(n566), .A2(n537), .ZN(n676) );
  INV_X1 U591 ( .A(n676), .ZN(n501) );
  NOR2_X2 U592 ( .A1(n502), .A2(n501), .ZN(n571) );
  INV_X1 U593 ( .A(KEYINPUT16), .ZN(n503) );
  XNOR2_X1 U594 ( .A(n503), .B(G122), .ZN(n504) );
  INV_X1 U595 ( .A(n507), .ZN(n514) );
  XNOR2_X1 U596 ( .A(n509), .B(n508), .ZN(n512) );
  NAND2_X1 U597 ( .A1(n463), .A2(G224), .ZN(n510) );
  XNOR2_X1 U598 ( .A(n510), .B(KEYINPUT88), .ZN(n511) );
  XNOR2_X1 U599 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U600 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U601 ( .A(n748), .B(n515), .ZN(n650) );
  NAND2_X1 U602 ( .A1(n650), .A2(n629), .ZN(n521) );
  NAND2_X1 U603 ( .A1(n531), .A2(n516), .ZN(n522) );
  NAND2_X1 U604 ( .A1(n522), .A2(G210), .ZN(n519) );
  INV_X1 U605 ( .A(KEYINPUT89), .ZN(n517) );
  XNOR2_X1 U606 ( .A(n517), .B(KEYINPUT90), .ZN(n518) );
  XNOR2_X1 U607 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U608 ( .A(n521), .B(n520), .ZN(n546) );
  INV_X1 U609 ( .A(n546), .ZN(n523) );
  NAND2_X1 U610 ( .A1(n522), .A2(G214), .ZN(n708) );
  XNOR2_X2 U611 ( .A(n524), .B(KEYINPUT85), .ZN(n607) );
  NAND2_X1 U612 ( .A1(n571), .A2(n607), .ZN(n526) );
  XOR2_X1 U613 ( .A(KEYINPUT36), .B(KEYINPUT84), .Z(n525) );
  XNOR2_X1 U614 ( .A(n526), .B(n525), .ZN(n533) );
  NAND2_X1 U615 ( .A1(n463), .A2(G227), .ZN(n527) );
  XNOR2_X1 U616 ( .A(n527), .B(G140), .ZN(n528) );
  XNOR2_X1 U617 ( .A(n529), .B(n528), .ZN(n530) );
  INV_X1 U618 ( .A(G469), .ZN(n532) );
  INV_X1 U619 ( .A(n699), .ZN(n617) );
  NAND2_X1 U620 ( .A1(n533), .A2(n617), .ZN(n534) );
  INV_X1 U621 ( .A(n540), .ZN(n615) );
  BUF_X1 U622 ( .A(n536), .Z(n624) );
  INV_X1 U623 ( .A(n624), .ZN(n548) );
  XNOR2_X1 U624 ( .A(n607), .B(KEYINPUT19), .ZN(n583) );
  OR2_X1 U625 ( .A1(n678), .A2(n676), .ZN(n538) );
  INV_X1 U626 ( .A(n714), .ZN(n539) );
  NAND2_X1 U627 ( .A1(n554), .A2(KEYINPUT47), .ZN(n552) );
  NAND2_X1 U628 ( .A1(n708), .A2(n540), .ZN(n542) );
  NOR2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n588) );
  OR2_X1 U630 ( .A1(n613), .A2(n694), .ZN(n698) );
  INV_X1 U631 ( .A(n698), .ZN(n544) );
  NAND2_X1 U632 ( .A1(n544), .A2(n543), .ZN(n558) );
  INV_X1 U633 ( .A(n558), .ZN(n545) );
  NAND2_X1 U634 ( .A1(n588), .A2(n545), .ZN(n547) );
  NOR2_X1 U635 ( .A1(n547), .A2(n576), .ZN(n549) );
  NAND2_X1 U636 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U637 ( .A1(n561), .A2(n550), .ZN(n640) );
  INV_X1 U638 ( .A(n640), .ZN(n551) );
  NAND2_X1 U639 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U640 ( .A(n553), .B(KEYINPUT79), .ZN(n555) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT38), .ZN(n709) );
  NOR2_X1 U642 ( .A1(n624), .A2(n558), .ZN(n559) );
  NAND2_X1 U643 ( .A1(n709), .A2(n559), .ZN(n560) );
  NOR2_X1 U644 ( .A1(n561), .A2(n560), .ZN(n563) );
  INV_X1 U645 ( .A(KEYINPUT39), .ZN(n562) );
  XNOR2_X1 U646 ( .A(n563), .B(n562), .ZN(n570) );
  AND2_X1 U647 ( .A1(n676), .A2(n570), .ZN(n564) );
  NAND2_X1 U648 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U649 ( .A1(n566), .A2(n565), .ZN(n711) );
  NOR2_X1 U650 ( .A1(n713), .A2(n711), .ZN(n567) );
  XNOR2_X1 U651 ( .A(n567), .B(KEYINPUT41), .ZN(n706) );
  NOR2_X1 U652 ( .A1(n706), .A2(n568), .ZN(n569) );
  XNOR2_X1 U653 ( .A(n569), .B(KEYINPUT42), .ZN(n766) );
  NAND2_X1 U654 ( .A1(n570), .A2(n678), .ZN(n682) );
  BUF_X1 U655 ( .A(n571), .Z(n572) );
  NAND2_X1 U656 ( .A1(n572), .A2(n708), .ZN(n573) );
  OR2_X1 U657 ( .A1(n573), .A2(n617), .ZN(n575) );
  XOR2_X1 U658 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n574) );
  XNOR2_X1 U659 ( .A(n575), .B(n574), .ZN(n577) );
  NAND2_X1 U660 ( .A1(n577), .A2(n576), .ZN(n683) );
  NAND2_X1 U661 ( .A1(n682), .A2(n683), .ZN(n578) );
  XNOR2_X1 U662 ( .A(KEYINPUT86), .B(KEYINPUT0), .ZN(n603) );
  INV_X1 U663 ( .A(KEYINPUT91), .ZN(n580) );
  XNOR2_X1 U664 ( .A(n580), .B(G898), .ZN(n746) );
  NAND2_X1 U665 ( .A1(n746), .A2(G953), .ZN(n581) );
  NAND2_X1 U666 ( .A1(n582), .A2(n581), .ZN(n594) );
  BUF_X1 U667 ( .A(n585), .Z(n612) );
  INV_X1 U668 ( .A(KEYINPUT35), .ZN(n589) );
  INV_X1 U669 ( .A(n603), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n595), .A2(KEYINPUT19), .ZN(n590) );
  NOR2_X1 U671 ( .A1(n594), .A2(n590), .ZN(n592) );
  NOR2_X1 U672 ( .A1(n595), .A2(KEYINPUT19), .ZN(n591) );
  NOR2_X1 U673 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U674 ( .A1(n607), .A2(n593), .ZN(n600) );
  INV_X1 U675 ( .A(n711), .ZN(n598) );
  INV_X1 U676 ( .A(n594), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n602), .A2(n595), .ZN(n596) );
  NOR2_X1 U678 ( .A1(n694), .A2(n596), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U680 ( .A1(n600), .A2(n599), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n603), .A2(KEYINPUT19), .ZN(n601) );
  NAND2_X1 U682 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U683 ( .A1(n603), .A2(KEYINPUT19), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n611) );
  XNOR2_X1 U687 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n610) );
  XNOR2_X1 U688 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n615), .A2(n613), .ZN(n616) );
  NOR2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n639) );
  INV_X1 U692 ( .A(n627), .ZN(n620) );
  OR2_X1 U693 ( .A1(n621), .A2(n615), .ZN(n703) );
  XNOR2_X1 U694 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n623), .B(n622), .ZN(n679) );
  NOR2_X1 U696 ( .A1(n624), .A2(n698), .ZN(n625) );
  INV_X1 U697 ( .A(n740), .ZN(n628) );
  NAND2_X1 U698 ( .A1(n659), .A2(G472), .ZN(n634) );
  BUF_X1 U699 ( .A(n630), .Z(n632) );
  XNOR2_X1 U700 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(n636) );
  NOR2_X2 U703 ( .A1(n636), .A2(n739), .ZN(n638) );
  INV_X1 U704 ( .A(KEYINPUT63), .ZN(n637) );
  XNOR2_X1 U705 ( .A(n638), .B(n637), .ZN(G57) );
  XNOR2_X1 U706 ( .A(n639), .B(G110), .ZN(G12) );
  XOR2_X1 U707 ( .A(G143), .B(n640), .Z(G45) );
  XNOR2_X1 U708 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n641) );
  XNOR2_X1 U709 ( .A(n643), .B(n360), .ZN(n645) );
  INV_X1 U710 ( .A(n739), .ZN(n644) );
  XNOR2_X1 U711 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n647), .B(n646), .ZN(G60) );
  XNOR2_X1 U713 ( .A(n648), .B(G119), .ZN(G21) );
  NAND2_X1 U714 ( .A1(n659), .A2(G210), .ZN(n652) );
  XNOR2_X1 U715 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X2 U718 ( .A1(n653), .A2(n739), .ZN(n656) );
  XNOR2_X1 U719 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n654) );
  XNOR2_X1 U720 ( .A(n654), .B(KEYINPUT82), .ZN(n655) );
  XNOR2_X1 U721 ( .A(n656), .B(n655), .ZN(G51) );
  XOR2_X1 U722 ( .A(G122), .B(KEYINPUT127), .Z(n658) );
  XNOR2_X1 U723 ( .A(n657), .B(n658), .ZN(G24) );
  NAND2_X1 U724 ( .A1(n735), .A2(G217), .ZN(n662) );
  INV_X1 U725 ( .A(n660), .ZN(n661) );
  NOR2_X1 U726 ( .A1(n663), .A2(n739), .ZN(G66) );
  NAND2_X1 U727 ( .A1(n665), .A2(n676), .ZN(n664) );
  XNOR2_X1 U728 ( .A(n664), .B(G104), .ZN(G6) );
  XOR2_X1 U729 ( .A(KEYINPUT111), .B(KEYINPUT26), .Z(n667) );
  NAND2_X1 U730 ( .A1(n665), .A2(n678), .ZN(n666) );
  XNOR2_X1 U731 ( .A(n667), .B(n666), .ZN(n669) );
  XOR2_X1 U732 ( .A(G107), .B(KEYINPUT27), .Z(n668) );
  XNOR2_X1 U733 ( .A(n669), .B(n668), .ZN(G9) );
  XOR2_X1 U734 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n671) );
  NAND2_X1 U735 ( .A1(n673), .A2(n678), .ZN(n670) );
  XNOR2_X1 U736 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U737 ( .A(G128), .B(n672), .ZN(G30) );
  XOR2_X1 U738 ( .A(G146), .B(KEYINPUT113), .Z(n675) );
  NAND2_X1 U739 ( .A1(n673), .A2(n676), .ZN(n674) );
  XNOR2_X1 U740 ( .A(n675), .B(n674), .ZN(G48) );
  NAND2_X1 U741 ( .A1(n679), .A2(n676), .ZN(n677) );
  XNOR2_X1 U742 ( .A(n677), .B(G113), .ZN(G15) );
  NAND2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U744 ( .A(n680), .B(KEYINPUT114), .ZN(n681) );
  XNOR2_X1 U745 ( .A(G116), .B(n681), .ZN(G18) );
  XNOR2_X1 U746 ( .A(G134), .B(n682), .ZN(G36) );
  XOR2_X1 U747 ( .A(n683), .B(G140), .Z(n684) );
  XNOR2_X1 U748 ( .A(n684), .B(KEYINPUT115), .ZN(G42) );
  XNOR2_X1 U749 ( .A(KEYINPUT78), .B(KEYINPUT2), .ZN(n685) );
  NOR2_X1 U750 ( .A1(n356), .A2(n685), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n686), .B(KEYINPUT77), .ZN(n687) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n692) );
  INV_X1 U753 ( .A(n689), .ZN(n717) );
  NOR2_X1 U754 ( .A1(n706), .A2(n717), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n690), .A2(G953), .ZN(n691) );
  NAND2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n727) );
  NAND2_X1 U757 ( .A1(G952), .A2(n693), .ZN(n724) );
  NAND2_X1 U758 ( .A1(n613), .A2(n694), .ZN(n695) );
  XNOR2_X1 U759 ( .A(n695), .B(KEYINPUT49), .ZN(n696) );
  NOR2_X1 U760 ( .A1(n540), .A2(n696), .ZN(n697) );
  XNOR2_X1 U761 ( .A(KEYINPUT116), .B(n697), .ZN(n702) );
  NAND2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U763 ( .A(n700), .B(KEYINPUT50), .ZN(n701) );
  NAND2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U765 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U766 ( .A(KEYINPUT51), .B(n705), .ZN(n707) );
  NOR2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n720) );
  NOR2_X1 U768 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U770 ( .A(KEYINPUT117), .B(n712), .Z(n716) );
  NOR2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U772 ( .A1(n716), .A2(n715), .ZN(n718) );
  NOR2_X1 U773 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U774 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U775 ( .A(KEYINPUT52), .B(n721), .ZN(n722) );
  XNOR2_X1 U776 ( .A(KEYINPUT118), .B(n722), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U778 ( .A(KEYINPUT119), .B(n725), .Z(n726) );
  NOR2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U780 ( .A(KEYINPUT53), .B(n728), .ZN(G75) );
  NAND2_X1 U781 ( .A1(n735), .A2(G469), .ZN(n733) );
  XOR2_X1 U782 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n730) );
  XNOR2_X1 U783 ( .A(n730), .B(KEYINPUT121), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n729), .B(n731), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U786 ( .A1(n739), .A2(n734), .ZN(G54) );
  NAND2_X1 U787 ( .A1(n735), .A2(G478), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U789 ( .A1(n739), .A2(n738), .ZN(G63) );
  NAND2_X1 U790 ( .A1(n740), .A2(n463), .ZN(n745) );
  XOR2_X1 U791 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n742) );
  NAND2_X1 U792 ( .A1(G224), .A2(G953), .ZN(n741) );
  XNOR2_X1 U793 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U794 ( .A1(n743), .A2(n746), .ZN(n744) );
  NAND2_X1 U795 ( .A1(n745), .A2(n744), .ZN(n752) );
  NOR2_X1 U796 ( .A1(n746), .A2(n463), .ZN(n747) );
  NOR2_X1 U797 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U798 ( .A(n749), .B(KEYINPUT124), .Z(n750) );
  XNOR2_X1 U799 ( .A(KEYINPUT125), .B(n750), .ZN(n751) );
  XNOR2_X1 U800 ( .A(n752), .B(n751), .ZN(G69) );
  XNOR2_X1 U801 ( .A(n755), .B(n754), .ZN(n758) );
  XNOR2_X1 U802 ( .A(n756), .B(n758), .ZN(n757) );
  NAND2_X1 U803 ( .A1(n757), .A2(n463), .ZN(n763) );
  XOR2_X1 U804 ( .A(G227), .B(n758), .Z(n759) );
  XNOR2_X1 U805 ( .A(n759), .B(KEYINPUT126), .ZN(n760) );
  NAND2_X1 U806 ( .A1(n760), .A2(G900), .ZN(n761) );
  NAND2_X1 U807 ( .A1(n761), .A2(G953), .ZN(n762) );
  NAND2_X1 U808 ( .A1(n763), .A2(n762), .ZN(G72) );
  XOR2_X1 U809 ( .A(G125), .B(KEYINPUT37), .Z(n764) );
  XNOR2_X1 U810 ( .A(n765), .B(n764), .ZN(G27) );
  XOR2_X1 U811 ( .A(G137), .B(n766), .Z(G39) );
  XOR2_X1 U812 ( .A(G131), .B(n767), .Z(G33) );
  XNOR2_X1 U813 ( .A(G101), .B(n768), .ZN(G3) );
endmodule

