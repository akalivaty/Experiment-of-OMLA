//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT68), .A2(G116), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT68), .A2(G116), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT69), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(KEYINPUT69), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n191), .B1(new_n195), .B2(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT70), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT2), .B(G113), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n191), .B(new_n199), .C1(new_n195), .C2(new_n190), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n196), .A2(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(G137), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n204), .B(new_n209), .C1(new_n205), .C2(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G131), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(new_n213), .A3(new_n208), .A4(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT65), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G143), .B(G146), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT0), .A4(G128), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n220), .A2(new_n221), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n222), .A2(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n215), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n208), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n205), .A2(G137), .ZN(new_n232));
  OAI21_X1  g046(.A(G131), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n214), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n218), .B(G146), .C1(new_n235), .C2(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n216), .A3(G143), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G128), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n236), .B(new_n237), .C1(new_n220), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n230), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n203), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n240), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n234), .B2(KEYINPUT67), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n214), .A2(new_n233), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n245), .A2(new_n248), .B1(new_n215), .B2(new_n229), .ZN(new_n249));
  MUX2_X1   g063(.A(new_n249), .B(new_n242), .S(KEYINPUT30), .Z(new_n250));
  AOI21_X1  g064(.A(new_n243), .B1(new_n250), .B2(new_n203), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(G101), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT71), .A2(G237), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT71), .A2(G237), .ZN(new_n256));
  AOI21_X1  g070(.A(G953), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n253), .B(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n251), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT29), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n243), .A2(new_n262), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n203), .A2(new_n242), .A3(KEYINPUT28), .ZN(new_n264));
  INV_X1    g078(.A(new_n203), .ZN(new_n265));
  OAI22_X1  g079(.A1(new_n263), .A2(new_n264), .B1(new_n265), .B2(new_n249), .ZN(new_n266));
  INV_X1    g080(.A(new_n259), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n261), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n263), .A2(new_n264), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n230), .A2(new_n241), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n269), .A2(KEYINPUT29), .A3(new_n259), .A4(new_n272), .ZN(new_n273));
  OR2_X1    g087(.A1(new_n273), .A2(KEYINPUT72), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(KEYINPUT72), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n268), .A2(new_n274), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G472), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n266), .A2(new_n267), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n270), .A2(KEYINPUT30), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n280), .B(new_n203), .C1(new_n249), .C2(KEYINPUT30), .ZN(new_n281));
  INV_X1    g095(.A(new_n243), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n259), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT31), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n281), .A2(new_n285), .A3(new_n282), .A4(new_n259), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n279), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n288), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT32), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n278), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n187), .A2(G128), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT73), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n235), .A2(G119), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT24), .B(G110), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n295), .A2(KEYINPUT75), .A3(KEYINPUT23), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n297), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n235), .A2(KEYINPUT23), .A3(G119), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT74), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n300), .B1(new_n308), .B2(G110), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G140), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n311), .A3(KEYINPUT76), .ZN(new_n315));
  OR3_X1    g129(.A1(new_n310), .A2(KEYINPUT76), .A3(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n312), .B1(new_n317), .B2(KEYINPUT16), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G146), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n314), .A2(new_n311), .A3(KEYINPUT77), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT77), .B1(new_n314), .B2(new_n311), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n216), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n309), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n318), .B(G146), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n308), .A2(G110), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(new_n298), .C2(new_n299), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n309), .A2(KEYINPUT78), .A3(new_n319), .A4(new_n322), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT22), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(G137), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(KEYINPUT79), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n330), .B2(new_n335), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n325), .A2(new_n328), .A3(new_n329), .A4(new_n334), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  OAI22_X1  g157(.A1(new_n337), .A2(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n294), .B1(new_n344), .B2(G902), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n336), .B(KEYINPUT79), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n340), .B(new_n341), .ZN(new_n347));
  INV_X1    g161(.A(new_n294), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n346), .A2(new_n275), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n345), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G217), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(G234), .B2(new_n275), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(G902), .ZN(new_n355));
  XOR2_X1   g169(.A(new_n355), .B(KEYINPUT82), .Z(new_n356));
  NAND3_X1  g170(.A1(new_n346), .A2(new_n356), .A3(new_n347), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n293), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G122), .ZN(new_n362));
  XOR2_X1   g176(.A(KEYINPUT83), .B(G101), .Z(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G107), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G104), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT3), .B1(new_n364), .B2(G107), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n363), .A2(new_n365), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n368), .A3(new_n365), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G101), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n372), .A3(KEYINPUT4), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n372), .A2(KEYINPUT4), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n203), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n367), .A2(G104), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n365), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G101), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n365), .B2(new_n377), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT84), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n370), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT5), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n197), .B2(new_n200), .ZN(new_n386));
  OAI21_X1  g200(.A(G113), .B1(new_n194), .B2(KEYINPUT5), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n202), .B(new_n384), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  AOI211_X1 g202(.A(KEYINPUT89), .B(new_n362), .C1(new_n375), .C2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n375), .A2(new_n388), .A3(new_n362), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT6), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT89), .B1(new_n375), .B2(new_n388), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n394));
  INV_X1    g208(.A(new_n362), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  MUX2_X1   g210(.A(new_n240), .B(new_n229), .S(G125), .Z(new_n397));
  INV_X1    g211(.A(G224), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G953), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n397), .B(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n392), .A2(KEYINPUT90), .A3(new_n396), .A4(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT90), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n396), .B1(new_n389), .B2(new_n391), .ZN(new_n404));
  INV_X1    g218(.A(new_n401), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n397), .B1(KEYINPUT92), .B2(new_n400), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT7), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n407), .B1(new_n408), .B2(new_n399), .ZN(new_n409));
  INV_X1    g223(.A(new_n387), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n196), .B2(new_n385), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n202), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n384), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n362), .B(KEYINPUT91), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT8), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n202), .B1(new_n386), .B2(new_n387), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n413), .B(new_n415), .C1(new_n416), .C2(new_n384), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT7), .B(new_n400), .C1(new_n397), .C2(KEYINPUT92), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n409), .A2(new_n417), .A3(new_n390), .A4(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n419), .A2(new_n275), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n402), .A2(new_n406), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n402), .A2(new_n406), .A3(new_n422), .A4(new_n420), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(KEYINPUT93), .A3(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n425), .A2(KEYINPUT93), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n318), .B(new_n216), .ZN(new_n429));
  AND2_X1   g243(.A1(KEYINPUT71), .A2(G237), .ZN(new_n430));
  OAI211_X1 g244(.A(G214), .B(new_n331), .C1(new_n430), .C2(new_n254), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n218), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT71), .B(G237), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(G143), .A3(G214), .A4(new_n331), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n213), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT17), .ZN(new_n436));
  INV_X1    g250(.A(new_n435), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n434), .A3(new_n213), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n429), .B(new_n436), .C1(KEYINPUT17), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT18), .A2(G131), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n432), .A2(new_n434), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n314), .A2(new_n311), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT77), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n314), .A2(new_n311), .A3(KEYINPUT77), .ZN(new_n447));
  AOI21_X1  g261(.A(G146), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n315), .A2(G146), .A3(new_n316), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT18), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n451), .B(new_n213), .C1(new_n432), .C2(new_n434), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n441), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n322), .B1(new_n216), .B2(new_n317), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT94), .A4(new_n443), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(G113), .B(G122), .Z(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT96), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n364), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n440), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT19), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n320), .B2(new_n321), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT19), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n216), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n319), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n439), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n457), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT95), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n453), .A2(new_n456), .B1(new_n466), .B2(new_n439), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT95), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n461), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(G475), .A2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT20), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n472), .ZN(new_n477));
  INV_X1    g291(.A(new_n460), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n471), .B2(KEYINPUT95), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n440), .A2(new_n457), .ZN(new_n480));
  OAI22_X1  g294(.A1(new_n477), .A2(new_n479), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n474), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT97), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n476), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n481), .A2(KEYINPUT97), .A3(new_n482), .A4(new_n474), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n331), .A2(G952), .ZN(new_n488));
  NAND2_X1  g302(.A1(G234), .A2(G237), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT21), .B(G898), .Z(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(G902), .A3(G953), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT9), .B(G234), .Z(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n495), .A2(new_n352), .A3(G953), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT68), .B(G116), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G122), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n192), .A2(G122), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n367), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G128), .B(G143), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(G134), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT14), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n498), .B2(G122), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n506), .B1(new_n508), .B2(new_n500), .ZN(new_n509));
  INV_X1    g323(.A(G122), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n188), .B2(new_n189), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n507), .ZN(new_n512));
  OAI211_X1 g326(.A(KEYINPUT98), .B(new_n501), .C1(new_n511), .C2(new_n507), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI211_X1 g328(.A(new_n503), .B(new_n505), .C1(new_n514), .C2(G107), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n499), .A2(new_n501), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G107), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n517), .A2(new_n502), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n504), .A2(new_n205), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n504), .A2(KEYINPUT13), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n218), .A2(G128), .ZN(new_n521));
  OAI21_X1  g335(.A(G134), .B1(new_n521), .B2(KEYINPUT13), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n519), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n497), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n514), .A2(G107), .ZN(new_n526));
  INV_X1    g340(.A(new_n505), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n502), .A3(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n518), .A2(new_n523), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n496), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n275), .ZN(new_n532));
  INV_X1    g346(.A(G478), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n532), .B(new_n534), .Z(new_n535));
  XNOR2_X1  g349(.A(new_n480), .B(new_n460), .ZN(new_n536));
  OAI21_X1  g350(.A(G475), .B1(new_n536), .B2(G902), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n487), .A2(new_n493), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G214), .B1(G237), .B2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n428), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G221), .B1(new_n495), .B2(G902), .ZN(new_n543));
  XNOR2_X1  g357(.A(G110), .B(G140), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n331), .A2(G227), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n215), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT10), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n244), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n384), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n220), .A2(KEYINPUT1), .A3(new_n235), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n236), .A2(KEYINPUT85), .A3(new_n237), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT85), .B1(new_n236), .B2(new_n237), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n549), .B1(new_n555), .B2(new_n383), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n229), .A2(new_n374), .A3(new_n373), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT86), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT86), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n551), .A2(new_n556), .A3(new_n560), .A4(new_n557), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n548), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n556), .A2(new_n548), .A3(new_n557), .A4(new_n551), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n547), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n383), .A2(new_n244), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n383), .B2(new_n555), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n215), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n563), .A2(new_n546), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(G902), .B1(new_n565), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G469), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n275), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n546), .B1(new_n570), .B2(new_n563), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n562), .A2(new_n571), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT87), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n568), .A2(new_n569), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT12), .B1(new_n567), .B2(new_n215), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n563), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n547), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT87), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n586), .B(new_n587), .C1(new_n562), .C2(new_n571), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n575), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n543), .B1(new_n579), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT88), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n361), .A2(new_n542), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n593), .B(new_n363), .Z(G3));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n287), .A2(new_n275), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n287), .B2(new_n275), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n592), .A2(new_n359), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n541), .B1(new_n424), .B2(new_n425), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n493), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n533), .A2(G902), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n525), .A2(new_n604), .A3(new_n530), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n604), .B1(new_n525), .B2(new_n530), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n532), .A2(new_n533), .ZN(new_n610));
  OAI211_X1 g424(.A(KEYINPUT100), .B(new_n603), .C1(new_n605), .C2(new_n606), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT101), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n485), .A2(new_n486), .A3(new_n537), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n602), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n600), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(new_n535), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n476), .A2(new_n483), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n537), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n602), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n600), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n330), .B(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n356), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n351), .B2(new_n353), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n542), .A2(new_n592), .A3(new_n599), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT37), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G110), .ZN(G12));
  AND2_X1   g451(.A1(new_n634), .A2(new_n601), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n492), .A2(G900), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n490), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n625), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n638), .A2(new_n293), .A3(new_n592), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  AND3_X1   g458(.A1(new_n617), .A2(new_n540), .A3(new_n623), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n633), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT103), .Z(new_n647));
  AND2_X1   g461(.A1(new_n428), .A2(KEYINPUT38), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n428), .A2(KEYINPUT38), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n251), .A2(new_n267), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n282), .A2(new_n267), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n275), .B1(new_n653), .B2(new_n271), .ZN(new_n654));
  OAI21_X1  g468(.A(G472), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n292), .A2(new_n289), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT102), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n640), .B(KEYINPUT39), .Z(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n592), .A2(KEYINPUT40), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(KEYINPUT40), .B1(new_n592), .B2(new_n659), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n651), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n218), .ZN(G45));
  NOR2_X1   g478(.A1(new_n618), .A2(new_n641), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n638), .A2(new_n293), .A3(new_n592), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  OR2_X1    g481(.A1(new_n574), .A2(new_n575), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n543), .A3(new_n576), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n360), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n619), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT41), .B(G113), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n626), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G116), .ZN(G18));
  INV_X1    g489(.A(new_n539), .ZN(new_n676));
  INV_X1    g490(.A(new_n669), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n638), .A2(new_n293), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G119), .ZN(G21));
  AND2_X1   g493(.A1(new_n269), .A2(new_n272), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n284), .B(new_n286), .C1(new_n680), .C2(new_n259), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n287), .A2(new_n275), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(G472), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n288), .A2(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n359), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n424), .A2(new_n425), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n645), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n685), .A2(new_n493), .A3(new_n677), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G122), .ZN(G24));
  NAND4_X1  g503(.A1(new_n638), .A2(new_n665), .A3(new_n677), .A4(new_n684), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G125), .ZN(G27));
  AOI21_X1  g505(.A(new_n541), .B1(new_n426), .B2(new_n427), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n580), .A2(new_n581), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n579), .B1(G469), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n543), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n692), .A2(KEYINPUT105), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT105), .B1(new_n692), .B2(new_n696), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n361), .B(new_n665), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n692), .A2(new_n696), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n692), .A2(KEYINPUT105), .A3(new_n696), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n289), .A2(KEYINPUT106), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n289), .A2(KEYINPUT106), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n278), .A2(new_n292), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n359), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n706), .A2(KEYINPUT42), .A3(new_n665), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n701), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G131), .ZN(G33));
  INV_X1    g528(.A(new_n642), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n360), .B(new_n715), .C1(new_n704), .C2(new_n705), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n205), .ZN(G36));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n617), .B1(new_n614), .B2(new_n615), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n485), .A2(new_n486), .A3(new_n537), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n616), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(KEYINPUT110), .A3(KEYINPUT43), .ZN(new_n724));
  INV_X1    g538(.A(new_n632), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n599), .B1(new_n354), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n721), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n721), .A2(new_n724), .A3(KEYINPUT44), .A4(new_n726), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n732), .A2(new_n692), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n727), .A2(KEYINPUT111), .A3(new_n728), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT112), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n582), .A2(new_n588), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n575), .B1(new_n693), .B2(KEYINPUT45), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n740), .B1(new_n738), .B2(new_n739), .ZN(new_n742));
  OAI211_X1 g556(.A(KEYINPUT46), .B(new_n578), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n576), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n578), .B1(new_n741), .B2(new_n742), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n747), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n743), .A2(KEYINPUT108), .A3(new_n576), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n746), .A2(new_n750), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n754), .A2(new_n543), .A3(new_n659), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n731), .A2(new_n733), .A3(new_n756), .A4(new_n734), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n736), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  INV_X1    g573(.A(new_n692), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n760), .A2(new_n359), .A3(new_n293), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n754), .A2(new_n543), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n762), .B1(new_n754), .B2(new_n543), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n665), .B(new_n761), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  INV_X1    g580(.A(new_n650), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n657), .A2(new_n358), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n723), .A2(new_n695), .A3(new_n541), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n668), .A2(new_n576), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT49), .Z(new_n771));
  NAND4_X1  g585(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n716), .B1(new_n701), .B2(new_n712), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n428), .A2(new_n541), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n618), .B1(new_n535), .B2(new_n617), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n600), .A2(new_n774), .A3(new_n493), .A4(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(new_n635), .A3(new_n593), .A4(new_n678), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n671), .A2(new_n674), .A3(new_n688), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n633), .A2(new_n641), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n618), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(new_n684), .C1(new_n697), .C2(new_n698), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n538), .A2(new_n624), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n692), .A2(new_n592), .A3(new_n293), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n781), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n773), .A2(new_n779), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n633), .A2(new_n640), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n657), .A2(new_n687), .A3(new_n696), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n643), .A2(new_n666), .A3(new_n690), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n791), .B(KEYINPUT114), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n643), .A2(new_n666), .A3(new_n690), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT52), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(KEYINPUT115), .A3(new_n798), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n788), .A2(new_n801), .A3(KEYINPUT53), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n786), .A2(new_n777), .A3(new_n778), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n773), .ZN(new_n806));
  INV_X1    g620(.A(new_n799), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n803), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  AND4_X1   g625(.A1(KEYINPUT53), .A2(new_n799), .A3(new_n805), .A4(new_n773), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n788), .A2(new_n801), .A3(new_n802), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n812), .B1(new_n813), .B2(new_n804), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n763), .A2(new_n764), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n543), .B2(new_n770), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n490), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n685), .A2(new_n821), .A3(new_n724), .A4(new_n721), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n760), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n818), .A2(new_n819), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n822), .A2(new_n669), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n541), .A3(new_n767), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT50), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n760), .A2(new_n490), .A3(new_n669), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n634), .A2(new_n684), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n724), .A2(new_n829), .A3(new_n721), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n768), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n832), .A2(new_n616), .A3(new_n617), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n828), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n825), .A2(KEYINPUT51), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n818), .A2(new_n823), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT51), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n829), .A2(new_n711), .A3(new_n724), .A4(new_n721), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT48), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n829), .A2(new_n782), .A3(new_n768), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n826), .A2(new_n601), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n488), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n816), .A2(new_n835), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(G952), .A2(G953), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n772), .B1(new_n843), .B2(new_n844), .ZN(G75));
  NOR2_X1   g659(.A1(new_n331), .A2(G952), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n275), .B1(new_n803), .B2(new_n808), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT56), .B1(new_n848), .B2(G210), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n848), .A2(G210), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n404), .B(KEYINPUT118), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT55), .Z(new_n856));
  XOR2_X1   g670(.A(KEYINPUT119), .B(KEYINPUT120), .Z(new_n857));
  XNOR2_X1  g671(.A(new_n401), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n856), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n859), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n849), .A2(new_n850), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n851), .B1(new_n860), .B2(new_n862), .ZN(G51));
  NAND2_X1  g677(.A1(new_n565), .A2(new_n573), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n578), .A2(KEYINPUT57), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n803), .A2(new_n810), .A3(new_n808), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n810), .B1(new_n803), .B2(new_n808), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n578), .A2(KEYINPUT57), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n741), .A2(new_n742), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n848), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n846), .B1(new_n870), .B2(new_n872), .ZN(G54));
  NAND3_X1  g687(.A1(new_n848), .A2(KEYINPUT58), .A3(G475), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n874), .A2(new_n473), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n473), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n875), .A2(new_n876), .A3(new_n846), .ZN(G60));
  OR2_X1    g691(.A1(new_n605), .A2(new_n606), .ZN(new_n878));
  NAND2_X1  g692(.A1(G478), .A2(G902), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT59), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n878), .B1(new_n816), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n866), .A2(new_n867), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n880), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n881), .A2(new_n884), .A3(new_n846), .ZN(G63));
  NAND2_X1  g699(.A1(new_n803), .A2(new_n808), .ZN(new_n886));
  NAND2_X1  g700(.A1(G217), .A2(G902), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT60), .Z(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n344), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n631), .A3(new_n888), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n847), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n890), .A2(KEYINPUT61), .A3(new_n847), .A4(new_n891), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(G66));
  INV_X1    g710(.A(new_n491), .ZN(new_n897));
  OAI21_X1  g711(.A(G953), .B1(new_n897), .B2(new_n398), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n779), .B2(G953), .ZN(new_n899));
  INV_X1    g713(.A(G898), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n855), .B1(new_n900), .B2(G953), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n899), .B(new_n901), .Z(G69));
  NAND2_X1  g716(.A1(new_n463), .A2(new_n464), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n250), .B(new_n903), .Z(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT122), .ZN(new_n905));
  INV_X1    g719(.A(new_n765), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n797), .B(KEYINPUT62), .C1(new_n651), .C2(new_n662), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n663), .B2(new_n794), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n361), .A2(new_n775), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(new_n592), .A3(new_n659), .A4(new_n692), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n758), .A2(KEYINPUT123), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT123), .B1(new_n758), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n905), .B1(new_n915), .B2(new_n331), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n765), .A2(new_n713), .A3(new_n797), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n709), .A2(new_n687), .A3(new_n359), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n754), .A2(new_n918), .A3(new_n543), .A4(new_n659), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(KEYINPUT124), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(KEYINPUT124), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n716), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n917), .A2(new_n331), .A3(new_n758), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(G900), .A2(G953), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n904), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT125), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n924), .A3(new_n904), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n758), .A2(new_n912), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n758), .A2(KEYINPUT123), .A3(new_n912), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(G953), .B1(new_n933), .B2(new_n910), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n927), .B(new_n928), .C1(new_n934), .C2(new_n905), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n331), .B1(G227), .B2(G900), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n926), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n926), .B2(new_n935), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G72));
  NAND4_X1  g753(.A1(new_n917), .A2(new_n758), .A3(new_n779), .A4(new_n922), .ZN(new_n940));
  NAND2_X1  g754(.A1(G472), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT63), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n940), .A2(new_n945), .A3(new_n942), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n944), .A2(new_n267), .A3(new_n251), .A4(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n283), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n942), .B1(new_n260), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT127), .Z(new_n950));
  OAI211_X1 g764(.A(new_n947), .B(new_n847), .C1(new_n814), .C2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n933), .A2(new_n779), .A3(new_n910), .ZN(new_n952));
  AOI211_X1 g766(.A(new_n267), .B(new_n251), .C1(new_n952), .C2(new_n942), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(G57));
endmodule


