//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(KEYINPUT69), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n476), .A3(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n477), .A2(G137), .A3(new_n478), .A4(new_n467), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT69), .B(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n473), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n477), .A2(new_n467), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n478), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n467), .A2(new_n469), .A3(new_n478), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n494), .A2(new_n496), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n477), .A2(new_n478), .A3(new_n467), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n477), .A2(new_n467), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT70), .A2(G114), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT70), .A2(G114), .ZN(new_n504));
  OAI21_X1  g079(.A(G2105), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT71), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n502), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n500), .B1(new_n510), .B2(new_n512), .ZN(G164));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT72), .B(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT5), .B(G543), .Z(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT73), .B(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT72), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT72), .A2(G651), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT6), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n514), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G50), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G62), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n517), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(new_n515), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n520), .A2(new_n527), .A3(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT75), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n536));
  XNOR2_X1  g111(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n518), .A2(G89), .ZN(new_n538));
  INV_X1    g113(.A(new_n517), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n526), .A2(G51), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n537), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n517), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n546), .A2(new_n515), .B1(new_n526), .B2(G52), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n518), .A2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n517), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(new_n515), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n518), .A2(G81), .B1(G43), .B2(new_n526), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n555), .A2(KEYINPUT76), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(KEYINPUT76), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n517), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n524), .A2(new_n525), .ZN(new_n570));
  AND4_X1   g145(.A1(new_n569), .A2(new_n570), .A3(G53), .A4(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n569), .B1(new_n526), .B2(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n574), .B1(new_n516), .B2(new_n517), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n539), .A3(KEYINPUT77), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(G91), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n575), .A2(KEYINPUT78), .A3(new_n576), .A4(G91), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n573), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT79), .ZN(G299));
  NAND3_X1  g157(.A1(new_n575), .A2(G87), .A3(new_n576), .ZN(new_n583));
  INV_X1    g158(.A(G651), .ZN(new_n584));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n584), .B1(new_n517), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(G49), .B2(new_n526), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT80), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n583), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G288));
  NAND3_X1  g168(.A1(new_n575), .A2(G86), .A3(new_n576), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n517), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(new_n515), .B1(new_n526), .B2(G48), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n517), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n515), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n526), .A2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n570), .A2(new_n539), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n607), .A2(KEYINPUT81), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n607), .A2(KEYINPUT81), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n603), .B1(new_n608), .B2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n612));
  OAI21_X1  g187(.A(G54), .B1(new_n526), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g188(.A1(new_n516), .A2(KEYINPUT82), .A3(new_n521), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n539), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n615));
  OAI22_X1  g190(.A1(new_n613), .A2(new_n614), .B1(new_n615), .B2(new_n584), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n575), .A2(new_n576), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G92), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n617), .A2(KEYINPUT10), .A3(G92), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n611), .B1(new_n622), .B2(G868), .ZN(G284));
  XNOR2_X1  g198(.A(G284), .B(KEYINPUT83), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n581), .B(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n625), .B1(new_n627), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n625), .B1(new_n627), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n622), .B1(new_n630), .B2(G860), .ZN(G148));
  OR2_X1    g206(.A1(new_n558), .A2(G868), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n622), .A2(new_n630), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT84), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n633), .B1(new_n635), .B2(G868), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g212(.A1(new_n495), .A2(new_n480), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n486), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n488), .A2(G123), .ZN(new_n643));
  OR2_X1    g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(G2104), .C1(G111), .C2(new_n478), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n641), .A2(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n652), .B(new_n658), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(G14), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n660), .ZN(G401));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT85), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT86), .Z(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n669), .B(KEYINPUT17), .Z(new_n673));
  INV_X1    g248(.A(new_n670), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n667), .B2(new_n669), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n676));
  OAI22_X1  g251(.A1(new_n673), .A2(new_n666), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n676), .B2(new_n675), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n667), .A2(new_n674), .ZN(new_n679));
  AOI211_X1 g254(.A(new_n672), .B(new_n678), .C1(new_n673), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2096), .B(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(new_n693), .B(new_n692), .S(new_n685), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(G229));
  NAND2_X1  g278(.A1(G301), .A2(G16), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G5), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G1961), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G168), .A2(new_n705), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n705), .B2(G21), .ZN(new_n711));
  INV_X1    g286(.A(G1966), .ZN(new_n712));
  OAI22_X1  g287(.A1(new_n711), .A2(new_n712), .B1(new_n707), .B2(new_n708), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n709), .B(new_n713), .C1(new_n712), .C2(new_n711), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NOR2_X1   g290(.A1(G164), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G27), .B2(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(G2078), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G34), .ZN(new_n721));
  AOI21_X1  g296(.A(G29), .B1(new_n721), .B2(KEYINPUT24), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(KEYINPUT24), .B2(new_n721), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n483), .B2(new_n715), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT31), .B(G11), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT99), .ZN(new_n729));
  INV_X1    g304(.A(G28), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n731));
  AOI21_X1  g306(.A(G29), .B1(new_n730), .B2(KEYINPUT30), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n727), .B(new_n733), .C1(new_n715), .C2(new_n646), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n720), .A2(new_n726), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n715), .A2(G33), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n486), .A2(G139), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT97), .Z(new_n741));
  INV_X1    g316(.A(new_n470), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n742), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n478), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n736), .B1(new_n745), .B2(new_n715), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G2072), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n714), .A2(new_n719), .A3(new_n735), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n715), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n715), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT29), .Z(new_n751));
  INV_X1    g326(.A(G2090), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G1348), .ZN(new_n754));
  NOR2_X1   g329(.A1(G4), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n622), .B2(G16), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n753), .A2(KEYINPUT100), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(KEYINPUT100), .B2(new_n753), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n715), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n486), .A2(G141), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n488), .A2(G129), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT26), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n481), .A2(G105), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n761), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n760), .B1(new_n769), .B2(new_n715), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT27), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1996), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n754), .B2(new_n757), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n748), .A2(new_n759), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n751), .A2(new_n752), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G19), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n559), .B2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n775), .B1(G1341), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n715), .A2(G26), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT28), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n486), .A2(G140), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n488), .A2(G128), .ZN(new_n782));
  OR2_X1    g357(.A1(G104), .A2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n783), .B(G2104), .C1(G116), .C2(new_n478), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT95), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n780), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT96), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G2067), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n778), .B(new_n792), .C1(G1341), .C2(new_n777), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(G2067), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n746), .A2(G2072), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT98), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n705), .A2(G20), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT23), .Z(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G299), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1956), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n774), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G23), .B(new_n588), .S(G16), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT92), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT33), .B(G1976), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n804), .A2(new_n806), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n705), .A2(G22), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT93), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G303), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1971), .Z(new_n812));
  AND2_X1   g387(.A1(new_n705), .A2(G6), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G305), .B2(G16), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT32), .B(G1981), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n814), .A2(new_n816), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n812), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n807), .A2(new_n808), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT94), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT34), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(G290), .A2(KEYINPUT91), .ZN(new_n824));
  NAND2_X1  g399(.A1(G290), .A2(KEYINPUT91), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n705), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G24), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n705), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1986), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n715), .A2(G25), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n486), .A2(G131), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT90), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n478), .A2(G107), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n488), .A2(G119), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n830), .B1(new_n838), .B2(new_n715), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT35), .B(G1991), .Z(new_n840));
  XOR2_X1   g415(.A(new_n839), .B(new_n840), .Z(new_n841));
  NOR2_X1   g416(.A1(new_n829), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n821), .A2(new_n822), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n823), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n823), .A2(new_n842), .A3(new_n846), .A4(new_n843), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n802), .B1(new_n845), .B2(new_n847), .ZN(G311));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n847), .ZN(new_n849));
  INV_X1    g424(.A(new_n802), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(G150));
  NAND2_X1  g426(.A1(new_n622), .A2(G559), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT38), .Z(new_n853));
  NAND2_X1  g428(.A1(G80), .A2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G67), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n517), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n515), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n526), .A2(G55), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n605), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n558), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n863), .B(new_n554), .C1(new_n557), .C2(new_n556), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n853), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g445(.A(G860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n864), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT102), .ZN(G145));
  XNOR2_X1  g451(.A(new_n837), .B(new_n639), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n769), .B1(new_n787), .B2(new_n788), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n486), .A2(G142), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n488), .A2(G130), .ZN(new_n881));
  OR2_X1    g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n882), .B(G2104), .C1(G118), .C2(new_n478), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n787), .A2(new_n788), .A3(new_n769), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n884), .ZN(new_n887));
  INV_X1    g462(.A(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n888), .B2(new_n878), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n877), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n877), .B1(new_n889), .B2(new_n886), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n745), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n886), .A2(new_n889), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n837), .B(new_n639), .Z(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n745), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n890), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n500), .A2(new_n509), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n492), .B(G160), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT103), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n646), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n893), .A2(new_n898), .A3(new_n900), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n905), .B1(new_n902), .B2(new_n906), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT104), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n902), .A2(new_n906), .ZN(new_n912));
  INV_X1    g487(.A(new_n905), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n907), .A4(new_n908), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n911), .A2(new_n916), .A3(new_n918), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(G395));
  XNOR2_X1  g497(.A(new_n635), .B(new_n868), .ZN(new_n923));
  NAND2_X1  g498(.A1(G299), .A2(new_n622), .ZN(new_n924));
  INV_X1    g499(.A(new_n622), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n627), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n926), .A3(KEYINPUT41), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT41), .B1(new_n924), .B2(new_n926), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n923), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n926), .A3(KEYINPUT106), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n926), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n923), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n588), .B(KEYINPUT107), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G303), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n588), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(G166), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(G290), .A2(new_n594), .A3(new_n598), .ZN(new_n942));
  OAI211_X1 g517(.A(G305), .B(new_n603), .C1(new_n608), .C2(new_n609), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n937), .A2(new_n940), .A3(new_n943), .A4(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(KEYINPUT108), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  AND4_X1   g529(.A1(new_n930), .A2(new_n935), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n930), .A2(new_n935), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G868), .B2(new_n863), .ZN(G295));
  OAI21_X1  g533(.A(new_n957), .B1(G868), .B2(new_n863), .ZN(G331));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  XNOR2_X1  g537(.A(G171), .B(G286), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n865), .A2(new_n963), .A3(new_n866), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n865), .B2(new_n866), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT109), .B1(new_n868), .B2(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n928), .B2(new_n929), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n964), .A2(new_n965), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n932), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n951), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n908), .ZN(new_n973));
  INV_X1    g548(.A(new_n968), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n934), .A2(new_n931), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI22_X1  g551(.A1(new_n928), .A2(new_n929), .B1(new_n965), .B2(new_n964), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n951), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n961), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n968), .B1(new_n931), .B2(new_n934), .ZN(new_n980));
  INV_X1    g555(.A(new_n929), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n970), .B1(new_n981), .B2(new_n927), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n950), .B(new_n949), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n983), .A2(KEYINPUT110), .A3(new_n908), .A4(new_n972), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n960), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n969), .A2(new_n971), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n951), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n973), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT43), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT44), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT43), .B1(new_n987), .B2(new_n973), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n960), .A3(new_n983), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n991), .A2(new_n996), .ZN(G397));
  OAI211_X1 g572(.A(KEYINPUT113), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n473), .A2(G40), .A3(new_n482), .A4(new_n479), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n497), .A2(new_n499), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n502), .A2(new_n511), .A3(new_n508), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n511), .B1(new_n502), .B2(new_n508), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1001), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1001), .B(new_n1006), .C1(new_n500), .C2(new_n509), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT113), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n998), .B(new_n1000), .C1(new_n1007), .C2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT114), .B1(new_n1011), .B2(G2090), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n999), .B1(new_n1014), .B2(new_n1009), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n752), .A4(new_n998), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT111), .B(G1384), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT45), .B(new_n1018), .C1(new_n500), .C2(new_n509), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1000), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1012), .B(new_n1017), .C1(G1971), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G303), .A2(G8), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1023), .A2(G8), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1006), .B1(new_n500), .B2(new_n509), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(new_n999), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n588), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT52), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n518), .A2(G86), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n598), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G1981), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n594), .A2(new_n1042), .A3(new_n598), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1041), .A2(KEYINPUT49), .A3(new_n1043), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1035), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1038), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n592), .B2(G1976), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1037), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1049), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1031), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1014), .A2(new_n1009), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1057), .A2(new_n725), .A3(new_n1000), .A4(new_n998), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n999), .B1(new_n1032), .B2(new_n1021), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n712), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1034), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1023), .A2(G8), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1030), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1056), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1061), .B1(new_n1011), .B2(G2084), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G8), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G286), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1022), .A2(G1971), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n999), .B1(new_n1032), .B2(KEYINPUT50), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(G2090), .ZN(new_n1074));
  OAI21_X1  g649(.A(G8), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1065), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1031), .A2(new_n1055), .A3(new_n1070), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT63), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1067), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1055), .A2(G8), .A3(new_n1023), .A4(new_n1030), .ZN(new_n1082));
  AOI211_X1 g657(.A(G1976), .B(G288), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1043), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1035), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT117), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1082), .A2(KEYINPUT117), .A3(new_n1085), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1080), .B(new_n1081), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1086), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1056), .A2(new_n1066), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT118), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1011), .A2(new_n708), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1000), .A2(new_n1019), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G164), .A2(G1384), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(KEYINPUT45), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1093), .B1(new_n1096), .B2(G2078), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n718), .A2(KEYINPUT53), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1092), .B(new_n1097), .C1(new_n1060), .C2(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n579), .A2(new_n580), .ZN(new_n1103));
  INV_X1    g678(.A(new_n573), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n1106));
  INV_X1    g681(.A(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1073), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n581), .B2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(G2072), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1094), .B(new_n1113), .C1(new_n1095), .C2(KEYINPUT45), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1106), .A2(new_n1108), .A3(new_n1111), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1011), .A2(new_n754), .ZN(new_n1116));
  INV_X1    g691(.A(G2067), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1033), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n925), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1111), .A2(new_n1106), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1115), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  AND4_X1   g697(.A1(new_n1108), .A2(new_n1106), .A3(new_n1114), .A4(new_n1111), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(new_n1120), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1116), .A2(new_n925), .A3(KEYINPUT60), .A4(new_n1118), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1108), .A2(new_n1114), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(KEYINPUT61), .A3(new_n1115), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1096), .A2(G1996), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT58), .B(G1341), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1033), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1130), .B(new_n559), .C1(new_n1131), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1996), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1133), .B1(new_n1022), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT59), .B1(new_n1136), .B2(new_n558), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1124), .A2(new_n1125), .A3(new_n1129), .A4(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1116), .A2(KEYINPUT60), .A3(new_n1118), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT60), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n925), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1121), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G301), .B(KEYINPUT54), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT45), .B1(new_n901), .B2(new_n1018), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(new_n1098), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1144), .B1(new_n1146), .B2(new_n1094), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1097), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1149), .B2(new_n1092), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1011), .A2(KEYINPUT125), .A3(new_n708), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1150), .A2(new_n1151), .B1(new_n1099), .B2(new_n1144), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1102), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(G286), .A2(G8), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT121), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1154), .A2(KEYINPUT121), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1069), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1062), .A2(KEYINPUT123), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT51), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1068), .A2(new_n1158), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1068), .A2(KEYINPUT122), .A3(G8), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT51), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1062), .A2(KEYINPUT122), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT124), .B1(new_n1162), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT51), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1165), .B1(new_n1062), .B2(KEYINPUT123), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1069), .A2(new_n1159), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1069), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1178), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1175), .A2(new_n1176), .A3(new_n1163), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1171), .A2(new_n1180), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1153), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1100), .A2(KEYINPUT62), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1171), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1056), .A2(new_n1076), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1088), .B(new_n1091), .C1(new_n1182), .C2(new_n1186), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1145), .A2(new_n1000), .ZN(new_n1188));
  INV_X1    g763(.A(G290), .ZN(new_n1189));
  INV_X1    g764(.A(G1986), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT112), .Z(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(new_n1190), .B2(new_n1189), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n789), .B(new_n1117), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n768), .B(new_n1135), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n837), .B(new_n840), .Z(new_n1197));
  NOR2_X1   g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1188), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1187), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1188), .A2(new_n1135), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT46), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT126), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1188), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1206), .B1(new_n1194), .B2(new_n769), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1207), .B1(new_n1203), .B2(new_n1202), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT47), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT48), .ZN(new_n1211));
  OR3_X1    g786(.A1(new_n1192), .A2(new_n1211), .A3(new_n1206), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1211), .B1(new_n1192), .B2(new_n1206), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1212), .B(new_n1213), .C1(new_n1206), .C2(new_n1198), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n838), .A2(new_n840), .ZN(new_n1215));
  OAI22_X1  g790(.A1(new_n1196), .A2(new_n1215), .B1(G2067), .B2(new_n789), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n1188), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1210), .A2(new_n1214), .A3(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT127), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1201), .A2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g795(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1222));
  AND3_X1   g796(.A1(new_n917), .A2(new_n1222), .A3(new_n994), .ZN(G308));
  NAND3_X1  g797(.A1(new_n917), .A2(new_n1222), .A3(new_n994), .ZN(G225));
endmodule


