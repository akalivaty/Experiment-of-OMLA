//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT67), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT69), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n452), .B2(G2106), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT70), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n462), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(new_n470), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n462), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n477), .B1(new_n479), .B2(G124), .ZN(new_n480));
  INV_X1    g055(.A(new_n466), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G138), .B(new_n462), .C1(new_n469), .C2(new_n470), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(new_n462), .A3(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT71), .B1(new_n478), .B2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n487), .A2(new_n462), .A3(G138), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n465), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n486), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n479), .B2(G126), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n493), .B2(new_n498), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(G164));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT74), .Z(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT75), .B(G89), .Z(new_n523));
  OAI221_X1 g098(.A(new_n521), .B1(new_n508), .B2(new_n522), .C1(new_n506), .C2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n519), .A2(new_n524), .ZN(G168));
  NAND2_X1  g100(.A1(G77), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n503), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n514), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n533), .B1(new_n532), .B2(new_n531), .ZN(new_n534));
  AND2_X1   g109(.A1(KEYINPUT6), .A2(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT6), .A2(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n529), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(G90), .B1(new_n540), .B2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n514), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n538), .A2(G81), .B1(new_n540), .B2(G43), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(new_n506), .A2(KEYINPUT78), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT78), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n504), .A2(new_n505), .A3(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G91), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n540), .A2(KEYINPUT77), .A3(G53), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n508), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n558), .A2(new_n561), .A3(KEYINPUT9), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n514), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n557), .A2(new_n562), .A3(new_n563), .A4(new_n565), .ZN(G299));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G74), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n514), .B1(new_n529), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(G49), .B2(new_n540), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n553), .A2(G87), .A3(new_n555), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(G288));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  INV_X1    g148(.A(G73), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n574), .B2(new_n539), .ZN(new_n575));
  NAND3_X1  g150(.A1(KEYINPUT79), .A2(G73), .A3(G543), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n529), .C2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n540), .B2(G48), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n553), .A2(G86), .A3(new_n555), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n538), .A2(G85), .B1(new_n540), .B2(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n514), .B2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G54), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n586), .A2(new_n514), .B1(new_n587), .B2(new_n508), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n556), .A2(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n556), .A2(KEYINPUT10), .A3(G92), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n585), .B1(new_n593), .B2(G868), .ZN(G284));
  XOR2_X1   g169(.A(G284), .B(KEYINPUT80), .Z(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G168), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT81), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n599), .A2(KEYINPUT82), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(new_n599), .B2(KEYINPUT82), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(G297));
  OAI21_X1  g177(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(G280));
  INV_X1    g178(.A(new_n593), .ZN(new_n604));
  INV_X1    g179(.A(G860), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(G559), .B2(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT83), .Z(G148));
  OAI21_X1  g182(.A(KEYINPUT84), .B1(new_n547), .B2(G868), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n604), .A2(G559), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  MUX2_X1   g185(.A(KEYINPUT84), .B(new_n608), .S(new_n610), .Z(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n465), .A2(new_n463), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  INV_X1    g190(.A(G2100), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n479), .A2(G123), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n481), .A2(G135), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT85), .ZN(new_n621));
  NOR3_X1   g196(.A1(new_n621), .A2(new_n462), .A3(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n462), .B2(G111), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(G2104), .A3(new_n624), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n619), .B(new_n620), .C1(new_n622), .C2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n617), .A2(new_n618), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  INV_X1    g205(.A(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT86), .B(KEYINPUT14), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT87), .ZN(new_n645));
  INV_X1    g220(.A(G14), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n642), .B2(new_n643), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n645), .A2(new_n647), .ZN(G401));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT88), .B(G2100), .Z(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n652), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(new_n627), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(KEYINPUT90), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(KEYINPUT90), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n662), .A2(new_n663), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g248(.A(new_n673), .B(new_n672), .S(new_n668), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G229));
  NAND3_X1  g257(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT25), .Z(new_n684));
  INV_X1    g259(.A(G139), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n466), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT94), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(new_n462), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT95), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  MUX2_X1   g266(.A(G33), .B(new_n691), .S(G29), .Z(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(G2072), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT96), .Z(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G4), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n593), .B2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G1348), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(G20), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT23), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n599), .B2(new_n695), .ZN(new_n702));
  INV_X1    g277(.A(G1956), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n694), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G19), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n547), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT93), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(G1341), .Z(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G35), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G162), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G2090), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G27), .A2(G29), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G164), .B2(G29), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(G2078), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(G2078), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n709), .A2(new_n716), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n710), .A2(G32), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n463), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n479), .A2(G129), .ZN(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT26), .Z(new_n726));
  NAND3_X1  g301(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT97), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n722), .B1(new_n732), .B2(new_n710), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(G160), .A2(G29), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT24), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G34), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n710), .B1(new_n737), .B2(G34), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT30), .B(G28), .ZN(new_n744));
  OR2_X1    g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n744), .A2(new_n710), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n743), .B(new_n747), .C1(new_n710), .C2(new_n626), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n742), .B(new_n748), .C1(new_n692), .C2(G2072), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n695), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n695), .ZN(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n695), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n695), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(G1966), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(G1966), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n710), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n481), .A2(G140), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n479), .A2(G128), .ZN(new_n761));
  OR2_X1    g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n756), .A2(new_n757), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n735), .A2(new_n749), .A3(new_n753), .A4(new_n768), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n705), .A2(new_n721), .A3(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G6), .B(G305), .S(G16), .Z(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT32), .B(G1981), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n771), .B(new_n772), .Z(new_n773));
  AND2_X1   g348(.A1(new_n695), .A2(G22), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G303), .B2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G1971), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n695), .A2(G23), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n570), .A2(new_n571), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n695), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n775), .A2(new_n776), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n773), .A2(new_n777), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT34), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(KEYINPUT34), .ZN(new_n786));
  OR2_X1    g361(.A1(G95), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT91), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n481), .A2(G131), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n479), .A2(G119), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G29), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G25), .B2(G29), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT35), .B(G1991), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT92), .ZN(new_n798));
  MUX2_X1   g373(.A(G24), .B(G290), .S(G16), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1986), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n795), .A2(new_n796), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n785), .A2(new_n786), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n770), .A2(new_n805), .A3(new_n806), .ZN(G150));
  XOR2_X1   g382(.A(G150), .B(KEYINPUT99), .Z(G311));
  NAND2_X1  g383(.A1(new_n593), .A2(G559), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT102), .B(G93), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n538), .A2(new_n812), .B1(new_n540), .B2(G55), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT101), .B1(new_n814), .B2(new_n514), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n814), .A2(KEYINPUT101), .A3(new_n514), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(new_n547), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n811), .B(new_n819), .Z(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT103), .ZN(new_n822));
  AOI21_X1  g397(.A(G860), .B1(new_n820), .B2(KEYINPUT39), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n818), .A2(new_n605), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT37), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(G145));
  XNOR2_X1  g402(.A(new_n731), .B(new_n764), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n479), .A2(G130), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n462), .A2(G118), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G142), .B2(new_n481), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n828), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n493), .A2(new_n498), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT104), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n691), .B(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n792), .B(new_n614), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n834), .B(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n483), .B(G160), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n626), .ZN(new_n842));
  AOI21_X1  g417(.A(G37), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n840), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g420(.A(new_n596), .B1(new_n816), .B2(new_n817), .ZN(new_n846));
  XOR2_X1   g421(.A(G303), .B(G290), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n779), .B(G305), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n847), .B(new_n848), .Z(new_n849));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(KEYINPUT106), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(KEYINPUT106), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n851), .B(new_n852), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n609), .B(new_n819), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n593), .B(new_n599), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n855), .B(KEYINPUT41), .Z(new_n858));
  OAI211_X1 g433(.A(new_n857), .B(KEYINPUT105), .C1(new_n858), .C2(new_n854), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(KEYINPUT105), .B2(new_n857), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n853), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n846), .B1(new_n861), .B2(new_n596), .ZN(G295));
  OAI21_X1  g437(.A(new_n846), .B1(new_n861), .B2(new_n596), .ZN(G331));
  NAND2_X1  g438(.A1(G301), .A2(KEYINPUT107), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n819), .B(new_n864), .Z(new_n865));
  OAI21_X1  g440(.A(G168), .B1(G301), .B2(KEYINPUT107), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n819), .B(new_n864), .ZN(new_n868));
  INV_X1    g443(.A(new_n866), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT108), .B1(new_n871), .B2(new_n858), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n855), .A3(new_n870), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n849), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n849), .B1(new_n872), .B2(new_n873), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT43), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n872), .A2(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(new_n849), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n875), .A4(new_n874), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(KEYINPUT109), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n887));
  NAND3_X1  g462(.A1(new_n878), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(G397));
  NAND2_X1  g464(.A1(G160), .A2(G40), .ZN(new_n890));
  AOI21_X1  g465(.A(G1384), .B1(new_n493), .B2(new_n498), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT45), .ZN(new_n892));
  INV_X1    g467(.A(G1996), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT46), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n764), .B(new_n766), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n732), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n892), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n896), .B1(new_n732), .B2(new_n893), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(new_n893), .B2(new_n732), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n793), .A3(new_n796), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n764), .A2(G2067), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n898), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n792), .B(new_n796), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n892), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n898), .A2(G1986), .A3(G290), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(KEYINPUT48), .Z(new_n914));
  AOI21_X1  g489(.A(new_n909), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n903), .A2(new_n904), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G8), .ZN(new_n917));
  INV_X1    g492(.A(G40), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n468), .A2(new_n473), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n891), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1981), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n579), .A2(new_n580), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n575), .A2(new_n576), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n577), .B1(new_n502), .B2(new_n503), .ZN(new_n925));
  OAI21_X1  g500(.A(G651), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n540), .A2(G48), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n504), .A2(new_n505), .A3(G86), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G1981), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT49), .B1(new_n923), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n921), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n923), .A2(new_n930), .A3(KEYINPUT49), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n933), .A2(KEYINPUT113), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(KEYINPUT113), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1976), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n779), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n921), .B1(new_n938), .B2(new_n923), .ZN(new_n939));
  XNOR2_X1  g514(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(G166), .B2(new_n917), .ZN(new_n942));
  NAND3_X1  g517(.A1(G303), .A2(G8), .A3(new_n940), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n945), .B(G1384), .C1(new_n493), .C2(new_n498), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n499), .B2(new_n500), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n948), .B2(new_n945), .ZN(new_n949));
  AOI21_X1  g524(.A(G1971), .B1(new_n949), .B2(new_n919), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n890), .B1(new_n891), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n835), .A2(KEYINPUT72), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n493), .A2(new_n498), .A3(new_n494), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n713), .B(new_n952), .C1(new_n955), .C2(new_n951), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n944), .B(G8), .C1(new_n950), .C2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT52), .B1(G288), .B2(new_n937), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n570), .A2(new_n571), .A3(G1976), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n920), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT112), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n920), .A3(new_n964), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n920), .A2(new_n961), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT111), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n920), .A2(new_n969), .A3(new_n961), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n970), .A3(KEYINPUT52), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n966), .A2(new_n936), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n939), .B1(new_n959), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n944), .ZN(new_n974));
  INV_X1    g549(.A(new_n946), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n975), .B(new_n919), .C1(new_n955), .C2(KEYINPUT45), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n919), .B1(new_n891), .B2(new_n951), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n955), .B2(new_n951), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n976), .A2(new_n776), .B1(new_n978), .B2(new_n713), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n974), .B1(new_n979), .B2(new_n917), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n835), .A2(new_n947), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n890), .B1(new_n981), .B2(new_n945), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n948), .B2(new_n945), .ZN(new_n983));
  INV_X1    g558(.A(G1966), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n741), .B(new_n952), .C1(new_n955), .C2(new_n951), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n917), .B(G286), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n980), .A2(new_n972), .A3(new_n987), .A4(new_n958), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT63), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n985), .A2(new_n986), .ZN(new_n991));
  AND4_X1   g566(.A1(KEYINPUT63), .A2(new_n991), .A3(G8), .A4(G168), .ZN(new_n992));
  OAI21_X1  g567(.A(G8), .B1(new_n950), .B2(new_n957), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n974), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n958), .A2(new_n992), .A3(new_n994), .A4(new_n972), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n973), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n952), .B1(new_n955), .B2(new_n951), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n919), .B1(new_n891), .B2(KEYINPUT45), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n955), .B2(KEYINPUT45), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(G2078), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n752), .A2(new_n997), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1000), .B1(new_n976), .B2(G2078), .ZN(new_n1003));
  AOI21_X1  g578(.A(G301), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n980), .A2(new_n958), .A3(new_n972), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n985), .A2(G168), .A3(new_n986), .ZN(new_n1006));
  AND2_X1   g581(.A1(KEYINPUT119), .A2(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT51), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1010), .A3(new_n1007), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n991), .A2(G8), .A3(G286), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1004), .B(new_n1005), .C1(new_n1013), .C2(KEYINPUT62), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT122), .B1(new_n1013), .B2(KEYINPUT62), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n996), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n835), .A2(new_n951), .A3(new_n947), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n919), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(KEYINPUT50), .B2(new_n948), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT120), .B1(new_n1021), .B2(G1961), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n997), .A2(new_n1023), .A3(new_n752), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n982), .A2(new_n975), .A3(new_n1001), .ZN(new_n1025));
  AND4_X1   g600(.A1(new_n1003), .A2(new_n1022), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1004), .B1(new_n1026), .B2(G301), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1013), .B(new_n1005), .C1(new_n1027), .C2(KEYINPUT54), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1002), .A2(G301), .A3(new_n1003), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1002), .A2(new_n1003), .A3(KEYINPUT121), .A4(G301), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1003), .A2(new_n1022), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(G171), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1028), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT61), .ZN(new_n1039));
  XOR2_X1   g614(.A(G299), .B(KEYINPUT57), .Z(new_n1040));
  INV_X1    g615(.A(new_n977), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n948), .B2(KEYINPUT50), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n703), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT56), .B(G2072), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n949), .A2(new_n919), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1040), .B1(new_n1045), .B2(new_n1043), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1039), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n891), .A2(new_n919), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n997), .A2(new_n698), .B1(new_n766), .B2(new_n1051), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1052), .A2(new_n604), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n604), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT60), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1056));
  XNOR2_X1  g631(.A(G299), .B(KEYINPUT57), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(KEYINPUT61), .A3(new_n1046), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1052), .A2(new_n1060), .A3(new_n593), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1049), .A2(new_n1055), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT58), .B(G1341), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1051), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n890), .A2(G1996), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n975), .B(new_n1066), .C1(new_n955), .C2(KEYINPUT45), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n949), .A2(KEYINPUT115), .A3(new_n1066), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n547), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g648(.A(KEYINPUT116), .B(new_n1065), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1063), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1076));
  XOR2_X1   g651(.A(new_n1076), .B(KEYINPUT118), .Z(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1063), .B(new_n1077), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1062), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1048), .B1(new_n1046), .B2(new_n1054), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT114), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1038), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1018), .A2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(G290), .B(G1986), .Z(new_n1086));
  NAND3_X1  g661(.A1(new_n906), .A2(new_n910), .A3(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1087), .A2(new_n892), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT123), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1091), .B(new_n1088), .C1(new_n1018), .C2(new_n1084), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n916), .B1(new_n1090), .B2(new_n1092), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g668(.A(G227), .ZN(new_n1095));
  NAND2_X1  g669(.A1(G319), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g670(.A(new_n1096), .B1(new_n645), .B2(new_n647), .ZN(new_n1097));
  NAND2_X1  g671(.A1(new_n1097), .A2(new_n681), .ZN(new_n1098));
  XNOR2_X1  g672(.A(new_n1098), .B(KEYINPUT126), .ZN(new_n1099));
  AND3_X1   g673(.A1(new_n1099), .A2(new_n884), .A3(new_n844), .ZN(G308));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n884), .A3(new_n844), .ZN(G225));
endmodule


