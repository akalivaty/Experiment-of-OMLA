//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT71), .B1(new_n194), .B2(G104), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n191), .A3(G107), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT72), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n192), .A2(new_n197), .A3(new_n195), .A4(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT72), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(G101), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT73), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n196), .A2(new_n200), .A3(new_n210), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n211), .A2(new_n206), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n202), .A2(new_n204), .A3(G101), .A4(new_n207), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT2), .B(G113), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G116), .B(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(G116), .B(G119), .Z(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n215), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT5), .ZN(new_n223));
  INV_X1    g037(.A(G119), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G116), .ZN(new_n225));
  OAI211_X1 g039(.A(G113), .B(new_n225), .C1(new_n219), .C2(new_n223), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n218), .ZN(new_n227));
  XOR2_X1   g041(.A(G104), .B(G107), .Z(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G101), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n203), .B2(G101), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT75), .B1(new_n222), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT75), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n227), .A2(new_n230), .ZN(new_n234));
  AOI211_X1 g048(.A(new_n233), .B(new_n234), .C1(new_n214), .C2(new_n221), .ZN(new_n235));
  OAI211_X1 g049(.A(KEYINPUT6), .B(new_n190), .C1(new_n232), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n231), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n233), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n234), .B1(new_n214), .B2(new_n221), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT75), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n189), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n189), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT6), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n236), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G143), .B(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT0), .B(G128), .Z(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G125), .ZN(new_n251));
  INV_X1    g065(.A(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n254), .A3(G143), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n256), .B(G146), .C1(new_n252), .C2(KEYINPUT1), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G125), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n251), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G224), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n251), .A2(new_n266), .A3(new_n263), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n245), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT79), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n267), .A2(KEYINPUT7), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n268), .B2(new_n270), .ZN(new_n277));
  AOI211_X1 g091(.A(KEYINPUT7), .B(new_n267), .C1(new_n251), .C2(new_n263), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n227), .B2(new_n230), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n231), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n189), .B(KEYINPUT8), .ZN(new_n283));
  OR3_X1    g097(.A1(new_n227), .A2(new_n230), .A3(KEYINPUT76), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT77), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n285), .B(KEYINPUT77), .C1(new_n277), .C2(new_n278), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n242), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n275), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT78), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n273), .A2(new_n274), .A3(new_n290), .A4(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n272), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n190), .B1(new_n232), .B2(new_n235), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n243), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n297), .B2(new_n236), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT78), .B(new_n292), .C1(new_n298), .C2(new_n289), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n273), .A2(new_n291), .A3(new_n290), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT79), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n188), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n305), .B1(new_n224), .B2(G128), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n252), .A2(KEYINPUT23), .A3(G119), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n306), .B(new_n307), .C1(G119), .C2(new_n252), .ZN(new_n308));
  XNOR2_X1  g122(.A(G119), .B(G128), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT24), .B(G110), .Z(new_n310));
  AOI22_X1  g124(.A1(new_n308), .A2(G110), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n262), .A2(KEYINPUT16), .A3(G140), .ZN(new_n312));
  XNOR2_X1  g126(.A(G125), .B(G140), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(new_n313), .B2(KEYINPUT16), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G146), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n314), .A2(G146), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT68), .B(G110), .Z(new_n319));
  OAI22_X1  g133(.A1(new_n308), .A2(new_n319), .B1(new_n309), .B2(new_n310), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n254), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(KEYINPUT69), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT69), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n318), .B2(new_n322), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT22), .ZN(new_n328));
  INV_X1    g142(.A(G137), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n324), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n330), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n323), .A2(KEYINPUT69), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n275), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT25), .ZN(new_n335));
  INV_X1    g149(.A(G217), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(G234), .B2(new_n275), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n338), .B(new_n275), .C1(new_n331), .C2(new_n333), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n337), .A2(G902), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n331), .B2(new_n333), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G472), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT11), .ZN(new_n345));
  INV_X1    g159(.A(G134), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(G137), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n329), .A2(KEYINPUT11), .A3(G134), .ZN(new_n348));
  INV_X1    g162(.A(G131), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(G137), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n350), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n346), .A2(G137), .ZN(new_n353));
  OAI21_X1  g167(.A(G131), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n261), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n261), .A2(KEYINPUT65), .A3(new_n351), .A4(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n347), .A2(new_n350), .A3(new_n348), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G131), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n351), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n250), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT64), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT30), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT64), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n366), .A3(new_n250), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n359), .A2(new_n364), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT66), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n362), .A2(new_n369), .A3(new_n250), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n369), .B1(new_n362), .B2(new_n250), .ZN(new_n371));
  INV_X1    g185(.A(new_n355), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n368), .B1(new_n373), .B2(new_n365), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n221), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT31), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n363), .A2(KEYINPUT66), .ZN(new_n377));
  INV_X1    g191(.A(new_n221), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n362), .A2(new_n369), .A3(new_n250), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n355), .ZN(new_n380));
  XOR2_X1   g194(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n381));
  INV_X1    g195(.A(G237), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n265), .A3(G210), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n381), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G101), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n375), .A2(new_n376), .A3(new_n380), .A4(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n359), .A2(new_n367), .A3(new_n364), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n221), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n389), .B1(new_n391), .B2(new_n380), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n363), .A2(new_n378), .A3(new_n355), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n393), .A2(new_n389), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n388), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n387), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n380), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n374), .B2(new_n221), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n376), .B1(new_n398), .B2(new_n386), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n344), .B(new_n275), .C1(new_n396), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT32), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n386), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT31), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n387), .A3(new_n395), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT32), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n344), .A4(new_n275), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n398), .A2(new_n388), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n386), .B1(new_n392), .B2(new_n394), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n377), .A2(new_n379), .A3(new_n355), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n221), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n380), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n394), .B1(new_n413), .B2(KEYINPUT28), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT29), .A3(new_n386), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n275), .ZN(new_n416));
  OAI21_X1  g230(.A(G472), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n343), .B1(new_n407), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n316), .A2(new_n317), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n382), .A2(new_n265), .A3(G214), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(new_n256), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT17), .A3(G131), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(G131), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n420), .B(G143), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n349), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n419), .B(new_n422), .C1(new_n426), .C2(KEYINPUT17), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n424), .B1(new_n428), .B2(new_n349), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n313), .B(new_n254), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n429), .B(new_n430), .C1(new_n428), .C2(new_n423), .ZN(new_n431));
  XOR2_X1   g245(.A(G113), .B(G122), .Z(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT80), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n191), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n427), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n427), .B2(new_n431), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n275), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G475), .ZN(new_n439));
  INV_X1    g253(.A(new_n434), .ZN(new_n440));
  INV_X1    g254(.A(new_n426), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n313), .B(KEYINPUT19), .Z(new_n442));
  OAI21_X1  g256(.A(new_n315), .B1(new_n442), .B2(G146), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n431), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(G475), .B1(new_n445), .B2(new_n435), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n446), .A2(new_n447), .A3(new_n275), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n447), .B1(new_n446), .B2(new_n275), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n439), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G952), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  NAND2_X1  g267(.A1(G234), .A2(G237), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT21), .B(G898), .Z(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT83), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(G902), .A3(G953), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G128), .B(G143), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n346), .B1(new_n461), .B2(KEYINPUT13), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n256), .A2(G128), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(KEYINPUT13), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n346), .ZN(new_n466));
  XNOR2_X1  g280(.A(G116), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n194), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n465), .A2(new_n466), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n461), .B(new_n346), .ZN(new_n471));
  INV_X1    g285(.A(G116), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT14), .A3(G122), .ZN(new_n473));
  INV_X1    g287(.A(new_n467), .ZN(new_n474));
  OAI211_X1 g288(.A(G107), .B(new_n473), .C1(new_n474), .C2(KEYINPUT14), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n471), .B(new_n475), .C1(G107), .C2(new_n474), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT9), .B(G234), .Z(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(G217), .A3(new_n265), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n479), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n470), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n275), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(G478), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(G478), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n483), .A2(new_n484), .A3(new_n275), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n460), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G469), .ZN(new_n492));
  XNOR2_X1  g306(.A(G110), .B(G140), .ZN(new_n493));
  INV_X1    g307(.A(G227), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(G953), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n493), .B(new_n495), .Z(new_n496));
  NAND2_X1  g310(.A1(new_n214), .A2(new_n250), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n211), .A2(new_n261), .A3(new_n229), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT10), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n499), .A2(KEYINPUT10), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n362), .ZN(new_n503));
  INV_X1    g317(.A(new_n362), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n497), .A2(new_n504), .A3(new_n500), .A4(new_n501), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n496), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n261), .B1(new_n211), .B2(new_n229), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT74), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n508), .B2(new_n498), .ZN(new_n509));
  AOI211_X1 g323(.A(KEYINPUT74), .B(new_n261), .C1(new_n211), .C2(new_n229), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n362), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT12), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n513), .B(new_n362), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  AND4_X1   g328(.A1(new_n505), .A2(new_n512), .A3(new_n496), .A4(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n492), .B(new_n275), .C1(new_n506), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(G469), .A2(G902), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n505), .A2(new_n514), .A3(new_n512), .ZN(new_n518));
  INV_X1    g332(.A(new_n496), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n503), .A2(new_n505), .A3(new_n496), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(G469), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n478), .ZN(new_n524));
  OAI21_X1  g338(.A(G221), .B1(new_n524), .B2(G902), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n525), .B(KEYINPUT70), .Z(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n304), .A2(new_n418), .A3(new_n491), .A4(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT84), .B(G101), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(G3));
  OAI21_X1  g346(.A(new_n275), .B1(new_n396), .B2(new_n399), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G472), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n534), .A2(new_n400), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n536), .A2(new_n343), .A3(new_n528), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT85), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n292), .B1(new_n298), .B2(new_n289), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n188), .B1(new_n302), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G478), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT86), .B1(new_n470), .B2(new_n476), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n483), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n542), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n482), .A3(new_n480), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n541), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n483), .A2(new_n541), .A3(new_n275), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n541), .A2(new_n275), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n551), .A2(new_n459), .A3(new_n450), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n540), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n538), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT34), .B(G104), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(G6));
  AND3_X1   g370(.A1(new_n540), .A2(new_n459), .A3(new_n439), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT87), .B1(new_n448), .B2(new_n449), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(KEYINPUT87), .B2(new_n449), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n559), .A2(new_n490), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n538), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT35), .B(G107), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(G9));
  NAND3_X1  g379(.A1(new_n304), .A2(new_n491), .A3(new_n529), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n330), .A2(KEYINPUT36), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n323), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n341), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n340), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n566), .A2(new_n536), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT90), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT37), .B(G110), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G12));
  AOI21_X1  g391(.A(new_n528), .B1(new_n407), .B2(new_n417), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n455), .B(KEYINPUT91), .Z(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(G900), .B2(new_n458), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT92), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n439), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n559), .A2(new_n490), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n578), .A2(new_n540), .A3(new_n572), .A4(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G128), .ZN(G30));
  NAND3_X1  g400(.A1(new_n303), .A2(new_n299), .A3(new_n294), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT93), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT38), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n582), .B(KEYINPUT96), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT39), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n529), .A2(new_n591), .ZN(new_n592));
  AOI211_X1 g406(.A(new_n188), .B(new_n572), .C1(new_n592), .C2(KEYINPUT40), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n411), .A2(KEYINPUT30), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n378), .B1(new_n594), .B2(new_n368), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n386), .B1(new_n595), .B2(new_n397), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n412), .A2(new_n380), .A3(new_n388), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(new_n275), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT94), .B1(new_n599), .B2(G472), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n601), .B(new_n344), .C1(new_n596), .C2(new_n598), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n407), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT95), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n490), .A2(new_n450), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n592), .B2(KEYINPUT40), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n589), .A2(new_n593), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G143), .ZN(G45));
  AND3_X1   g426(.A1(new_n551), .A2(new_n450), .A3(new_n582), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n578), .A2(new_n540), .A3(new_n572), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G146), .ZN(G48));
  OAI21_X1  g429(.A(new_n275), .B1(new_n506), .B2(new_n515), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(G469), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n617), .A2(new_n527), .A3(new_n516), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n418), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n553), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(KEYINPUT97), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n619), .B2(new_n553), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G113), .ZN(G15));
  NAND2_X1  g441(.A1(new_n561), .A2(new_n620), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G116), .ZN(G18));
  NAND2_X1  g443(.A1(new_n302), .A2(new_n539), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n630), .A2(new_n618), .A3(new_n187), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n407), .A2(new_n417), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n491), .A4(new_n572), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G119), .ZN(G21));
  OAI21_X1  g448(.A(new_n387), .B1(new_n386), .B2(new_n414), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n344), .B(new_n275), .C1(new_n635), .C2(new_n399), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n534), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n343), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n188), .B(new_n607), .C1(new_n302), .C2(new_n539), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n459), .A3(new_n618), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G122), .ZN(G24));
  NAND4_X1  g457(.A1(new_n631), .A2(new_n572), .A3(new_n613), .A4(new_n637), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G125), .ZN(G27));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n289), .B1(new_n245), .B2(new_n272), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n274), .B1(new_n647), .B2(new_n291), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n300), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n516), .A2(new_n517), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n520), .A2(new_n521), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT98), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n521), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(G469), .A3(new_n655), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n526), .B(new_n188), .C1(new_n651), .C2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n418), .A2(new_n649), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n613), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n646), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n632), .A2(new_n638), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT99), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n418), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(KEYINPUT42), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n649), .A2(new_n657), .A3(new_n613), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n660), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G131), .ZN(G33));
  NAND4_X1  g482(.A1(new_n418), .A2(new_n649), .A3(new_n657), .A4(new_n584), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT100), .B(G134), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G36));
  NAND2_X1  g485(.A1(new_n649), .A2(new_n187), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n551), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n450), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT43), .Z(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n536), .A3(new_n572), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n673), .B1(new_n679), .B2(KEYINPUT44), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n653), .A2(KEYINPUT45), .A3(new_n655), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n652), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n681), .A2(G469), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n517), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n684), .A2(KEYINPUT46), .A3(new_n517), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n516), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n689), .A2(new_n527), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n591), .B(new_n690), .C1(new_n678), .C2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n680), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT101), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n329), .ZN(G39));
  XOR2_X1   g509(.A(new_n690), .B(KEYINPUT47), .Z(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n659), .A3(new_n672), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n632), .A2(new_n638), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G140), .ZN(G42));
  INV_X1    g514(.A(new_n589), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n526), .A2(new_n188), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n606), .A2(new_n638), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n617), .A2(new_n516), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n706), .A2(KEYINPUT49), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n675), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(KEYINPUT49), .B2(new_n706), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n701), .A2(new_n702), .A3(new_n704), .A4(new_n709), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n187), .B(new_n552), .C1(new_n300), .C2(new_n648), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT102), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n587), .A2(new_n713), .A3(new_n187), .A4(new_n552), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n537), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n530), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n715), .A2(KEYINPUT103), .A3(new_n530), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n574), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n490), .ZN(new_n721));
  AND4_X1   g535(.A1(new_n721), .A2(new_n559), .A3(new_n572), .A4(new_n583), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n649), .A2(new_n578), .A3(new_n722), .A4(new_n187), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n534), .A2(new_n572), .A3(new_n636), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n649), .A2(new_n657), .A3(new_n613), .A4(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n669), .A2(new_n723), .A3(new_n725), .A4(KEYINPUT104), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n669), .A2(new_n723), .A3(new_n725), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n667), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  AND4_X1   g544(.A1(new_n625), .A2(new_n642), .A3(new_n633), .A4(new_n628), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n649), .A2(new_n460), .A3(new_n188), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n490), .A3(new_n537), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n720), .A2(new_n730), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n644), .A2(new_n585), .A3(new_n614), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n340), .A2(new_n527), .A3(new_n571), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n651), .B2(new_n656), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n605), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n630), .A2(new_n187), .A3(new_n582), .A4(new_n608), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT105), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n603), .B1(new_n401), .B2(new_n406), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n340), .A2(new_n527), .A3(new_n571), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n654), .B1(new_n520), .B2(new_n521), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n521), .A2(new_n654), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n492), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n742), .B1(new_n745), .B2(new_n650), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n641), .A4(new_n582), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n740), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT52), .B1(new_n735), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n644), .A2(new_n585), .A3(new_n614), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n740), .A2(new_n749), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT53), .B1(new_n734), .B2(new_n756), .ZN(new_n757));
  OR3_X1    g571(.A1(new_n566), .A2(new_n536), .A3(new_n573), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n715), .A2(KEYINPUT103), .A3(new_n530), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT103), .B1(new_n715), .B2(new_n530), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n758), .B(new_n733), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n625), .A2(new_n642), .A3(new_n633), .A4(new_n628), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n667), .A2(new_n729), .A3(new_n726), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n751), .B2(new_n755), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n735), .A2(new_n750), .A3(KEYINPUT52), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n754), .B1(new_n752), .B2(new_n753), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(KEYINPUT107), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n764), .A2(new_n765), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n757), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n677), .A2(new_n776), .A3(new_n579), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT109), .B1(new_n676), .B2(new_n580), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n639), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n631), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n673), .A2(new_n618), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n703), .A2(new_n781), .A3(new_n455), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n674), .A2(new_n451), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n453), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n777), .A2(new_n778), .ZN(new_n786));
  INV_X1    g600(.A(new_n781), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n662), .A2(new_n664), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n788), .A2(KEYINPUT48), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT48), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n785), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n765), .B1(new_n734), .B2(new_n756), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT106), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(KEYINPUT106), .B(new_n765), .C1(new_n734), .C2(new_n756), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n761), .A2(new_n762), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n771), .A2(new_n797), .A3(KEYINPUT53), .A4(new_n730), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT108), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT108), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n764), .A2(new_n771), .A3(new_n800), .A4(KEYINPUT53), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n795), .A2(new_n796), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n775), .B(new_n792), .C1(new_n802), .C2(new_n774), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n618), .A2(new_n188), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT110), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n701), .A2(new_n779), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT111), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n806), .A2(new_n809), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n810), .A2(KEYINPUT112), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT112), .B1(new_n810), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n696), .B1(new_n527), .B2(new_n706), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n673), .A3(new_n779), .ZN(new_n816));
  INV_X1    g630(.A(new_n788), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n551), .A2(new_n450), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n817), .A2(new_n724), .B1(new_n782), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n810), .A2(new_n811), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n803), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(G952), .A2(G953), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n710), .B1(new_n824), .B2(new_n825), .ZN(G75));
  NOR2_X1   g640(.A1(new_n245), .A2(new_n272), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n298), .ZN(new_n828));
  XOR2_X1   g642(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT114), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n828), .B(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n757), .A2(new_n772), .A3(G210), .A4(G902), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n452), .A2(G953), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT117), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n832), .A2(new_n831), .A3(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n836), .A2(new_n839), .A3(new_n841), .ZN(G51));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n757), .A2(new_n772), .A3(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n775), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n773), .A2(KEYINPUT118), .A3(new_n774), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n517), .B(KEYINPUT57), .Z(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n506), .B2(new_n515), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n773), .A2(new_n275), .A3(new_n684), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n839), .B1(new_n849), .B2(new_n850), .ZN(G54));
  NOR2_X1   g665(.A1(new_n773), .A2(new_n275), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n445), .A2(new_n435), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(KEYINPUT58), .A2(G475), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n852), .A2(KEYINPUT119), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n757), .A2(new_n772), .A3(G902), .A4(new_n855), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n853), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n858), .A2(KEYINPUT120), .A3(new_n853), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT120), .B1(new_n858), .B2(new_n853), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n838), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT121), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n861), .A2(new_n862), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n856), .A2(new_n859), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n838), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n864), .A2(new_n868), .ZN(G60));
  NAND2_X1  g683(.A1(new_n544), .A2(new_n546), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n775), .B1(new_n802), .B2(new_n774), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n550), .B(KEYINPUT59), .Z(new_n873));
  AOI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n871), .A2(new_n845), .A3(new_n846), .A4(new_n873), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n874), .A2(new_n875), .A3(new_n839), .ZN(G63));
  NOR2_X1   g690(.A1(new_n331), .A2(new_n333), .ZN(new_n877));
  XNOR2_X1  g691(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n336), .A2(new_n275), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n877), .B1(new_n773), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n839), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n757), .A2(new_n772), .A3(new_n570), .A4(new_n880), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT61), .A4(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n886), .A2(new_n888), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n882), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n839), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n887), .B1(new_n892), .B2(KEYINPUT61), .ZN(G66));
  AOI21_X1  g707(.A(new_n265), .B1(new_n457), .B2(G224), .ZN(new_n894));
  INV_X1    g708(.A(new_n797), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(new_n265), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n297), .B(new_n236), .C1(G898), .C2(new_n265), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n896), .B(new_n897), .Z(G69));
  XNOR2_X1  g712(.A(new_n442), .B(KEYINPUT125), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n374), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(G900), .A2(G953), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n693), .B1(new_n697), .B2(new_n698), .ZN(new_n902));
  INV_X1    g716(.A(new_n789), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n690), .A2(new_n903), .A3(new_n591), .A4(new_n641), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n667), .A2(new_n669), .A3(new_n735), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n900), .B(new_n901), .C1(new_n906), .C2(G953), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n265), .B1(G227), .B2(G900), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n900), .B(KEYINPUT126), .Z(new_n910));
  NAND2_X1  g724(.A1(new_n611), .A2(new_n735), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT62), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n911), .B(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n912), .A2(KEYINPUT62), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n672), .A2(new_n592), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n721), .A2(new_n450), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n916), .B(new_n418), .C1(new_n783), .C2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n914), .A2(new_n902), .A3(new_n915), .A4(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n910), .B1(new_n919), .B2(new_n265), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n908), .A2(new_n909), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n909), .B1(new_n908), .B2(new_n920), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(G72));
  INV_X1    g737(.A(new_n802), .ZN(new_n924));
  NAND2_X1  g738(.A1(G472), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT63), .Z(new_n926));
  NAND4_X1  g740(.A1(new_n924), .A2(new_n408), .A3(new_n596), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n919), .B2(new_n895), .ZN(new_n928));
  INV_X1    g742(.A(new_n596), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n839), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n926), .B1(new_n906), .B2(new_n895), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n398), .A3(new_n388), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n927), .A2(new_n930), .A3(new_n932), .ZN(G57));
endmodule


