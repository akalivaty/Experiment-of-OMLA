//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NAND2_X1  g0010(.A1(G50), .A2(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  AOI211_X1 g0016(.A(new_n214), .B(new_n216), .C1(G77), .C2(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n207), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n203), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n210), .B(new_n227), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n221), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  INV_X1    g0044(.A(G50), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G58), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT68), .B1(new_n207), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n259), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(new_n228), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n253), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n256), .B1(new_n263), .B2(new_n252), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT7), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n212), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n229), .A2(new_n257), .ZN(new_n274));
  INV_X1    g0074(.A(G159), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT77), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT77), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(G159), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(G58), .B(G68), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT76), .B1(new_n281), .B2(G20), .ZN(new_n282));
  AND2_X1   g0082(.A1(G58), .A2(G68), .ZN(new_n283));
  OAI211_X1 g0083(.A(KEYINPUT76), .B(G20), .C1(new_n283), .C2(new_n203), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n280), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT78), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(G20), .B1(new_n283), .B2(new_n203), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT76), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n284), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(KEYINPUT78), .A3(new_n280), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n273), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n261), .B1(new_n294), .B2(KEYINPUT16), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT16), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(new_n286), .B2(new_n273), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n264), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT67), .ZN(new_n299));
  INV_X1    g0099(.A(G41), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT66), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT66), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G41), .ZN(new_n303));
  AOI21_X1  g0103(.A(G45), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n299), .B1(new_n304), .B2(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G1), .A3(G13), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT66), .B(G41), .ZN(new_n308));
  OAI211_X1 g0108(.A(KEYINPUT67), .B(new_n253), .C1(new_n308), .C2(G45), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n305), .A2(G274), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n307), .A2(G232), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT80), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n307), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G223), .A2(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G1698), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(G226), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n271), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G87), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT79), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n315), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n310), .A2(new_n314), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G200), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n298), .A2(KEYINPUT17), .A3(new_n324), .A4(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n273), .ZN(new_n328));
  AOI221_X4 g0128(.A(new_n287), .B1(new_n276), .B2(new_n279), .C1(new_n291), .C2(new_n284), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT78), .B1(new_n292), .B2(new_n280), .ZN(new_n330));
  OAI211_X1 g0130(.A(KEYINPUT16), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n258), .A2(new_n228), .A3(new_n260), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n332), .A3(new_n297), .ZN(new_n333));
  INV_X1    g0133(.A(new_n264), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n333), .A2(new_n324), .A3(new_n326), .A4(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n323), .A2(G169), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n310), .A2(new_n314), .A3(new_n322), .A4(G179), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT18), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT18), .ZN(new_n343));
  AOI221_X4 g0143(.A(new_n343), .B1(new_n339), .B2(new_n340), .C1(new_n333), .C2(new_n334), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n327), .B(new_n337), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT81), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n335), .B(KEYINPUT17), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n338), .A2(new_n341), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n343), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n338), .A2(new_n341), .A3(KEYINPUT18), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(new_n352), .A3(KEYINPUT81), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n307), .A2(G238), .A3(new_n311), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n236), .A2(G1698), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(G226), .B2(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n357), .B2(new_n271), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n354), .B1(new_n358), .B2(new_n315), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n310), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT13), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n310), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(KEYINPUT74), .A3(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n363), .A2(KEYINPUT74), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(KEYINPUT75), .B2(KEYINPUT14), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n361), .A2(new_n363), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G179), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n364), .A2(new_n365), .A3(new_n367), .A4(new_n369), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n254), .B(KEYINPUT69), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n376), .A2(new_n261), .A3(new_n262), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT12), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n212), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n212), .A2(G20), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n229), .A2(G33), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n381), .B1(new_n382), .B2(new_n202), .C1(new_n245), .C2(new_n274), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n332), .ZN(new_n384));
  XOR2_X1   g0184(.A(new_n384), .B(KEYINPUT11), .Z(new_n385));
  NOR3_X1   g0185(.A1(new_n376), .A2(new_n378), .A3(G68), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n255), .A2(KEYINPUT12), .ZN(new_n387));
  NOR4_X1   g0187(.A1(new_n380), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n375), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n307), .A2(G226), .A3(new_n311), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n317), .A2(G222), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G223), .A2(G1698), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n266), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n315), .C1(G77), .C2(new_n266), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n310), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n396), .A2(G179), .ZN(new_n397));
  INV_X1    g0197(.A(G150), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n252), .A2(new_n382), .B1(new_n398), .B2(new_n274), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n229), .B1(new_n201), .B2(new_n203), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n332), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n255), .A2(new_n245), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n401), .B(new_n402), .C1(new_n245), .C2(new_n263), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n396), .A2(new_n366), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n347), .A2(new_n353), .A3(new_n390), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT9), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT71), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n396), .A2(G200), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(KEYINPUT73), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n412), .A2(KEYINPUT10), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n396), .A2(new_n325), .ZN(new_n415));
  OR3_X1    g0215(.A1(new_n403), .A2(KEYINPUT72), .A3(new_n407), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT72), .B1(new_n403), .B2(new_n407), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n411), .A2(new_n414), .A3(new_n415), .A4(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n409), .A2(new_n410), .A3(new_n418), .A4(new_n415), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n413), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n406), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n372), .A2(G190), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n364), .A2(G200), .A3(new_n365), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n388), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n377), .A2(G77), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT69), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n254), .B(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n202), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT15), .B(G87), .Z(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n382), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n252), .A2(new_n274), .B1(new_n229), .B2(new_n202), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n332), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n427), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G238), .A2(G1698), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n266), .B(new_n438), .C1(new_n236), .C2(G1698), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(new_n315), .C1(G107), .C2(new_n266), .ZN(new_n440));
  INV_X1    g0240(.A(G179), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n307), .A2(G244), .A3(new_n311), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n310), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT70), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n444), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n437), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n310), .A2(new_n442), .A3(new_n440), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n366), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n448), .A2(new_n325), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(G200), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n437), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n426), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n268), .A2(new_n270), .A3(G244), .A4(new_n317), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT4), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT4), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n266), .A2(new_n458), .A3(G244), .A4(new_n317), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT82), .ZN(new_n462));
  AND4_X1   g0262(.A1(G250), .A2(new_n268), .A3(new_n270), .A4(G1698), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n460), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n315), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n301), .A2(new_n303), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n300), .A2(KEYINPUT5), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n468), .A2(G274), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G257), .A3(new_n307), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n466), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G200), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n254), .A2(G97), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n254), .B1(G1), .B2(new_n257), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n332), .A2(new_n223), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT7), .B1(new_n271), .B2(new_n229), .ZN(new_n480));
  AOI211_X1 g0280(.A(new_n265), .B(G20), .C1(new_n268), .C2(new_n270), .ZN(new_n481));
  OAI21_X1  g0281(.A(G107), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  INV_X1    g0283(.A(G107), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n223), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(KEYINPUT6), .A3(G97), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n229), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n277), .A2(G77), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n482), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI211_X1 g0292(.A(new_n477), .B(new_n479), .C1(new_n492), .C2(new_n332), .ZN(new_n493));
  INV_X1    g0293(.A(new_n472), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n465), .B2(new_n315), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G190), .A3(new_n474), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n476), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n219), .B1(new_n470), .B2(G1), .ZN(new_n498));
  INV_X1    g0298(.A(G274), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n253), .A2(new_n499), .A3(G45), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n307), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n213), .A2(new_n317), .ZN(new_n502));
  INV_X1    g0302(.A(G244), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G1698), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n268), .A2(new_n502), .A3(new_n270), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G116), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n501), .B1(new_n507), .B2(new_n315), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT83), .B1(new_n508), .B2(new_n441), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n307), .A2(new_n498), .A3(new_n500), .ZN(new_n510));
  INV_X1    g0310(.A(new_n506), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G238), .A2(G1698), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n503), .B2(G1698), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n513), .B2(new_n266), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n441), .B(new_n510), .C1(new_n514), .C2(new_n307), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n508), .B2(G169), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n509), .B1(new_n516), .B2(KEYINPUT83), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n268), .A2(new_n270), .A3(new_n229), .A4(G68), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT84), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n266), .A2(KEYINPUT84), .A3(new_n229), .A4(G68), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT19), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n229), .B1(new_n355), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n486), .A2(new_n218), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n229), .A2(G33), .A3(G97), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n523), .A2(new_n524), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n332), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n429), .A2(new_n432), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n332), .A2(new_n478), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n431), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n307), .B1(new_n505), .B2(new_n506), .ZN(new_n533));
  OAI21_X1  g0333(.A(G200), .B1(new_n533), .B2(new_n501), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(G87), .ZN(new_n535));
  AND4_X1   g0335(.A1(new_n529), .A2(new_n528), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT85), .B1(new_n508), .B2(G190), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT85), .ZN(new_n538));
  NOR4_X1   g0338(.A1(new_n533), .A2(new_n538), .A3(new_n501), .A4(new_n325), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n517), .A2(new_n532), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n477), .ZN(new_n542));
  INV_X1    g0342(.A(new_n479), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n484), .B1(new_n267), .B2(new_n272), .ZN(new_n544));
  INV_X1    g0344(.A(new_n491), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n544), .A2(new_n545), .A3(new_n489), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n542), .B(new_n543), .C1(new_n546), .C2(new_n261), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n466), .A2(new_n441), .A3(new_n472), .A4(new_n474), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n463), .B1(new_n457), .B2(new_n459), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n307), .B1(new_n549), .B2(new_n462), .ZN(new_n550));
  INV_X1    g0350(.A(new_n474), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n550), .A2(new_n494), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n547), .B(new_n548), .C1(new_n552), .C2(G169), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT24), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n268), .A2(new_n270), .A3(new_n229), .A4(G87), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT22), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n266), .A2(KEYINPUT22), .A3(new_n229), .A4(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT23), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(new_n484), .A3(G20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT87), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT87), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n560), .A3(new_n484), .A4(G20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n506), .A2(new_n560), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(new_n229), .B1(KEYINPUT23), .B2(G107), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n554), .B1(new_n559), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n570), .A2(G20), .B1(new_n560), .B2(new_n484), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n562), .B2(new_n564), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n572), .A2(KEYINPUT24), .A3(new_n557), .A4(new_n558), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n569), .A2(new_n332), .A3(new_n573), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n332), .A2(new_n484), .A3(new_n478), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT88), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT25), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n576), .B(new_n577), .C1(new_n255), .C2(new_n484), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  NOR2_X1   g0379(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n580));
  NOR4_X1   g0380(.A1(new_n579), .A2(new_n254), .A3(G107), .A4(new_n580), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n575), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n473), .A2(G264), .A3(new_n307), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n219), .A2(new_n317), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n224), .A2(G1698), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n268), .A2(new_n585), .A3(new_n270), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G294), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n315), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n584), .A2(new_n590), .A3(new_n472), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n366), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n591), .A2(G179), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n583), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n497), .A2(new_n541), .A3(new_n553), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(G200), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n584), .A2(new_n590), .A3(G190), .A4(new_n472), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n574), .A2(new_n596), .A3(new_n597), .A4(new_n582), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT89), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT20), .ZN(new_n601));
  AOI21_X1  g0401(.A(G20), .B1(new_n257), .B2(G97), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n462), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n220), .A2(G20), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n332), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n601), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n462), .A2(new_n602), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n607), .A2(KEYINPUT20), .A3(new_n332), .A4(new_n604), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n220), .B1(new_n253), .B2(G33), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n376), .A2(new_n261), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n429), .A2(new_n220), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n473), .A2(G270), .A3(new_n307), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n317), .A2(G257), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G264), .A2(G1698), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n266), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g0419(.A(KEYINPUT86), .B(G303), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n271), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n621), .A3(new_n315), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n616), .A2(new_n472), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n615), .A2(new_n623), .A3(KEYINPUT21), .A4(G169), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT21), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n613), .B1(new_n606), .B2(new_n608), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(G169), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n623), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n615), .A2(G179), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(G190), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n623), .A2(G200), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n624), .A2(new_n628), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n595), .A2(new_n600), .A3(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n423), .A2(new_n455), .A3(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n405), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n419), .A2(KEYINPUT90), .A3(new_n421), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT90), .B1(new_n419), .B2(new_n421), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n450), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n389), .A2(new_n375), .B1(new_n641), .B2(new_n426), .ZN(new_n642));
  INV_X1    g0442(.A(new_n348), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n352), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n637), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n423), .A2(new_n455), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n536), .A2(new_n540), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n574), .A2(new_n582), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n650), .A2(new_n599), .A3(new_n597), .A4(new_n596), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n598), .A2(KEYINPUT89), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n594), .A2(new_n624), .A3(new_n628), .A4(new_n630), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n497), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n649), .B1(new_n655), .B2(new_n553), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n528), .A2(new_n529), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n516), .B1(new_n657), .B2(new_n531), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n541), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n553), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n661), .B2(new_n648), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n645), .B1(new_n646), .B2(new_n663), .ZN(G369));
  NAND3_X1  g0464(.A1(new_n624), .A2(new_n628), .A3(new_n630), .ZN(new_n665));
  INV_X1    g0465(.A(G13), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G20), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n253), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n626), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n665), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n634), .B2(new_n675), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n594), .A2(new_n673), .ZN(new_n678));
  INV_X1    g0478(.A(new_n652), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n598), .A2(KEYINPUT89), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n679), .A2(new_n680), .B1(new_n650), .B2(new_n674), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n681), .B2(new_n594), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n665), .A2(new_n674), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI211_X1 g0484(.A(G330), .B(new_n677), .C1(new_n682), .C2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n678), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n650), .A2(new_n674), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n651), .B2(new_n652), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(new_n665), .A3(new_n594), .A4(new_n674), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n686), .A3(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n208), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n308), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n524), .A2(G116), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G1), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n232), .B2(new_n693), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n698), .B(new_n674), .C1(new_n656), .C2(new_n662), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n653), .A2(new_n654), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n497), .A2(new_n647), .A3(new_n553), .A4(new_n659), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n659), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n553), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(KEYINPUT26), .A3(new_n647), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n661), .B2(KEYINPUT26), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n673), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n699), .B1(new_n707), .B2(new_n698), .ZN(new_n708));
  INV_X1    g0508(.A(G330), .ZN(new_n709));
  NOR4_X1   g0509(.A1(new_n595), .A2(new_n600), .A3(new_n634), .A4(new_n673), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n510), .B1(new_n514), .B2(new_n307), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT92), .ZN(new_n713));
  AND4_X1   g0513(.A1(new_n441), .A2(new_n475), .A3(new_n623), .A4(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT91), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n584), .A2(new_n590), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n712), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n495), .A3(new_n474), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n508), .A2(KEYINPUT91), .A3(new_n590), .A4(new_n584), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n629), .A2(new_n719), .A3(G179), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT30), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n616), .A2(G179), .A3(new_n622), .A4(new_n472), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n716), .A2(new_n712), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(KEYINPUT91), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(new_n725), .A3(new_n552), .A4(new_n717), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n591), .A2(new_n714), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT93), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n673), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n721), .A2(new_n726), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n552), .A2(new_n629), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n441), .A3(new_n591), .A4(new_n713), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n730), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n710), .A2(new_n711), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n727), .A2(new_n711), .A3(new_n674), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n709), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n708), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n697), .B1(new_n738), .B2(G1), .ZN(G364));
  OAI21_X1  g0539(.A(G20), .B1(KEYINPUT96), .B2(G169), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(KEYINPUT96), .A2(G169), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n228), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n325), .A2(G179), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n229), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n229), .A2(new_n441), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G294), .A2(new_n746), .B1(new_n750), .B2(G326), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT98), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G190), .A2(G200), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n747), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n752), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n229), .A2(G179), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(new_n325), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(G283), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(G303), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n758), .A2(new_n754), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n266), .B1(new_n766), .B2(G329), .ZN(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n747), .A2(G190), .A3(new_n749), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n747), .A2(new_n325), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT97), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n747), .A2(KEYINPUT97), .A3(new_n325), .A4(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT99), .B(G317), .Z(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT33), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n767), .B1(new_n768), .B2(new_n769), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  NOR4_X1   g0578(.A1(new_n757), .A2(new_n761), .A3(new_n764), .A4(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n774), .A2(G68), .B1(G97), .B2(new_n746), .ZN(new_n780));
  INV_X1    g0580(.A(G58), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(new_n769), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n759), .A2(new_n484), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G77), .B2(new_n755), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n271), .B1(new_n750), .B2(G50), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(new_n218), .C2(new_n762), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n766), .A2(G159), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT32), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n782), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n743), .B1(new_n779), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n266), .A2(G355), .A3(new_n208), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n247), .A2(new_n470), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n691), .A2(new_n266), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n232), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n791), .B1(G116), .B2(new_n208), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n743), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n798), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n790), .B(new_n800), .C1(new_n677), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n667), .A2(G45), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT95), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(KEYINPUT95), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(G1), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n692), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT94), .B1(new_n677), .B2(G330), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n677), .A2(G330), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n809), .B(new_n810), .Z(new_n811));
  OAI21_X1  g0611(.A(new_n808), .B1(new_n811), .B2(new_n807), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT100), .Z(G396));
  NAND2_X1  g0613(.A1(new_n450), .A2(KEYINPUT101), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT101), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n447), .A2(new_n815), .A3(new_n449), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n453), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n436), .A2(new_n673), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n817), .A2(new_n818), .B1(new_n641), .B2(new_n673), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n663), .B2(new_n673), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n674), .B(new_n817), .C1(new_n656), .C2(new_n662), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n600), .A2(new_n634), .ZN(new_n823));
  INV_X1    g0623(.A(new_n595), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n823), .A2(new_n824), .A3(new_n674), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n728), .B1(new_n730), .B2(new_n732), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n674), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n727), .A2(new_n728), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n825), .A2(KEYINPUT31), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(G330), .B1(new_n829), .B2(new_n735), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n822), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n807), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n737), .A2(new_n820), .A3(new_n821), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n819), .A2(new_n796), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n743), .A2(new_n796), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n202), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n775), .A2(new_n760), .B1(new_n223), .B2(new_n745), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n765), .A2(new_n753), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n759), .A2(new_n218), .ZN(new_n840));
  INV_X1    g0640(.A(G294), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n271), .B1(new_n762), .B2(new_n484), .C1(new_n841), .C2(new_n769), .ZN(new_n842));
  NOR4_X1   g0642(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n750), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n220), .B2(new_n756), .C1(new_n763), .C2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n769), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G137), .A2(new_n750), .B1(new_n846), .B2(G143), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n847), .B1(new_n275), .B2(new_n756), .C1(new_n775), .C2(new_n398), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT34), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n849), .B1(new_n245), .B2(new_n762), .C1(new_n212), .C2(new_n759), .ZN(new_n850));
  INV_X1    g0650(.A(G132), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n266), .B1(new_n765), .B2(new_n851), .C1(new_n745), .C2(new_n781), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n845), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n743), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n835), .A2(new_n807), .A3(new_n837), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n834), .A2(new_n855), .ZN(G384));
  INV_X1    g0656(.A(new_n826), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n857), .A2(new_n828), .A3(KEYINPUT31), .A4(new_n673), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n711), .B1(new_n635), .B2(new_n674), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n733), .A2(new_n826), .A3(new_n674), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n423), .A2(new_n455), .A3(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT106), .Z(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  INV_X1    g0664(.A(new_n671), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n331), .A2(new_n332), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n294), .A2(KEYINPUT16), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n334), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n345), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n339), .A2(new_n340), .A3(new_n671), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n338), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n872), .A3(new_n335), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n868), .A2(new_n870), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n874), .A2(new_n335), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n875), .B2(new_n872), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n869), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n389), .A2(new_n673), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n880), .A2(new_n426), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT105), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n375), .A2(new_n882), .A3(new_n389), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n375), .B2(new_n389), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n375), .A2(new_n389), .A3(new_n673), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n819), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n861), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n864), .B1(new_n879), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n345), .A2(new_n338), .A3(new_n865), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n871), .A2(new_n335), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n873), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n876), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n819), .B1(new_n734), .B2(new_n858), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n900), .A4(new_n887), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n890), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n863), .B(new_n902), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(G330), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT38), .B1(new_n891), .B2(new_n894), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n877), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n869), .A2(new_n876), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n896), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n883), .A2(new_n884), .A3(new_n673), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n907), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n352), .A2(new_n865), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n898), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n814), .A2(new_n674), .A3(new_n816), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n821), .A2(new_n915), .B1(new_n885), .B2(new_n886), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n708), .A2(new_n423), .A3(new_n455), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n645), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  XNOR2_X1  g0721(.A(new_n904), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n253), .B2(new_n667), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n232), .A2(new_n202), .A3(new_n283), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT103), .Z(new_n925));
  INV_X1    g0725(.A(new_n201), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n212), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(G1), .A3(new_n666), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT104), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n487), .A2(new_n488), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n220), .B1(new_n930), .B2(KEYINPUT35), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(new_n230), .C1(KEYINPUT35), .C2(new_n930), .ZN(new_n932));
  XOR2_X1   g0732(.A(KEYINPUT102), .B(KEYINPUT36), .Z(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n923), .A2(new_n929), .A3(new_n934), .ZN(G367));
  NAND2_X1  g0735(.A1(new_n704), .A2(new_n673), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n547), .A2(new_n673), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n497), .A2(new_n553), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(KEYINPUT107), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT107), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n936), .B2(new_n938), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n940), .A2(new_n594), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n674), .B1(new_n943), .B2(new_n704), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n689), .A2(new_n938), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT42), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n657), .A2(new_n535), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n673), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n659), .A2(new_n647), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n659), .B2(new_n948), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n944), .A2(new_n946), .A3(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(KEYINPUT108), .B(KEYINPUT109), .Z(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n944), .A2(new_n946), .A3(new_n951), .A4(new_n953), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n950), .B(KEYINPUT43), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n944), .A2(new_n946), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n955), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n940), .A2(new_n942), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(new_n685), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n959), .B(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n806), .ZN(new_n964));
  INV_X1    g0764(.A(new_n738), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n677), .A2(G330), .ZN(new_n967));
  INV_X1    g0767(.A(new_n594), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n686), .B1(new_n688), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n967), .A2(new_n969), .A3(new_n683), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n685), .A2(new_n970), .A3(new_n689), .ZN(new_n971));
  INV_X1    g0771(.A(new_n706), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n674), .B1(new_n972), .B2(new_n702), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT29), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n830), .A2(new_n971), .A3(new_n974), .A4(new_n699), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n689), .A2(new_n686), .ZN(new_n977));
  INV_X1    g0777(.A(new_n939), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(KEYINPUT44), .B(new_n939), .C1(new_n689), .C2(new_n686), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n977), .B2(new_n978), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n689), .A2(KEYINPUT45), .A3(new_n686), .A4(new_n939), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n966), .B1(new_n975), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n981), .A2(new_n985), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n738), .A2(KEYINPUT110), .A3(new_n971), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n965), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n692), .B(KEYINPUT41), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n964), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n963), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n793), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n799), .B1(new_n208), .B2(new_n432), .C1(new_n242), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n759), .A2(new_n223), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n844), .A2(new_n753), .B1(new_n620), .B2(new_n769), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(G107), .C2(new_n746), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n774), .A2(G294), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n762), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(G116), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT46), .ZN(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n271), .B1(new_n765), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G283), .B2(new_n755), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .A4(new_n1006), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n750), .A2(G143), .ZN(new_n1008));
  INV_X1    g0808(.A(G137), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n762), .A2(new_n781), .B1(new_n765), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT111), .Z(new_n1011));
  INV_X1    g0811(.A(new_n759), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n271), .B1(new_n1012), .B2(G77), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n755), .A2(new_n926), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n745), .A2(new_n212), .B1(new_n769), .B2(new_n398), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G159), .B2(new_n774), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1007), .B1(new_n1008), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT47), .Z(new_n1019));
  INV_X1    g0819(.A(new_n743), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n807), .B(new_n996), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n950), .A2(new_n801), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n994), .A2(new_n1024), .ZN(G387));
  NAND2_X1  g0825(.A1(new_n239), .A2(G45), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT113), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n252), .A2(G50), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n694), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1027), .A2(new_n793), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n266), .A2(new_n208), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(G107), .B2(new_n208), .C1(new_n694), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1034), .A2(new_n799), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n969), .A2(new_n798), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n807), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n750), .A2(G159), .B1(G150), .B2(new_n766), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n202), .B2(new_n762), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n997), .B(new_n1039), .C1(G68), .C2(new_n755), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n252), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n774), .A2(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n432), .A2(new_n745), .B1(new_n245), .B2(new_n769), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT114), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n266), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n620), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n774), .A2(G311), .B1(new_n1046), .B2(new_n755), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n1004), .B2(new_n769), .C1(new_n768), .C2(new_n844), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT48), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n760), .B2(new_n745), .C1(new_n841), .C2(new_n762), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT49), .Z(new_n1051));
  AOI21_X1  g0851(.A(new_n266), .B1(new_n766), .B2(G326), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n220), .B2(new_n759), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1045), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1035), .B(new_n1037), .C1(new_n1054), .C2(new_n743), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n975), .A2(new_n692), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT115), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n971), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1056), .A2(KEYINPUT115), .B1(new_n965), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1055), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n971), .A2(new_n806), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT112), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(G393));
  INV_X1    g0863(.A(new_n685), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n988), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n981), .A2(new_n685), .A3(new_n985), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1065), .A2(new_n1066), .B1(new_n738), .B2(new_n971), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT118), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1067), .A2(new_n1068), .B1(new_n987), .B2(new_n989), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT119), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1066), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n685), .B1(new_n981), .B2(new_n985), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n975), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n693), .B1(new_n1073), .B2(KEYINPUT118), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n1069), .A2(new_n1070), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1070), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1065), .A2(KEYINPUT116), .A3(new_n1066), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n806), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n832), .B1(new_n961), .B2(new_n798), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n799), .B1(new_n223), .B2(new_n208), .C1(new_n250), .C2(new_n995), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n745), .A2(new_n202), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n844), .A2(new_n398), .B1(new_n275), .B2(new_n769), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT51), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n271), .B(new_n840), .C1(new_n774), .C2(new_n926), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1001), .A2(G68), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1041), .A2(new_n755), .B1(new_n766), .B2(G143), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n844), .A2(new_n1004), .B1(new_n753), .B2(new_n769), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n266), .B(new_n783), .C1(new_n774), .C2(new_n1046), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n746), .A2(G116), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G294), .A2(new_n755), .B1(new_n766), .B2(G322), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n762), .A2(new_n760), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1083), .A2(new_n1089), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n743), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1081), .A2(new_n1082), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT117), .B1(new_n1080), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1080), .A2(KEYINPUT117), .A3(new_n1099), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1075), .A2(new_n1076), .B1(new_n1100), .B2(new_n1101), .ZN(G390));
  INV_X1    g0902(.A(KEYINPUT120), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n821), .A2(new_n915), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n887), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n911), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n907), .A2(new_n910), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n737), .A2(new_n888), .A3(new_n887), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1106), .B1(new_n877), .B2(new_n906), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n674), .B(new_n817), .C1(new_n972), .C2(new_n702), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1110), .A2(new_n915), .B1(new_n885), .B2(new_n886), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  OR3_X1    g0912(.A1(new_n1107), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n887), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n861), .A2(G330), .A3(new_n888), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1107), .A2(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n423), .A2(G330), .A3(new_n455), .A4(new_n861), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n919), .A3(new_n645), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1115), .A2(new_n1114), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n887), .B1(new_n737), .B2(new_n888), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1104), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1115), .A2(new_n1114), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1123), .A2(new_n915), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1119), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1103), .B1(new_n1117), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n907), .A2(new_n910), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1112), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1120), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1107), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1125), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1119), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1136), .A2(new_n1113), .A3(KEYINPUT120), .A4(new_n1116), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1126), .A2(new_n692), .A3(new_n1133), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n836), .A2(new_n252), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n762), .A2(new_n398), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G159), .A2(new_n746), .B1(new_n846), .B2(G132), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n1009), .C2(new_n775), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n266), .B1(new_n759), .B2(new_n201), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT121), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1144), .A2(new_n1145), .B1(new_n750), .B2(G128), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1145), .B2(new_n1144), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT54), .B(G143), .Z(new_n1149));
  NAND2_X1  g0949(.A1(new_n755), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n766), .A2(G125), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n844), .A2(new_n760), .B1(new_n762), .B2(new_n218), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n756), .A2(new_n223), .B1(new_n212), .B2(new_n759), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n266), .B(new_n1083), .C1(G116), .C2(new_n846), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n766), .A2(G294), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n774), .A2(G107), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1020), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n832), .B(new_n1160), .C1(new_n1127), .C2(new_n796), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1117), .A2(new_n806), .B1(new_n1139), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1138), .A2(new_n1162), .ZN(G378));
  NAND3_X1  g0963(.A1(new_n890), .A2(new_n901), .A3(G330), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n403), .A2(new_n865), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n640), .B2(new_n405), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n638), .A2(new_n639), .A3(new_n637), .A4(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT123), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n912), .A2(new_n1171), .A3(new_n917), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n912), .B2(new_n917), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1164), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1171), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n918), .A2(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n890), .A2(G330), .A3(new_n901), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n912), .A2(new_n1171), .A3(new_n917), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1174), .A2(new_n1179), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n308), .B(new_n266), .C1(new_n1001), .C2(G77), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT122), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n759), .A2(new_n781), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n774), .B2(G97), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G68), .A2(new_n746), .B1(new_n750), .B2(G116), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n431), .B2(new_n755), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n484), .B2(new_n769), .C1(new_n760), .C2(new_n765), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT58), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n245), .B1(G33), .B2(G41), .C1(new_n308), .C2(new_n266), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n774), .A2(G132), .B1(G137), .B2(new_n755), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n750), .A2(G125), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n846), .A2(G128), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n746), .A2(G150), .B1(new_n1001), .B2(new_n1149), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT59), .Z(new_n1197));
  INV_X1    g0997(.A(G124), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n759), .A2(new_n275), .B1(new_n765), .B2(new_n1198), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1199), .A2(G33), .A3(G41), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1191), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1020), .B1(new_n1189), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1168), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1170), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n797), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1202), .B(new_n1205), .C1(new_n201), .C2(new_n836), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1180), .A2(new_n806), .B1(new_n807), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(KEYINPUT57), .A3(new_n1180), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n692), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1133), .A2(new_n1135), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(KEYINPUT57), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1207), .B1(new_n1210), .B2(new_n1212), .ZN(G375));
  AOI22_X1  g1013(.A1(new_n774), .A2(G116), .B1(G77), .B2(new_n1012), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n431), .A2(new_n746), .B1(new_n846), .B2(G283), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n763), .C2(new_n765), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n756), .A2(new_n484), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n762), .A2(new_n223), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n271), .B1(new_n844), .B2(new_n841), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n762), .A2(new_n275), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1183), .B(new_n1221), .C1(G128), .C2(new_n766), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n846), .A2(G137), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n774), .A2(new_n1149), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n266), .B1(new_n745), .B2(new_n245), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G132), .B2(new_n750), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G150), .B2(new_n755), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n743), .B1(new_n1220), .B2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n807), .B(new_n1229), .C1(new_n887), .C2(new_n797), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n212), .B2(new_n836), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1134), .B2(new_n806), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1122), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n991), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(new_n1125), .ZN(G381));
  NAND2_X1  g1035(.A1(new_n1069), .A2(new_n1074), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT119), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1069), .A2(new_n1070), .A3(new_n1074), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(G393), .A2(G396), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1023), .B1(new_n963), .B2(new_n993), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1100), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1080), .A2(KEYINPUT117), .A3(new_n1099), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1245), .A2(G384), .A3(G381), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1138), .A2(new_n1162), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1180), .A2(new_n806), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1206), .A2(new_n807), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n693), .B1(new_n1211), .B2(KEYINPUT57), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1208), .A2(new_n1180), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT57), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1250), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1246), .A2(new_n1247), .A3(new_n1255), .ZN(G407));
  NOR2_X1   g1056(.A1(new_n1246), .A2(new_n672), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1247), .ZN(new_n1258));
  OAI21_X1  g1058(.A(G213), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT124), .Z(G409));
  NAND2_X1  g1060(.A1(new_n672), .A2(G213), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1211), .A2(new_n991), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1138), .A2(new_n1262), .A3(new_n1162), .A4(new_n1207), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1261), .B(new_n1263), .C1(new_n1255), .C2(new_n1247), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1261), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1233), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1122), .A2(new_n1119), .A3(new_n1124), .A4(KEYINPUT60), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n1136), .A3(new_n692), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1232), .ZN(new_n1270));
  INV_X1    g1070(.A(G384), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(G384), .A3(new_n1232), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G2897), .B(new_n1265), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1265), .A2(G2897), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1272), .A2(KEYINPUT125), .A3(new_n1273), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT125), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1264), .A2(new_n1276), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G375), .A2(G378), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1274), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1282), .A2(new_n1283), .A3(new_n1261), .A4(new_n1263), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT63), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G390), .A2(G387), .ZN(new_n1288));
  INV_X1    g1088(.A(G396), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1240), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1239), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1288), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1287), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT126), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1297), .B(new_n1287), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1296), .A2(new_n1298), .B1(new_n1299), .B2(new_n1284), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1286), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT62), .B1(new_n1264), .B2(new_n1274), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1265), .B1(G375), .B2(G378), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1283), .A4(new_n1263), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1302), .A2(new_n1305), .A3(new_n1281), .A4(new_n1287), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1301), .A2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(new_n1282), .A2(new_n1258), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT127), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1311), .A3(new_n1283), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1282), .B(new_n1258), .C1(KEYINPUT127), .C2(new_n1274), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1307), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1314), .B(new_n1315), .ZN(G402));
endmodule


