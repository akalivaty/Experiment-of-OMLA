//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT66), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n209), .A2(new_n210), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT65), .ZN(new_n218));
  INV_X1    g0018(.A(new_n206), .ZN(new_n219));
  INV_X1    g0019(.A(G13), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR3_X1   g0021(.A1(new_n206), .A2(KEYINPUT65), .A3(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n217), .B(new_n226), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT69), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G41), .A2(G45), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n250), .B1(new_n251), .B2(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n255), .B(KEYINPUT69), .C1(G41), .C2(G45), .ZN(new_n256));
  AND3_X1   g0056(.A1(new_n252), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G226), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n254), .A3(G274), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT71), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n253), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n265), .A2(new_n264), .A3(new_n253), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(G223), .A3(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G77), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n270), .B(new_n271), .C1(new_n272), .C2(new_n268), .ZN(new_n273));
  AOI211_X1 g0073(.A(new_n266), .B(new_n267), .C1(new_n273), .C2(KEYINPUT70), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n263), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G50), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n227), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n255), .B2(G20), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n280), .B1(new_n283), .B2(G50), .ZN(new_n284));
  OAI21_X1  g0084(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT72), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G58), .ZN(new_n293));
  OR3_X1    g0093(.A1(new_n291), .A2(new_n293), .A3(KEYINPUT8), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n228), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n289), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n282), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n284), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n276), .B2(G169), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n278), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n276), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n301), .B(KEYINPUT9), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n276), .A2(G190), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n279), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT12), .B1(new_n314), .B2(KEYINPUT76), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(KEYINPUT76), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G50), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n288), .A2(new_n318), .B1(new_n228), .B2(G68), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n297), .A2(new_n272), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n282), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT11), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n321), .A2(new_n322), .B1(G68), .B2(new_n283), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n317), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n268), .A2(G226), .A3(new_n269), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G97), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n267), .A2(new_n266), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n262), .B(KEYINPUT75), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n257), .A2(G238), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n331), .A2(new_n332), .A3(new_n336), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(G169), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n335), .A2(G179), .A3(new_n337), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n339), .B1(new_n338), .B2(G169), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n325), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n325), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n338), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n304), .B1(new_n335), .B2(new_n337), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n295), .A2(new_n283), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n295), .B2(new_n279), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n268), .A2(new_n354), .A3(G20), .ZN(new_n355));
  INV_X1    g0155(.A(G33), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G33), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT7), .B1(new_n360), .B2(new_n228), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n293), .A2(new_n313), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n363), .B2(new_n201), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n287), .A2(G159), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n300), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n362), .A2(KEYINPUT16), .A3(new_n367), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n353), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n252), .A2(G232), .A3(new_n254), .A4(new_n256), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n262), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n357), .A2(new_n359), .A3(G226), .A4(G1698), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT77), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n268), .A2(KEYINPUT77), .A3(G226), .A4(G1698), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n268), .A2(G223), .A3(new_n269), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n374), .B1(new_n381), .B2(new_n330), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n277), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G169), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT18), .B1(new_n372), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n354), .B1(new_n268), .B2(G20), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n360), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n313), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n369), .B1(new_n388), .B2(new_n366), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n371), .A2(new_n389), .A3(new_n282), .ZN(new_n390));
  INV_X1    g0190(.A(new_n353), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n382), .A2(G169), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n383), .A4(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n385), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n382), .A2(G200), .ZN(new_n397));
  AOI211_X1 g0197(.A(G190), .B(new_n374), .C1(new_n381), .C2(new_n330), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n390), .B(new_n391), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n382), .A2(new_n346), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(G200), .B2(new_n382), .ZN(new_n403));
  XOR2_X1   g0203(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n372), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n268), .A2(G232), .A3(new_n269), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n409));
  INV_X1    g0209(.A(G107), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n409), .C1(new_n410), .C2(new_n268), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n330), .ZN(new_n412));
  INV_X1    g0212(.A(new_n254), .ZN(new_n413));
  INV_X1    g0213(.A(G274), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n257), .A2(G244), .B1(new_n415), .B2(new_n261), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n412), .A2(G190), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n416), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G200), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n283), .A2(G77), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT74), .ZN(new_n421));
  INV_X1    g0221(.A(new_n290), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT15), .B(G87), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(KEYINPUT73), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(KEYINPUT73), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n423), .B1(new_n428), .B2(new_n297), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n282), .B1(new_n272), .B2(new_n312), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n417), .A2(new_n419), .A3(new_n421), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n421), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n412), .A2(new_n277), .A3(new_n416), .ZN(new_n433));
  INV_X1    g0233(.A(G169), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n418), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n396), .A2(new_n407), .A3(new_n431), .A4(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n311), .A2(new_n351), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT4), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1698), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n440), .A2(new_n357), .A3(new_n359), .A4(G244), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT80), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n268), .A2(KEYINPUT80), .A3(G244), .A4(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n357), .A2(new_n359), .A3(G244), .A4(new_n269), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n439), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n357), .A2(new_n359), .A3(G250), .A4(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n446), .A2(KEYINPUT79), .A3(new_n439), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n445), .A2(new_n449), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n330), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT81), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(KEYINPUT81), .A3(new_n330), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n255), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT82), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n459), .A2(new_n460), .B1(KEYINPUT5), .B2(new_n259), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n260), .A2(G1), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(KEYINPUT82), .C1(KEYINPUT5), .C2(new_n259), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G257), .A3(new_n254), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n415), .A2(new_n463), .A3(new_n461), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n457), .A2(new_n458), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G200), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n455), .A2(new_n467), .A3(G190), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n470), .A2(KEYINPUT83), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT6), .ZN(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n410), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n410), .A2(KEYINPUT6), .A3(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n287), .ZN(new_n479));
  OAI21_X1  g0279(.A(G107), .B1(new_n355), .B2(new_n361), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n282), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n312), .A2(new_n473), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n255), .A2(G33), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n279), .A2(new_n484), .A3(new_n227), .A4(new_n281), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n473), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(KEYINPUT83), .B2(new_n470), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n469), .A2(new_n471), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n486), .B1(new_n481), .B2(new_n282), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n455), .A2(new_n467), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n434), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n465), .A2(new_n277), .A3(new_n466), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n457), .A2(new_n458), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n413), .B1(new_n461), .B2(new_n463), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n459), .A2(new_n460), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n463), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(G270), .A2(new_n499), .B1(new_n502), .B2(new_n415), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n360), .A2(G303), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n357), .A2(new_n359), .A3(G264), .A4(G1698), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n357), .A2(new_n359), .A3(G257), .A4(new_n269), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n504), .A2(KEYINPUT86), .A3(new_n505), .A4(new_n506), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n330), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n503), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G200), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n451), .B(new_n228), .C1(G33), .C2(new_n473), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G20), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n282), .A2(KEYINPUT88), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT88), .B1(new_n282), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT20), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(KEYINPUT20), .B(new_n514), .C1(new_n517), .C2(new_n518), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OR3_X1    g0323(.A1(new_n485), .A2(KEYINPUT87), .A3(new_n515), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT87), .B1(new_n485), .B2(new_n515), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n524), .A2(new_n525), .B1(new_n515), .B2(new_n312), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n513), .A2(KEYINPUT90), .A3(new_n523), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT90), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n304), .B1(new_n503), .B2(new_n511), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n523), .A2(new_n526), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n503), .A2(new_n511), .A3(G190), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n527), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n512), .A2(new_n277), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT21), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n523), .B2(new_n526), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n434), .B1(new_n503), .B2(new_n511), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n534), .A2(new_n530), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n530), .ZN(new_n539));
  XOR2_X1   g0339(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT23), .B1(new_n228), .B2(G107), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT23), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(new_n410), .A3(G20), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n228), .A2(G33), .A3(G116), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT91), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n544), .A2(new_n546), .A3(new_n547), .A4(KEYINPUT91), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n357), .A2(new_n359), .A3(new_n228), .A4(G87), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT22), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n268), .A2(new_n555), .A3(new_n228), .A4(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT24), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n552), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n300), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT25), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n279), .B2(G107), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n279), .A2(new_n563), .A3(G107), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n565), .A2(new_n566), .B1(new_n410), .B2(new_n485), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT92), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n561), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n560), .B1(new_n552), .B2(new_n557), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n282), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT92), .ZN(new_n572));
  INV_X1    g0372(.A(new_n567), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n268), .A2(G250), .A3(new_n269), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G294), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n330), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n464), .A2(G264), .A3(new_n254), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(new_n466), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G169), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n277), .B2(new_n581), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n568), .A2(new_n574), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n581), .A2(new_n346), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(G200), .B2(new_n581), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n562), .A2(new_n567), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n357), .A2(new_n359), .A3(G244), .A4(G1698), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n357), .A2(new_n359), .A3(G238), .A4(new_n269), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G116), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n330), .ZN(new_n593));
  INV_X1    g0393(.A(G250), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n260), .B2(G1), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n255), .A2(new_n414), .A3(G45), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n254), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G169), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(G179), .A3(new_n598), .ZN(new_n601));
  INV_X1    g0401(.A(new_n427), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n312), .B1(new_n602), .B2(new_n425), .ZN(new_n603));
  INV_X1    g0403(.A(new_n485), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n426), .A2(new_n604), .A3(new_n427), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n228), .B1(new_n328), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G87), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n475), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n357), .A2(new_n359), .A3(new_n228), .A4(G68), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n606), .B1(new_n297), .B2(new_n473), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n282), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n603), .A2(new_n605), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT84), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n600), .A2(new_n601), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n599), .A2(G200), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n279), .A2(new_n484), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n620), .A2(KEYINPUT85), .A3(new_n300), .A4(G87), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n485), .B2(new_n608), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n603), .A3(new_n614), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n346), .B(new_n597), .C1(new_n592), .C2(new_n330), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n617), .A2(new_n618), .B1(new_n619), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n584), .A2(new_n588), .A3(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n438), .A2(new_n498), .A3(new_n543), .A4(new_n629), .ZN(G372));
  NAND2_X1  g0430(.A1(new_n385), .A2(new_n395), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n344), .B1(new_n349), .B2(new_n436), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n407), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n309), .A2(new_n310), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n303), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n465), .A2(new_n466), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n330), .B2(new_n454), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n488), .B1(new_n638), .B2(G169), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n454), .A2(KEYINPUT81), .A3(new_n330), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT81), .B1(new_n454), .B2(new_n330), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n640), .A2(new_n641), .A3(new_n494), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n636), .B1(new_n643), .B2(new_n628), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n597), .B1(new_n592), .B2(new_n330), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n601), .B1(new_n434), .B2(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n627), .A2(new_n619), .B1(new_n646), .B2(new_n615), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n493), .A2(new_n647), .A3(new_n496), .A4(new_n636), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n615), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n583), .B1(new_n562), .B2(new_n567), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n538), .A3(new_n541), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n627), .A2(new_n619), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n649), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n586), .B2(new_n587), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n653), .A2(new_n490), .A3(new_n656), .A4(new_n497), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n635), .B1(new_n438), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT93), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n255), .A2(new_n228), .A3(G13), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n530), .A2(new_n666), .ZN(new_n667));
  MUX2_X1   g0467(.A(new_n542), .B(new_n543), .S(new_n667), .Z(new_n668));
  INV_X1    g0468(.A(KEYINPUT94), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n666), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n584), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n568), .A2(new_n574), .A3(new_n666), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n584), .A2(new_n673), .A3(new_n588), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n670), .A2(G330), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n542), .A2(new_n671), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n584), .A2(new_n588), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n652), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n671), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n681), .ZN(G399));
  NOR2_X1   g0482(.A1(new_n223), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n475), .A2(new_n608), .A3(new_n515), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n255), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n230), .B2(new_n684), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  INV_X1    g0490(.A(new_n657), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n628), .A2(new_n496), .A3(new_n493), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n649), .B(new_n648), .C1(new_n692), .C2(new_n636), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n690), .B(new_n671), .C1(new_n691), .C2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n493), .A2(new_n647), .A3(new_n496), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT26), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n628), .A2(new_n636), .A3(new_n496), .A4(new_n493), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n696), .A2(new_n649), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n584), .A2(new_n541), .A3(new_n538), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n497), .A3(new_n490), .A4(new_n656), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n666), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n694), .B1(new_n690), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n498), .A2(new_n543), .A3(new_n629), .A4(new_n671), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n645), .A2(G179), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n468), .A2(new_n512), .A3(new_n581), .A4(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  INV_X1    g0506(.A(new_n601), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n499), .A2(G264), .B1(new_n578), .B2(new_n330), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n503), .A3(new_n708), .A4(new_n511), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n706), .B1(new_n709), .B2(new_n492), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT30), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n706), .B(new_n712), .C1(new_n709), .C2(new_n492), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n705), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n666), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n703), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n702), .B1(G330), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n689), .B1(new_n720), .B2(G1), .ZN(G364));
  NAND2_X1  g0521(.A1(new_n670), .A2(G330), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n220), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n255), .B1(new_n724), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n683), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G330), .B2(new_n670), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n265), .B1(new_n228), .B2(G169), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT97), .Z(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n245), .A2(new_n260), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n224), .A2(new_n360), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n737), .B(new_n738), .C1(new_n260), .C2(new_n231), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n224), .A2(G355), .A3(new_n268), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G116), .B2(new_n224), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n736), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n727), .B(KEYINPUT96), .Z(new_n743));
  NOR2_X1   g0543(.A1(new_n228), .A2(new_n346), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(new_n277), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n608), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n360), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT99), .Z(new_n748));
  NOR2_X1   g0548(.A1(new_n228), .A2(G190), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(new_n277), .A3(new_n304), .ZN(new_n750));
  INV_X1    g0550(.A(G159), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT32), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n277), .A2(G200), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n744), .A2(KEYINPUT98), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT98), .B1(new_n744), .B2(new_n753), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n748), .B(new_n752), .C1(new_n293), .C2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n346), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n228), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n228), .A2(new_n277), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G97), .A2(new_n760), .B1(new_n763), .B2(G50), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n761), .A2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n749), .A2(new_n753), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n766), .A2(G68), .B1(new_n768), .B2(G77), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n749), .A2(new_n277), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G107), .ZN(new_n772));
  OR3_X1    g0572(.A1(new_n750), .A2(KEYINPUT32), .A3(new_n751), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n764), .A2(new_n769), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G283), .ZN(new_n775));
  INV_X1    g0575(.A(G329), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n770), .B1(new_n750), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n777), .B1(new_n766), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n360), .B1(new_n767), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n745), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(G303), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G322), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n779), .B(new_n783), .C1(new_n784), .C2(new_n756), .ZN(new_n785));
  INV_X1    g0585(.A(G294), .ZN(new_n786));
  INV_X1    g0586(.A(G326), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n759), .A2(new_n786), .B1(new_n762), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT100), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n757), .A2(new_n774), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n732), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n742), .A2(new_n743), .A3(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT101), .Z(new_n793));
  INV_X1    g0593(.A(new_n735), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n668), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n729), .A2(new_n795), .ZN(G396));
  AOI21_X1  g0596(.A(new_n666), .B1(new_n651), .B2(new_n657), .ZN(new_n797));
  INV_X1    g0597(.A(new_n436), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n671), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n432), .A2(new_n666), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n431), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n436), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n797), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n719), .A2(G330), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n727), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n763), .A2(G137), .B1(new_n768), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(new_n766), .ZN(new_n811));
  INV_X1    g0611(.A(G143), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n811), .B2(new_n286), .C1(new_n812), .C2(new_n756), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT34), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n268), .B1(new_n745), .B2(new_n318), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n313), .A2(new_n770), .B1(new_n750), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(G58), .C2(new_n760), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n762), .A2(new_n819), .B1(new_n750), .B2(new_n780), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G87), .B2(new_n771), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n360), .B1(new_n767), .B2(new_n515), .C1(new_n745), .C2(new_n410), .ZN(new_n822));
  XOR2_X1   g0622(.A(KEYINPUT103), .B(G283), .Z(new_n823));
  OAI22_X1  g0623(.A1(new_n811), .A2(new_n823), .B1(new_n473), .B2(new_n759), .ZN(new_n824));
  INV_X1    g0624(.A(new_n756), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n822), .B(new_n824), .C1(G294), .C2(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n814), .A2(new_n818), .B1(new_n821), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n731), .B1(new_n827), .B2(KEYINPUT104), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(KEYINPUT104), .B2(new_n827), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n731), .A2(new_n734), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT102), .Z(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n743), .C1(G77), .C2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n733), .B2(new_n803), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n809), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G384));
  OR2_X1    g0635(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n836), .A2(G116), .A3(new_n229), .A4(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT36), .Z(new_n839));
  OR3_X1    g0639(.A1(new_n230), .A2(new_n272), .A3(new_n363), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n318), .A2(G68), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n255), .B(G13), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  INV_X1    g0644(.A(new_n664), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n392), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n396), .B2(new_n407), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n392), .A2(new_n383), .A3(new_n394), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n848), .A2(new_n849), .A3(new_n399), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT105), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n392), .B2(new_n845), .ZN(new_n852));
  AOI211_X1 g0652(.A(KEYINPUT105), .B(new_n664), .C1(new_n390), .C2(new_n391), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n848), .A2(new_n399), .A3(new_n846), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n850), .A2(new_n854), .B1(new_n855), .B2(KEYINPUT37), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n844), .B1(new_n847), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n846), .A2(KEYINPUT105), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n392), .A2(new_n851), .A3(new_n845), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n848), .A2(new_n849), .A3(new_n399), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n846), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n401), .A2(new_n406), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(new_n631), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n863), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n857), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n344), .B(new_n350), .C1(new_n345), .C2(new_n671), .ZN(new_n869));
  INV_X1    g0669(.A(new_n343), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n341), .A3(new_n340), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n325), .B(new_n666), .C1(new_n871), .C2(new_n349), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n666), .B(new_n803), .C1(new_n651), .C2(new_n657), .ZN(new_n874));
  INV_X1    g0674(.A(new_n799), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n868), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n631), .A2(new_n664), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n854), .B1(new_n396), .B2(new_n407), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT108), .B1(new_n861), .B2(new_n862), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT108), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n850), .A2(new_n882), .A3(new_n854), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n399), .B1(new_n372), .B2(new_n384), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT107), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT107), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n848), .A2(new_n887), .A3(new_n399), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n854), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n880), .B1(new_n891), .B2(KEYINPUT109), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n881), .A2(new_n883), .B1(new_n889), .B2(KEYINPUT37), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT109), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n867), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n879), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n871), .A2(new_n325), .A3(new_n671), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT106), .Z(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n878), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n635), .B1(new_n702), .B2(new_n438), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n903), .B(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n803), .B1(new_n869), .B2(new_n872), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n868), .A2(new_n719), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n892), .A2(new_n895), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n897), .B1(new_n910), .B2(new_n844), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n719), .A2(new_n906), .A3(KEYINPUT40), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n438), .A2(new_n719), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(G330), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n905), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n255), .B2(new_n724), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n905), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n843), .B1(new_n919), .B2(new_n920), .ZN(G367));
  OAI211_X1 g0721(.A(new_n490), .B(new_n497), .C1(new_n491), .C2(new_n671), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n643), .A2(new_n666), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n679), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n625), .A2(new_n666), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n649), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n647), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n497), .B1(new_n922), .B2(new_n584), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n925), .A2(KEYINPUT42), .B1(new_n934), .B2(new_n671), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n929), .A2(new_n930), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n927), .B2(new_n928), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n933), .A2(new_n930), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n933), .A2(new_n930), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n676), .B1(new_n922), .B2(new_n923), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n936), .B2(new_n940), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n683), .B(KEYINPUT41), .Z(new_n945));
  NOR2_X1   g0745(.A1(new_n681), .A2(new_n924), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n681), .A2(new_n924), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT45), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT111), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n676), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n720), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n672), .A2(new_n677), .A3(new_n674), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT112), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n679), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n677), .A2(KEYINPUT112), .A3(new_n678), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n722), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n670), .B(G330), .C1(new_n958), .C2(new_n957), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n954), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n947), .A2(new_n950), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n963), .A2(KEYINPUT111), .A3(new_n723), .A4(new_n675), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n953), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n945), .B1(new_n965), .B2(new_n720), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n944), .B1(new_n966), .B2(new_n726), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n360), .B1(new_n823), .B2(new_n767), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n745), .A2(new_n515), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT46), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n968), .B(new_n970), .C1(G294), .C2(new_n766), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n771), .A2(G97), .ZN(new_n972));
  INV_X1    g0772(.A(G317), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n973), .B2(new_n750), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n759), .A2(new_n410), .B1(new_n762), .B2(new_n780), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n971), .B(new_n976), .C1(new_n819), .C2(new_n756), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n770), .A2(new_n272), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n268), .B1(new_n767), .B2(new_n318), .C1(new_n745), .C2(new_n293), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(G159), .C2(new_n766), .ZN(new_n980));
  INV_X1    g0780(.A(G137), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n750), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n759), .A2(new_n313), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(G143), .C2(new_n763), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n980), .B(new_n984), .C1(new_n286), .C2(new_n756), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n731), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n986), .B2(new_n987), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n933), .A2(new_n735), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n736), .B1(new_n224), .B2(new_n428), .C1(new_n237), .C2(new_n738), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n989), .A2(new_n743), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n967), .A2(new_n992), .ZN(G387));
  INV_X1    g0793(.A(new_n962), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n960), .A2(new_n954), .A3(new_n961), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n683), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n960), .A2(new_n961), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n726), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n675), .A2(new_n794), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n360), .B1(new_n770), .B2(new_n515), .C1(new_n787), .C2(new_n750), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n766), .A2(G311), .B1(new_n768), .B2(G303), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n784), .B2(new_n762), .C1(new_n973), .C2(new_n756), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT114), .Z(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n759), .A2(new_n823), .B1(new_n745), .B2(new_n786), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT49), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(KEYINPUT49), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n972), .B1(new_n286), .B2(new_n750), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n745), .A2(new_n272), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n360), .B(new_n1013), .C1(G68), .C2(new_n768), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n825), .A2(G50), .B1(new_n296), .B2(new_n766), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n428), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n760), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1012), .B(new_n1018), .C1(G159), .C2(new_n763), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n732), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n241), .A2(new_n260), .A3(new_n268), .ZN(new_n1021));
  OR3_X1    g0821(.A1(new_n290), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT50), .B1(new_n290), .B2(G50), .ZN(new_n1023));
  AOI21_X1  g0823(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n685), .B1(new_n1025), .B2(new_n360), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1021), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1027), .A2(new_n223), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n736), .B1(new_n224), .B2(new_n410), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1020), .B(new_n743), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n996), .B(new_n998), .C1(new_n999), .C2(new_n1030), .ZN(G393));
  NAND2_X1  g0831(.A1(new_n965), .A2(new_n683), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT115), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n676), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n676), .A2(new_n1033), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n951), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n963), .A2(new_n1033), .A3(new_n676), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(KEYINPUT117), .B1(new_n1038), .B2(new_n962), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT117), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n994), .A3(new_n1040), .A4(new_n1037), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1032), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1038), .A2(new_n726), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n736), .B1(new_n473), .B2(new_n224), .C1(new_n738), .C2(new_n248), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n743), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n360), .B1(new_n782), .B2(G68), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n608), .B2(new_n770), .C1(new_n812), .C2(new_n750), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1047), .A2(KEYINPUT116), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(KEYINPUT116), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n811), .A2(new_n318), .B1(new_n290), .B2(new_n767), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G77), .B2(new_n760), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n756), .A2(new_n751), .B1(new_n286), .B2(new_n762), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT51), .Z(new_n1054));
  OAI22_X1  g0854(.A1(new_n756), .A2(new_n780), .B1(new_n973), .B2(new_n762), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  OAI21_X1  g0856(.A(new_n772), .B1(new_n811), .B2(new_n819), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n360), .B1(new_n767), .B2(new_n786), .C1(new_n745), .C2(new_n823), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n759), .A2(new_n515), .B1(new_n750), .B2(new_n784), .ZN(new_n1059));
  OR3_X1    g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1052), .A2(new_n1054), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1045), .B1(new_n732), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n924), .B2(new_n794), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1043), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1042), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(G390));
  INV_X1    g0866(.A(new_n880), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n893), .B2(new_n894), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n884), .A2(new_n894), .A3(new_n890), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n844), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n867), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n802), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n666), .B(new_n1072), .C1(new_n698), .C2(new_n700), .ZN(new_n1073));
  OAI21_X1  g0873(.A(KEYINPUT118), .B1(new_n1073), .B2(new_n875), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n698), .A2(new_n700), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n671), .A3(new_n802), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT118), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n799), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1074), .A2(new_n873), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1071), .A2(new_n1079), .A3(new_n901), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n875), .B1(new_n797), .B2(new_n804), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n873), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n901), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1083), .B(new_n879), .C1(new_n896), .C2(new_n898), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n719), .A2(G330), .A3(new_n804), .A4(new_n873), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1080), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n899), .A2(new_n734), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(KEYINPUT54), .B(G143), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n268), .B1(new_n767), .B2(new_n1090), .C1(new_n318), .C2(new_n770), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n811), .A2(new_n981), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n750), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1091), .B(new_n1092), .C1(G125), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n782), .A2(G150), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT53), .ZN(new_n1096));
  INV_X1    g0896(.A(G128), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n759), .A2(new_n751), .B1(new_n762), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1094), .B(new_n1099), .C1(new_n816), .C2(new_n756), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n811), .A2(new_n410), .B1(new_n786), .B2(new_n750), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G283), .B2(new_n763), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n825), .A2(G116), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n268), .B(new_n746), .C1(G97), .C2(new_n768), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n760), .A2(G77), .B1(new_n771), .B2(G68), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n731), .B1(new_n1100), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n743), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n831), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1107), .B(new_n1108), .C1(new_n295), .C2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1088), .A2(new_n726), .B1(new_n1089), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1085), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1080), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n701), .A2(new_n690), .ZN(new_n1117));
  AOI211_X1 g0917(.A(KEYINPUT29), .B(new_n666), .C1(new_n651), .C2(new_n657), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n438), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n635), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n438), .A2(new_n719), .A3(G330), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(KEYINPUT119), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT119), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n904), .B2(new_n1121), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n719), .A2(G330), .A3(new_n804), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1082), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n1085), .A3(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1129), .A2(new_n1085), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n1081), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT120), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n683), .B1(new_n1116), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT120), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1081), .B1(new_n1129), .B2(new_n1085), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1122), .A2(KEYINPUT119), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n904), .A2(new_n1124), .A3(new_n1121), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1135), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1088), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1111), .B1(new_n1134), .B2(new_n1142), .ZN(G378));
  NAND3_X1  g0943(.A1(new_n311), .A2(new_n301), .A3(new_n845), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n301), .A2(new_n845), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n303), .B(new_n1145), .C1(new_n309), .C2(new_n310), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n912), .B1(new_n1070), .B2(new_n867), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n909), .A2(G330), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(G330), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n907), .B2(new_n908), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1158), .B(new_n1152), .C1(new_n911), .C2(new_n912), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n903), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n903), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1153), .A2(new_n733), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n727), .B1(new_n831), .B2(G50), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n360), .A2(new_n259), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1167), .B(new_n318), .C1(G33), .C2(G41), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n811), .A2(new_n473), .B1(new_n775), .B2(new_n750), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n762), .A2(new_n515), .B1(new_n770), .B2(new_n293), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1016), .A2(new_n768), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n825), .A2(G107), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n983), .A2(new_n1013), .A3(new_n1167), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1168), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT122), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n745), .A2(new_n1090), .B1(new_n767), .B2(new_n981), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G132), .B2(new_n766), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G150), .A2(new_n760), .B1(new_n763), .B2(G125), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n1097), .C2(new_n756), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G33), .B(G41), .C1(new_n1093), .C2(G124), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n751), .B2(new_n770), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1186), .B2(KEYINPUT59), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1178), .A2(new_n1176), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1181), .A2(new_n1182), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1166), .B1(new_n1192), .B2(new_n732), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1164), .A2(new_n726), .B1(new_n1165), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1140), .B1(new_n1088), .B2(new_n1132), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n903), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n899), .A2(new_n902), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n878), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1156), .A2(new_n1159), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n683), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1114), .A2(new_n1115), .A3(new_n1132), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1126), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1164), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1194), .B1(new_n1201), .B2(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n1082), .A2(new_n733), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n811), .A2(new_n1090), .B1(new_n816), .B2(new_n762), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G50), .B2(new_n760), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n268), .B1(new_n767), .B2(new_n286), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G159), .B2(new_n782), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n825), .A2(G137), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n771), .A2(G58), .B1(new_n1093), .B2(G128), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1208), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n762), .A2(new_n786), .B1(new_n750), .B2(new_n819), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n978), .B(new_n1214), .C1(G116), .C2(new_n766), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n825), .A2(G283), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n360), .B1(new_n767), .B2(new_n410), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G97), .B2(new_n782), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1017), .A3(new_n1216), .A4(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n731), .B1(new_n1213), .B2(new_n1219), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1220), .B(new_n1108), .C1(new_n313), .C2(new_n1109), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT123), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1132), .A2(new_n726), .B1(new_n1206), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n945), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1223), .B1(new_n1225), .B2(new_n1227), .ZN(G381));
  INV_X1    g1028(.A(G387), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1089), .A2(new_n1110), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1116), .B2(new_n725), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1142), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n684), .B1(new_n1088), .B2(new_n1141), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1231), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1229), .A2(new_n1065), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1236), .A2(G375), .ZN(G407));
  OAI21_X1  g1037(.A(G213), .B1(new_n1236), .B2(G375), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n665), .A2(G213), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(G375), .A2(G378), .A3(new_n1239), .ZN(new_n1240));
  OR3_X1    g1040(.A1(new_n1238), .A2(new_n1240), .A3(KEYINPUT124), .ZN(new_n1241));
  OAI21_X1  g1041(.A(KEYINPUT124), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(G409));
  NAND2_X1  g1043(.A1(G387), .A2(new_n1065), .ZN(new_n1244));
  XOR2_X1   g1044(.A(G393), .B(G396), .Z(new_n1245));
  OAI211_X1 g1045(.A(new_n967), .B(new_n992), .C1(new_n1042), .C2(new_n1064), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1245), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1194), .C1(new_n1201), .C2(new_n1204), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1203), .A2(new_n1224), .A3(new_n1164), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1194), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1234), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT60), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1226), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n1140), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n683), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(G384), .A3(new_n1223), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1258), .B2(new_n1223), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1254), .A2(new_n1239), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  XOR2_X1   g1064(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1265));
  AOI22_X1  g1065(.A1(new_n1250), .A2(new_n1253), .B1(G213), .B2(new_n665), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1255), .A2(new_n1226), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1257), .A2(new_n683), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1223), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n834), .ZN(new_n1270));
  INV_X1    g1070(.A(G2897), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1239), .A2(new_n1271), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1270), .A2(new_n1259), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1272), .B1(new_n1270), .B2(new_n1259), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1264), .B(new_n1265), .C1(new_n1266), .C2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(new_n1266), .B2(new_n1262), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1249), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1247), .A2(new_n1248), .A3(KEYINPUT61), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1254), .A2(new_n1239), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1262), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT125), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n1260), .A2(new_n1261), .B1(new_n1271), .B2(new_n1239), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1270), .A2(new_n1259), .A3(new_n1272), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1286), .A2(new_n1290), .A3(new_n1283), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1262), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1281), .A2(new_n1285), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1280), .A2(new_n1293), .ZN(G405));
  NAND2_X1  g1094(.A1(G375), .A2(new_n1234), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1284), .A2(new_n1250), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1284), .B1(new_n1295), .B2(new_n1250), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1249), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1298), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1301), .A3(new_n1296), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(G402));
endmodule


