

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n579), .A2(n516), .ZN(G164) );
  XNOR2_X2 U549 ( .A(n739), .B(KEYINPUT32), .ZN(n762) );
  NOR2_X1 U550 ( .A1(n770), .A2(n751), .ZN(n753) );
  NOR2_X1 U551 ( .A1(n742), .A2(n722), .ZN(n724) );
  OR2_X1 U552 ( .A1(n697), .A2(n970), .ZN(n698) );
  INV_X1 U553 ( .A(KEYINPUT64), .ZN(n752) );
  INV_X1 U554 ( .A(KEYINPUT23), .ZN(n518) );
  INV_X1 U555 ( .A(KEYINPUT101), .ZN(n700) );
  NAND2_X1 U556 ( .A1(n773), .A2(n772), .ZN(n805) );
  AND2_X1 U557 ( .A1(n771), .A2(n514), .ZN(n772) );
  NOR2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  NOR2_X2 U559 ( .A1(n533), .A2(n532), .ZN(G160) );
  XNOR2_X2 U560 ( .A(n527), .B(KEYINPUT67), .ZN(n575) );
  XOR2_X1 U561 ( .A(n729), .B(KEYINPUT31), .Z(n513) );
  OR2_X1 U562 ( .A1(n770), .A2(n769), .ZN(n514) );
  AND2_X1 U563 ( .A1(n813), .A2(n804), .ZN(n515) );
  XOR2_X1 U564 ( .A(n578), .B(KEYINPUT93), .Z(n516) );
  OR2_X1 U565 ( .A1(n721), .A2(n740), .ZN(n722) );
  INV_X1 U566 ( .A(KEYINPUT30), .ZN(n723) );
  INV_X1 U567 ( .A(KEYINPUT103), .ZN(n736) );
  INV_X1 U568 ( .A(KEYINPUT97), .ZN(n719) );
  NOR2_X1 U569 ( .A1(n684), .A2(n774), .ZN(n687) );
  INV_X1 U570 ( .A(n687), .ZN(n718) );
  INV_X1 U571 ( .A(KEYINPUT33), .ZN(n754) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n524) );
  XNOR2_X1 U573 ( .A(n524), .B(KEYINPUT68), .ZN(n525) );
  XNOR2_X1 U574 ( .A(n519), .B(n518), .ZN(n522) );
  NOR2_X1 U575 ( .A1(n632), .A2(G651), .ZN(n649) );
  NAND2_X1 U576 ( .A1(n520), .A2(G2104), .ZN(n517) );
  XNOR2_X1 U577 ( .A(n517), .B(KEYINPUT65), .ZN(n571) );
  NAND2_X1 U578 ( .A1(n571), .A2(G101), .ZN(n519) );
  INV_X1 U579 ( .A(G2105), .ZN(n520) );
  NOR2_X4 U580 ( .A1(n520), .A2(G2104), .ZN(n883) );
  NAND2_X1 U581 ( .A1(n883), .A2(G125), .ZN(n521) );
  NAND2_X1 U582 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U583 ( .A(n523), .B(KEYINPUT66), .ZN(n533) );
  XNOR2_X2 U584 ( .A(n526), .B(n525), .ZN(n622) );
  NAND2_X1 U585 ( .A1(n622), .A2(G137), .ZN(n529) );
  NAND2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  NAND2_X1 U587 ( .A1(G113), .A2(n575), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n531) );
  INV_X1 U589 ( .A(KEYINPUT69), .ZN(n530) );
  XNOR2_X1 U590 ( .A(n531), .B(n530), .ZN(n532) );
  NOR2_X1 U591 ( .A1(G543), .A2(G651), .ZN(n654) );
  NAND2_X1 U592 ( .A1(n654), .A2(G89), .ZN(n534) );
  XNOR2_X1 U593 ( .A(n534), .B(KEYINPUT4), .ZN(n536) );
  XOR2_X1 U594 ( .A(KEYINPUT0), .B(G543), .Z(n632) );
  INV_X1 U595 ( .A(G651), .ZN(n538) );
  NOR2_X1 U596 ( .A1(n632), .A2(n538), .ZN(n651) );
  NAND2_X1 U597 ( .A1(G76), .A2(n651), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n537), .B(KEYINPUT5), .ZN(n545) );
  NOR2_X1 U600 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(n539), .Z(n650) );
  NAND2_X1 U602 ( .A1(n650), .A2(G63), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(KEYINPUT78), .ZN(n542) );
  NAND2_X1 U604 ( .A1(G51), .A2(n649), .ZN(n541) );
  NAND2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U606 ( .A(KEYINPUT6), .B(n543), .Z(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U608 ( .A(n546), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U609 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U610 ( .A(KEYINPUT9), .B(KEYINPUT71), .ZN(n550) );
  NAND2_X1 U611 ( .A1(G90), .A2(n654), .ZN(n548) );
  NAND2_X1 U612 ( .A1(G77), .A2(n651), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n649), .A2(G52), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n551), .B(KEYINPUT70), .ZN(n553) );
  NAND2_X1 U617 ( .A1(G64), .A2(n650), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT72), .B(n556), .Z(G301) );
  INV_X1 U621 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U622 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U623 ( .A(G57), .ZN(G237) );
  NAND2_X1 U624 ( .A1(G132), .A2(G82), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT22), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(KEYINPUT88), .ZN(n559) );
  NOR2_X1 U627 ( .A1(G218), .A2(n559), .ZN(n560) );
  NAND2_X1 U628 ( .A1(G96), .A2(n560), .ZN(n826) );
  NAND2_X1 U629 ( .A1(n826), .A2(G2106), .ZN(n564) );
  NAND2_X1 U630 ( .A1(G108), .A2(G120), .ZN(n561) );
  NOR2_X1 U631 ( .A1(G237), .A2(n561), .ZN(n562) );
  NAND2_X1 U632 ( .A1(G69), .A2(n562), .ZN(n825) );
  NAND2_X1 U633 ( .A1(G567), .A2(n825), .ZN(n563) );
  AND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(G319) );
  NAND2_X1 U635 ( .A1(G85), .A2(n654), .ZN(n566) );
  NAND2_X1 U636 ( .A1(G72), .A2(n651), .ZN(n565) );
  NAND2_X1 U637 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G60), .A2(n650), .ZN(n568) );
  NAND2_X1 U639 ( .A1(G47), .A2(n649), .ZN(n567) );
  NAND2_X1 U640 ( .A1(n568), .A2(n567), .ZN(n569) );
  OR2_X1 U641 ( .A1(n570), .A2(n569), .ZN(G290) );
  BUF_X1 U642 ( .A(n571), .Z(n886) );
  NAND2_X1 U643 ( .A1(n886), .A2(G102), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G138), .A2(n622), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n883), .A2(G126), .ZN(n574) );
  XNOR2_X1 U647 ( .A(n574), .B(KEYINPUT92), .ZN(n577) );
  NAND2_X1 U648 ( .A1(G114), .A2(n575), .ZN(n576) );
  NAND2_X1 U649 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U650 ( .A1(G94), .A2(G452), .ZN(n580) );
  XNOR2_X1 U651 ( .A(n580), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n581) );
  XOR2_X1 U653 ( .A(n581), .B(KEYINPUT10), .Z(n917) );
  NAND2_X1 U654 ( .A1(n917), .A2(G567), .ZN(n582) );
  XOR2_X1 U655 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  NAND2_X1 U656 ( .A1(n650), .A2(G56), .ZN(n583) );
  XNOR2_X1 U657 ( .A(KEYINPUT14), .B(n583), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n654), .A2(G81), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U660 ( .A1(G68), .A2(n651), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U662 ( .A(KEYINPUT13), .B(n587), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U664 ( .A(n590), .B(KEYINPUT75), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n649), .A2(G43), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n980) );
  XOR2_X1 U667 ( .A(G860), .B(KEYINPUT76), .Z(n612) );
  NOR2_X1 U668 ( .A1(n980), .A2(n612), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT77), .ZN(G153) );
  NAND2_X1 U670 ( .A1(G301), .A2(G868), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G66), .A2(n650), .ZN(n595) );
  NAND2_X1 U672 ( .A1(G92), .A2(n654), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G79), .A2(n651), .ZN(n597) );
  NAND2_X1 U675 ( .A1(G54), .A2(n649), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U678 ( .A(KEYINPUT15), .B(n600), .ZN(n613) );
  INV_X1 U679 ( .A(G868), .ZN(n672) );
  NAND2_X1 U680 ( .A1(n613), .A2(n672), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n602), .A2(n601), .ZN(G284) );
  NAND2_X1 U682 ( .A1(G91), .A2(n654), .ZN(n604) );
  NAND2_X1 U683 ( .A1(G78), .A2(n651), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n649), .A2(G53), .ZN(n605) );
  XOR2_X1 U686 ( .A(KEYINPUT74), .B(n605), .Z(n606) );
  NOR2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n650), .A2(G65), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(G299) );
  NOR2_X1 U690 ( .A1(G286), .A2(n672), .ZN(n611) );
  NOR2_X1 U691 ( .A1(G868), .A2(G299), .ZN(n610) );
  NOR2_X1 U692 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n612), .A2(G559), .ZN(n614) );
  INV_X1 U694 ( .A(n613), .ZN(n970) );
  NAND2_X1 U695 ( .A1(n614), .A2(n970), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U697 ( .A1(G868), .A2(n980), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n970), .A2(G868), .ZN(n616) );
  NOR2_X1 U699 ( .A1(G559), .A2(n616), .ZN(n617) );
  NOR2_X1 U700 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U701 ( .A1(n883), .A2(G123), .ZN(n619) );
  XNOR2_X1 U702 ( .A(n619), .B(KEYINPUT18), .ZN(n621) );
  NAND2_X1 U703 ( .A1(G111), .A2(n575), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n886), .A2(G99), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G135), .A2(n622), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n924) );
  XNOR2_X1 U709 ( .A(G2096), .B(n924), .ZN(n627) );
  INV_X1 U710 ( .A(G2100), .ZN(n836) );
  NAND2_X1 U711 ( .A1(n627), .A2(n836), .ZN(G156) );
  NAND2_X1 U712 ( .A1(G49), .A2(n649), .ZN(n629) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U715 ( .A(KEYINPUT83), .B(n630), .Z(n631) );
  NOR2_X1 U716 ( .A1(n650), .A2(n631), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n632), .A2(G87), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U719 ( .A1(G61), .A2(n650), .ZN(n636) );
  NAND2_X1 U720 ( .A1(G86), .A2(n654), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n651), .A2(G73), .ZN(n637) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n637), .Z(n638) );
  NOR2_X1 U724 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n649), .A2(G48), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G88), .A2(n654), .ZN(n643) );
  NAND2_X1 U728 ( .A1(G75), .A2(n651), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n650), .A2(G62), .ZN(n644) );
  XOR2_X1 U731 ( .A(KEYINPUT84), .B(n644), .Z(n645) );
  NOR2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n649), .A2(G50), .ZN(n647) );
  NAND2_X1 U734 ( .A1(n648), .A2(n647), .ZN(G303) );
  INV_X1 U735 ( .A(G303), .ZN(G166) );
  NAND2_X1 U736 ( .A1(G55), .A2(n649), .ZN(n659) );
  NAND2_X1 U737 ( .A1(G67), .A2(n650), .ZN(n653) );
  NAND2_X1 U738 ( .A1(G80), .A2(n651), .ZN(n652) );
  NAND2_X1 U739 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n654), .A2(G93), .ZN(n655) );
  XOR2_X1 U741 ( .A(KEYINPUT80), .B(n655), .Z(n656) );
  NOR2_X1 U742 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U743 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U744 ( .A(n660), .B(KEYINPUT81), .Z(n828) );
  XNOR2_X1 U745 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n662) );
  XNOR2_X1 U746 ( .A(G290), .B(KEYINPUT19), .ZN(n661) );
  XNOR2_X1 U747 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U748 ( .A(n828), .B(n663), .ZN(n664) );
  XNOR2_X1 U749 ( .A(G305), .B(n664), .ZN(n665) );
  XNOR2_X1 U750 ( .A(G288), .B(n665), .ZN(n667) );
  XOR2_X1 U751 ( .A(G299), .B(G166), .Z(n666) );
  XNOR2_X1 U752 ( .A(n667), .B(n666), .ZN(n851) );
  XNOR2_X1 U753 ( .A(n851), .B(KEYINPUT87), .ZN(n670) );
  XNOR2_X1 U754 ( .A(n980), .B(KEYINPUT79), .ZN(n669) );
  NAND2_X1 U755 ( .A1(n970), .A2(G559), .ZN(n668) );
  XOR2_X1 U756 ( .A(n669), .B(n668), .Z(n827) );
  XOR2_X1 U757 ( .A(n670), .B(n827), .Z(n671) );
  NAND2_X1 U758 ( .A1(n671), .A2(G868), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n828), .A2(n672), .ZN(n673) );
  NAND2_X1 U760 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U761 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U762 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U763 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U764 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n678), .A2(G2072), .ZN(G158) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n679) );
  XNOR2_X1 U767 ( .A(KEYINPUT89), .B(n679), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n680), .A2(G319), .ZN(n681) );
  XOR2_X1 U769 ( .A(KEYINPUT90), .B(n681), .Z(n824) );
  NAND2_X1 U770 ( .A1(n824), .A2(G36), .ZN(n682) );
  XOR2_X1 U771 ( .A(KEYINPUT91), .B(n682), .Z(G176) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n775) );
  INV_X1 U773 ( .A(n775), .ZN(n684) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n774) );
  NAND2_X1 U775 ( .A1(G8), .A2(n718), .ZN(n770) );
  INV_X1 U776 ( .A(G1961), .ZN(n987) );
  NAND2_X1 U777 ( .A1(n718), .A2(n987), .ZN(n686) );
  INV_X1 U778 ( .A(n718), .ZN(n703) );
  XNOR2_X1 U779 ( .A(G2078), .B(KEYINPUT25), .ZN(n946) );
  NAND2_X1 U780 ( .A1(n703), .A2(n946), .ZN(n685) );
  NAND2_X1 U781 ( .A1(n686), .A2(n685), .ZN(n726) );
  NAND2_X1 U782 ( .A1(n726), .A2(G171), .ZN(n716) );
  NAND2_X1 U783 ( .A1(G1996), .A2(n687), .ZN(n688) );
  XNOR2_X1 U784 ( .A(n688), .B(KEYINPUT26), .ZN(n690) );
  NAND2_X1 U785 ( .A1(G1341), .A2(n718), .ZN(n689) );
  NAND2_X1 U786 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U787 ( .A(n691), .B(KEYINPUT100), .ZN(n692) );
  NOR2_X1 U788 ( .A1(n692), .A2(n980), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n697), .A2(n970), .ZN(n696) );
  NOR2_X1 U790 ( .A1(n703), .A2(G1348), .ZN(n694) );
  NOR2_X1 U791 ( .A1(G2067), .A2(n718), .ZN(n693) );
  NOR2_X1 U792 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U795 ( .A(n701), .B(n700), .ZN(n707) );
  NAND2_X1 U796 ( .A1(n703), .A2(G2072), .ZN(n702) );
  XNOR2_X1 U797 ( .A(n702), .B(KEYINPUT27), .ZN(n705) );
  XNOR2_X1 U798 ( .A(G1956), .B(KEYINPUT99), .ZN(n991) );
  NOR2_X1 U799 ( .A1(n991), .A2(n703), .ZN(n704) );
  NOR2_X1 U800 ( .A1(n705), .A2(n704), .ZN(n709) );
  INV_X1 U801 ( .A(G299), .ZN(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n712) );
  NOR2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U805 ( .A(n710), .B(KEYINPUT28), .Z(n711) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n714) );
  XOR2_X1 U807 ( .A(KEYINPUT102), .B(KEYINPUT29), .Z(n713) );
  XNOR2_X1 U808 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n730) );
  NOR2_X1 U810 ( .A1(n770), .A2(G1966), .ZN(n717) );
  XNOR2_X1 U811 ( .A(n717), .B(KEYINPUT98), .ZN(n742) );
  INV_X1 U812 ( .A(G8), .ZN(n721) );
  NOR2_X1 U813 ( .A1(n718), .A2(G2084), .ZN(n720) );
  XNOR2_X1 U814 ( .A(n720), .B(n719), .ZN(n740) );
  XNOR2_X1 U815 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U816 ( .A1(G168), .A2(n725), .ZN(n728) );
  NOR2_X1 U817 ( .A1(n726), .A2(G171), .ZN(n727) );
  NOR2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U819 ( .A1(n730), .A2(n513), .ZN(n741) );
  NAND2_X1 U820 ( .A1(n741), .A2(G286), .ZN(n735) );
  NOR2_X1 U821 ( .A1(G1971), .A2(n770), .ZN(n732) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n718), .ZN(n731) );
  NOR2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U824 ( .A1(n733), .A2(G303), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n737) );
  XNOR2_X1 U826 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n738), .A2(G8), .ZN(n739) );
  NAND2_X1 U828 ( .A1(G8), .A2(n740), .ZN(n745) );
  INV_X1 U829 ( .A(n741), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n763) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n966) );
  AND2_X1 U833 ( .A1(n763), .A2(n966), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n762), .A2(n746), .ZN(n750) );
  INV_X1 U835 ( .A(n966), .ZN(n748) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U838 ( .A1(n756), .A2(n747), .ZN(n978) );
  OR2_X1 U839 ( .A1(n748), .A2(n978), .ZN(n749) );
  AND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U841 ( .A(n753), .B(n752), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n755), .A2(n754), .ZN(n761) );
  NAND2_X1 U843 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  NOR2_X1 U844 ( .A1(n757), .A2(n770), .ZN(n759) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n962) );
  INV_X1 U846 ( .A(n962), .ZN(n758) );
  NOR2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n773) );
  NAND2_X1 U849 ( .A1(n763), .A2(n762), .ZN(n766) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n764) );
  NAND2_X1 U851 ( .A1(G8), .A2(n764), .ZN(n765) );
  NAND2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n767), .A2(n770), .ZN(n771) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n768) );
  XOR2_X1 U855 ( .A(n768), .B(KEYINPUT24), .Z(n769) );
  NOR2_X1 U856 ( .A1(n775), .A2(n774), .ZN(n817) );
  XNOR2_X1 U857 ( .A(G2067), .B(KEYINPUT37), .ZN(n776) );
  XNOR2_X1 U858 ( .A(n776), .B(KEYINPUT94), .ZN(n815) );
  NAND2_X1 U859 ( .A1(n886), .A2(G104), .ZN(n778) );
  NAND2_X1 U860 ( .A1(G140), .A2(n622), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U862 ( .A(KEYINPUT34), .B(n779), .ZN(n785) );
  NAND2_X1 U863 ( .A1(G128), .A2(n883), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G116), .A2(n575), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U866 ( .A(KEYINPUT95), .B(n782), .ZN(n783) );
  XNOR2_X1 U867 ( .A(KEYINPUT35), .B(n783), .ZN(n784) );
  NOR2_X1 U868 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U869 ( .A(KEYINPUT36), .B(n786), .ZN(n865) );
  NOR2_X1 U870 ( .A1(n815), .A2(n865), .ZN(n929) );
  NAND2_X1 U871 ( .A1(n817), .A2(n929), .ZN(n813) );
  NAND2_X1 U872 ( .A1(G107), .A2(n575), .ZN(n788) );
  NAND2_X1 U873 ( .A1(G131), .A2(n622), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U875 ( .A1(G119), .A2(n883), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G95), .A2(n886), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  OR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n892) );
  AND2_X1 U879 ( .A1(n892), .A2(G1991), .ZN(n802) );
  NAND2_X1 U880 ( .A1(G129), .A2(n883), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G141), .A2(n622), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n800) );
  NAND2_X1 U883 ( .A1(G105), .A2(n886), .ZN(n795) );
  XNOR2_X1 U884 ( .A(n795), .B(KEYINPUT38), .ZN(n796) );
  XNOR2_X1 U885 ( .A(n796), .B(KEYINPUT96), .ZN(n798) );
  NAND2_X1 U886 ( .A1(G117), .A2(n575), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n864) );
  INV_X1 U889 ( .A(G1996), .ZN(n844) );
  NOR2_X1 U890 ( .A1(n864), .A2(n844), .ZN(n801) );
  NOR2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n927) );
  XOR2_X1 U892 ( .A(G1986), .B(G290), .Z(n969) );
  NAND2_X1 U893 ( .A1(n927), .A2(n969), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n803), .A2(n817), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n805), .A2(n515), .ZN(n820) );
  AND2_X1 U896 ( .A1(n844), .A2(n864), .ZN(n919) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n892), .ZN(n806) );
  XOR2_X1 U898 ( .A(KEYINPUT105), .B(n806), .Z(n925) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n807) );
  XNOR2_X1 U900 ( .A(KEYINPUT104), .B(n807), .ZN(n808) );
  NOR2_X1 U901 ( .A1(n925), .A2(n808), .ZN(n810) );
  INV_X1 U902 ( .A(n927), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U904 ( .A1(n919), .A2(n811), .ZN(n812) );
  XNOR2_X1 U905 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U907 ( .A1(n815), .A2(n865), .ZN(n922) );
  NAND2_X1 U908 ( .A1(n816), .A2(n922), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U911 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n917), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(G188) );
  XOR2_X1 U917 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  NOR2_X1 U918 ( .A1(n826), .A2(n825), .ZN(G325) );
  XNOR2_X1 U919 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  NOR2_X1 U921 ( .A1(G860), .A2(n827), .ZN(n830) );
  XOR2_X1 U922 ( .A(n828), .B(KEYINPUT82), .Z(n829) );
  XNOR2_X1 U923 ( .A(n830), .B(n829), .ZN(G145) );
  INV_X1 U924 ( .A(G132), .ZN(G219) );
  INV_X1 U925 ( .A(G108), .ZN(G238) );
  INV_X1 U926 ( .A(G82), .ZN(G220) );
  XOR2_X1 U927 ( .A(G2096), .B(G2678), .Z(n832) );
  XNOR2_X1 U928 ( .A(G2072), .B(KEYINPUT43), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U930 ( .A(n833), .B(KEYINPUT42), .Z(n835) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2090), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n840) );
  XNOR2_X1 U933 ( .A(KEYINPUT110), .B(n836), .ZN(n838) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2084), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U937 ( .A(G1976), .B(G1971), .Z(n842) );
  XOR2_X1 U938 ( .A(G1986), .B(n987), .Z(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U940 ( .A(n843), .B(G2474), .Z(n846) );
  XOR2_X1 U941 ( .A(n844), .B(G1991), .Z(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(G1981), .Z(n848) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1956), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(G229) );
  XOR2_X1 U947 ( .A(n851), .B(G286), .Z(n853) );
  XOR2_X1 U948 ( .A(G171), .B(n970), .Z(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U950 ( .A(n854), .B(n980), .Z(n855) );
  NOR2_X1 U951 ( .A1(G37), .A2(n855), .ZN(G397) );
  NAND2_X1 U952 ( .A1(G124), .A2(n883), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n856), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U954 ( .A1(G100), .A2(n886), .ZN(n857) );
  XOR2_X1 U955 ( .A(KEYINPUT111), .B(n857), .Z(n858) );
  NAND2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U957 ( .A1(G112), .A2(n575), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G136), .A2(n622), .ZN(n860) );
  NAND2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U960 ( .A1(n863), .A2(n862), .ZN(G162) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n867) );
  XNOR2_X1 U962 ( .A(G164), .B(G160), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U964 ( .A(KEYINPUT115), .B(KEYINPUT112), .Z(n869) );
  XNOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U967 ( .A(n871), .B(n870), .Z(n882) );
  NAND2_X1 U968 ( .A1(G139), .A2(n622), .ZN(n872) );
  XNOR2_X1 U969 ( .A(KEYINPUT113), .B(n872), .ZN(n880) );
  NAND2_X1 U970 ( .A1(G127), .A2(n883), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G115), .A2(n575), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n875), .B(KEYINPUT47), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT114), .ZN(n878) );
  NAND2_X1 U975 ( .A1(n886), .A2(G103), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n930) );
  XNOR2_X1 U978 ( .A(n930), .B(n924), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n896) );
  NAND2_X1 U980 ( .A1(G130), .A2(n883), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G118), .A2(n575), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U983 ( .A1(n886), .A2(G106), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G142), .A2(n622), .ZN(n887) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U986 ( .A(n889), .B(KEYINPUT45), .Z(n890) );
  NOR2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(G162), .B(n894), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U991 ( .A1(G37), .A2(n897), .ZN(n898) );
  XNOR2_X1 U992 ( .A(KEYINPUT116), .B(n898), .ZN(G395) );
  XNOR2_X1 U993 ( .A(G2446), .B(G2443), .ZN(n908) );
  XOR2_X1 U994 ( .A(G2430), .B(KEYINPUT107), .Z(n900) );
  XNOR2_X1 U995 ( .A(G2454), .B(G2435), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U997 ( .A(G2438), .B(G2427), .Z(n902) );
  XNOR2_X1 U998 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1001 ( .A(KEYINPUT106), .B(G2451), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n909), .A2(G14), .ZN(n916) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n916), .ZN(n913) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n910) );
  XOR2_X1 U1007 ( .A(KEYINPUT49), .B(n910), .Z(n911) );
  XNOR2_X1 U1008 ( .A(n911), .B(KEYINPUT117), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G397), .A2(G395), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  INV_X1 U1015 ( .A(n916), .ZN(G401) );
  INV_X1 U1016 ( .A(n917), .ZN(G223) );
  XOR2_X1 U1017 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1019 ( .A(KEYINPUT51), .B(n920), .Z(n921) );
  XNOR2_X1 U1020 ( .A(n921), .B(KEYINPUT118), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n939) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n937) );
  XOR2_X1 U1025 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1028 ( .A(KEYINPUT50), .B(n933), .Z(n935) );
  XOR2_X1 U1029 ( .A(G160), .B(G2084), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n940), .ZN(n941) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n1019) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n1019), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n942), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1037 ( .A(G2090), .B(G35), .ZN(n955) );
  XOR2_X1 U1038 ( .A(G25), .B(G1991), .Z(n943) );
  NAND2_X1 U1039 ( .A1(n943), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1040 ( .A(G2067), .B(G26), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n950) );
  XOR2_X1 U1043 ( .A(n946), .B(G27), .Z(n948) );
  XNOR2_X1 U1044 ( .A(G1996), .B(G32), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n953), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1050 ( .A(G2084), .B(G34), .Z(n956) );
  XNOR2_X1 U1051 ( .A(KEYINPUT54), .B(n956), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n1020) );
  NOR2_X1 U1053 ( .A1(G29), .A2(KEYINPUT55), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n1020), .A2(n959), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(G11), .A2(n960), .ZN(n1024) );
  XNOR2_X1 U1056 ( .A(KEYINPUT56), .B(KEYINPUT119), .ZN(n961) );
  XOR2_X1 U1057 ( .A(G16), .B(n961), .Z(n986) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(KEYINPUT57), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT120), .B(n965), .ZN(n984) );
  XOR2_X1 U1062 ( .A(G299), .B(G1956), .Z(n967) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n976) );
  XOR2_X1 U1064 ( .A(G171), .B(n987), .Z(n974) );
  NAND2_X1 U1065 ( .A1(G1971), .A2(G303), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1067 ( .A(G1348), .B(n970), .Z(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT121), .B(n979), .Z(n982) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n980), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n1017) );
  INV_X1 U1077 ( .A(G16), .ZN(n1015) );
  XOR2_X1 U1078 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n1013) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G21), .ZN(n989) );
  XOR2_X1 U1080 ( .A(n987), .B(G5), .Z(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n1011) );
  XOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .Z(n990) );
  XNOR2_X1 U1083 ( .A(G4), .B(n990), .ZN(n999) );
  XOR2_X1 U1084 ( .A(G1981), .B(G6), .Z(n994) );
  XNOR2_X1 U1085 ( .A(G20), .B(n991), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(n992), .B(KEYINPUT122), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(G19), .B(G1341), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(n997), .B(KEYINPUT123), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1092 ( .A(KEYINPUT60), .B(n1000), .Z(n1009) );
  XOR2_X1 U1093 ( .A(G1971), .B(G22), .Z(n1003) );
  XOR2_X1 U1094 ( .A(G23), .B(KEYINPUT124), .Z(n1001) );
  XNOR2_X1 U1095 ( .A(n1001), .B(G1976), .ZN(n1002) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1097 ( .A(KEYINPUT125), .B(G1986), .Z(n1004) );
  XNOR2_X1 U1098 ( .A(G24), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1007), .Z(n1008) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(n1013), .B(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(n1018), .B(KEYINPUT127), .ZN(n1022) );
  OR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1027), .ZN(G150) );
  INV_X1 U1112 ( .A(G150), .ZN(G311) );
endmodule

