

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  XOR2_X1 U323 ( .A(n320), .B(n319), .Z(n291) );
  XOR2_X1 U324 ( .A(KEYINPUT65), .B(n379), .Z(n292) );
  XNOR2_X1 U325 ( .A(n315), .B(KEYINPUT78), .ZN(n316) );
  XNOR2_X1 U326 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U327 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n384) );
  XNOR2_X1 U328 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U329 ( .A(n328), .B(n327), .ZN(n376) );
  NOR2_X1 U330 ( .A1(n568), .A2(n572), .ZN(n570) );
  NOR2_X1 U331 ( .A1(n550), .A2(n568), .ZN(n545) );
  XNOR2_X1 U332 ( .A(n457), .B(KEYINPUT58), .ZN(n458) );
  XNOR2_X1 U333 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G36GAT), .B(G190GAT), .Z(n396) );
  XOR2_X1 U335 ( .A(KEYINPUT81), .B(n396), .Z(n296) );
  XOR2_X1 U336 ( .A(G162GAT), .B(KEYINPUT80), .Z(n294) );
  XNOR2_X1 U337 ( .A(G50GAT), .B(G218GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n429) );
  XNOR2_X1 U339 ( .A(G134GAT), .B(n429), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n306) );
  INV_X1 U341 ( .A(G85GAT), .ZN(n297) );
  NAND2_X1 U342 ( .A1(G92GAT), .A2(n297), .ZN(n300) );
  INV_X1 U343 ( .A(G92GAT), .ZN(n298) );
  NAND2_X1 U344 ( .A1(n298), .A2(G85GAT), .ZN(n299) );
  NAND2_X1 U345 ( .A1(n300), .A2(n299), .ZN(n302) );
  XNOR2_X1 U346 ( .A(G99GAT), .B(G106GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n317) );
  XOR2_X1 U348 ( .A(n317), .B(KEYINPUT82), .Z(n304) );
  NAND2_X1 U349 ( .A1(G232GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n306), .B(n305), .Z(n314) );
  XOR2_X1 U352 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n308) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(G29GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT70), .B(n309), .Z(n345) );
  XOR2_X1 U356 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n311) );
  XNOR2_X1 U357 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n345), .B(n312), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n563) );
  XNOR2_X1 U361 ( .A(n563), .B(KEYINPUT83), .ZN(n551) );
  AND2_X1 U362 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XOR2_X1 U363 ( .A(KEYINPUT32), .B(n318), .Z(n320) );
  XOR2_X1 U364 ( .A(G57GAT), .B(KEYINPUT13), .Z(n364) );
  XNOR2_X1 U365 ( .A(n364), .B(KEYINPUT31), .ZN(n319) );
  XOR2_X1 U366 ( .A(KEYINPUT76), .B(G64GAT), .Z(n322) );
  XNOR2_X1 U367 ( .A(G176GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n322), .B(n321), .ZN(n388) );
  XNOR2_X1 U369 ( .A(n291), .B(n388), .ZN(n328) );
  XOR2_X1 U370 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n324) );
  XNOR2_X1 U371 ( .A(KEYINPUT74), .B(KEYINPUT77), .ZN(n323) );
  XOR2_X1 U372 ( .A(n324), .B(n323), .Z(n326) );
  XOR2_X1 U373 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XOR2_X1 U374 ( .A(G148GAT), .B(G78GAT), .Z(n424) );
  XNOR2_X1 U375 ( .A(n442), .B(n424), .ZN(n325) );
  NAND2_X1 U376 ( .A1(n376), .A2(KEYINPUT41), .ZN(n330) );
  OR2_X1 U377 ( .A1(n376), .A2(KEYINPUT41), .ZN(n329) );
  NAND2_X1 U378 ( .A1(n330), .A2(n329), .ZN(n507) );
  XOR2_X1 U379 ( .A(G8GAT), .B(G197GAT), .Z(n332) );
  XNOR2_X1 U380 ( .A(G50GAT), .B(G36GAT), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U382 ( .A(n333), .B(G113GAT), .Z(n335) );
  XOR2_X1 U383 ( .A(G141GAT), .B(G22GAT), .Z(n425) );
  XNOR2_X1 U384 ( .A(G169GAT), .B(n425), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n341) );
  XOR2_X1 U386 ( .A(G1GAT), .B(KEYINPUT71), .Z(n337) );
  XNOR2_X1 U387 ( .A(G15GAT), .B(KEYINPUT72), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n366) );
  XOR2_X1 U389 ( .A(n366), .B(KEYINPUT29), .Z(n339) );
  NAND2_X1 U390 ( .A1(G229GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U392 ( .A(n341), .B(n340), .Z(n347) );
  XOR2_X1 U393 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n343) );
  XNOR2_X1 U394 ( .A(KEYINPUT73), .B(KEYINPUT69), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U397 ( .A(n347), .B(n346), .ZN(n578) );
  NOR2_X1 U398 ( .A1(n507), .A2(n578), .ZN(n350) );
  XOR2_X1 U399 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n348) );
  XNOR2_X1 U400 ( .A(KEYINPUT114), .B(n348), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n371) );
  XOR2_X1 U402 ( .A(KEYINPUT87), .B(KEYINPUT12), .Z(n352) );
  XNOR2_X1 U403 ( .A(KEYINPUT14), .B(KEYINPUT84), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n370) );
  XOR2_X1 U405 ( .A(G211GAT), .B(G155GAT), .Z(n354) );
  XNOR2_X1 U406 ( .A(G71GAT), .B(G127GAT), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U408 ( .A(KEYINPUT15), .B(KEYINPUT88), .Z(n356) );
  XNOR2_X1 U409 ( .A(G22GAT), .B(G78GAT), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U411 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U412 ( .A(KEYINPUT85), .B(G64GAT), .Z(n360) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U415 ( .A(KEYINPUT86), .B(n361), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U417 ( .A(n365), .B(n364), .Z(n368) );
  XOR2_X1 U418 ( .A(G8GAT), .B(G183GAT), .Z(n389) );
  XNOR2_X1 U419 ( .A(n366), .B(n389), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U421 ( .A(n370), .B(n369), .Z(n489) );
  NOR2_X1 U422 ( .A1(n371), .A2(n489), .ZN(n373) );
  INV_X1 U423 ( .A(KEYINPUT116), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n373), .B(n372), .ZN(n374) );
  NOR2_X1 U425 ( .A1(n563), .A2(n374), .ZN(n375) );
  XNOR2_X1 U426 ( .A(n375), .B(KEYINPUT47), .ZN(n383) );
  INV_X1 U427 ( .A(n376), .ZN(n582) );
  NAND2_X1 U428 ( .A1(n578), .A2(n582), .ZN(n380) );
  XNOR2_X1 U429 ( .A(KEYINPUT36), .B(n551), .ZN(n588) );
  INV_X1 U430 ( .A(n489), .ZN(n585) );
  NOR2_X1 U431 ( .A1(n588), .A2(n585), .ZN(n378) );
  XNOR2_X1 U432 ( .A(KEYINPUT117), .B(KEYINPUT45), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n379) );
  NOR2_X1 U434 ( .A1(n380), .A2(n292), .ZN(n381) );
  XOR2_X1 U435 ( .A(KEYINPUT118), .B(n381), .Z(n382) );
  AND2_X1 U436 ( .A1(n383), .A2(n382), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n533) );
  XOR2_X1 U438 ( .A(G211GAT), .B(KEYINPUT93), .Z(n387) );
  XNOR2_X1 U439 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n428) );
  XNOR2_X1 U441 ( .A(n428), .B(n388), .ZN(n400) );
  XOR2_X1 U442 ( .A(n389), .B(G92GAT), .Z(n394) );
  XOR2_X1 U443 ( .A(KEYINPUT90), .B(KEYINPUT17), .Z(n391) );
  XNOR2_X1 U444 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U446 ( .A(G169GAT), .B(n392), .Z(n453) );
  XNOR2_X1 U447 ( .A(n453), .B(G218GAT), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U449 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U452 ( .A(n400), .B(n399), .ZN(n465) );
  NOR2_X1 U453 ( .A1(n533), .A2(n465), .ZN(n401) );
  XNOR2_X1 U454 ( .A(n401), .B(KEYINPUT54), .ZN(n575) );
  XOR2_X1 U455 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n403) );
  XNOR2_X1 U456 ( .A(KEYINPUT94), .B(G155GAT), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U458 ( .A(KEYINPUT95), .B(n404), .Z(n439) );
  XOR2_X1 U459 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n406) );
  NAND2_X1 U460 ( .A1(G225GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U462 ( .A(KEYINPUT5), .B(n407), .ZN(n422) );
  XOR2_X1 U463 ( .A(G57GAT), .B(G148GAT), .Z(n409) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(G141GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U466 ( .A(KEYINPUT4), .B(KEYINPUT96), .Z(n411) );
  XNOR2_X1 U467 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U469 ( .A(n413), .B(n412), .Z(n420) );
  XOR2_X1 U470 ( .A(G85GAT), .B(G162GAT), .Z(n417) );
  XOR2_X1 U471 ( .A(G127GAT), .B(KEYINPUT0), .Z(n415) );
  XNOR2_X1 U472 ( .A(G113GAT), .B(G134GAT), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n443) );
  XNOR2_X1 U474 ( .A(G120GAT), .B(n443), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U476 ( .A(G29GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n439), .B(n423), .ZN(n521) );
  INV_X1 U480 ( .A(n521), .ZN(n574) );
  XOR2_X1 U481 ( .A(KEYINPUT22), .B(G106GAT), .Z(n427) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n435) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n431) );
  XNOR2_X1 U486 ( .A(G204GAT), .B(KEYINPUT92), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n469) );
  AND2_X1 U493 ( .A1(n574), .A2(n469), .ZN(n440) );
  NAND2_X1 U494 ( .A1(n575), .A2(n440), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n441), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U496 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U499 ( .A(G183GAT), .B(KEYINPUT20), .Z(n447) );
  XNOR2_X1 U500 ( .A(G176GAT), .B(KEYINPUT91), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U502 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U503 ( .A(G190GAT), .B(G99GAT), .Z(n451) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G15GAT), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n536) );
  NAND2_X1 U508 ( .A1(n456), .A2(n536), .ZN(n572) );
  NOR2_X1 U509 ( .A1(n551), .A2(n572), .ZN(n459) );
  INV_X1 U510 ( .A(G190GAT), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n480) );
  NOR2_X1 U512 ( .A1(n376), .A2(n578), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n460), .B(KEYINPUT79), .ZN(n494) );
  NAND2_X1 U514 ( .A1(n551), .A2(n489), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n461), .B(KEYINPUT89), .ZN(n462) );
  XNOR2_X1 U516 ( .A(KEYINPUT16), .B(n462), .ZN(n478) );
  XOR2_X1 U517 ( .A(KEYINPUT67), .B(KEYINPUT28), .Z(n463) );
  XNOR2_X1 U518 ( .A(n469), .B(n463), .ZN(n539) );
  XOR2_X1 U519 ( .A(n465), .B(KEYINPUT27), .Z(n471) );
  NAND2_X1 U520 ( .A1(n471), .A2(n521), .ZN(n532) );
  NOR2_X1 U521 ( .A1(n536), .A2(n532), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n539), .A2(n464), .ZN(n476) );
  INV_X1 U523 ( .A(n465), .ZN(n523) );
  NAND2_X1 U524 ( .A1(n523), .A2(n536), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n466), .A2(n469), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT25), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT99), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n469), .A2(n536), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT26), .ZN(n576) );
  NAND2_X1 U530 ( .A1(n471), .A2(n576), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n574), .A2(n474), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U534 ( .A(KEYINPUT100), .B(n477), .ZN(n491) );
  NAND2_X1 U535 ( .A1(n478), .A2(n491), .ZN(n509) );
  NOR2_X1 U536 ( .A1(n494), .A2(n509), .ZN(n486) );
  NAND2_X1 U537 ( .A1(n486), .A2(n521), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NAND2_X1 U540 ( .A1(n523), .A2(n486), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT102), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U544 ( .A1(n486), .A2(n536), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  XOR2_X1 U546 ( .A(G22GAT), .B(KEYINPUT103), .Z(n488) );
  INV_X1 U547 ( .A(n539), .ZN(n529) );
  NAND2_X1 U548 ( .A1(n486), .A2(n529), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n497) );
  NOR2_X1 U551 ( .A1(n489), .A2(n588), .ZN(n490) );
  NAND2_X1 U552 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n492), .ZN(n493) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(n493), .Z(n520) );
  NOR2_X1 U555 ( .A1(n520), .A2(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(KEYINPUT38), .B(n495), .ZN(n504) );
  NAND2_X1 U557 ( .A1(n504), .A2(n521), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U559 ( .A(G29GAT), .B(n498), .Z(G1328GAT) );
  NAND2_X1 U560 ( .A1(n504), .A2(n523), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(KEYINPUT106), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n502) );
  NAND2_X1 U564 ( .A1(n536), .A2(n504), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(KEYINPUT108), .ZN(n506) );
  NAND2_X1 U568 ( .A1(n529), .A2(n504), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n511) );
  XNOR2_X1 U571 ( .A(KEYINPUT110), .B(n507), .ZN(n568) );
  INV_X1 U572 ( .A(n568), .ZN(n508) );
  NAND2_X1 U573 ( .A1(n578), .A2(n508), .ZN(n519) );
  NOR2_X1 U574 ( .A1(n519), .A2(n509), .ZN(n516) );
  NAND2_X1 U575 ( .A1(n516), .A2(n521), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  XOR2_X1 U578 ( .A(G64GAT), .B(KEYINPUT111), .Z(n514) );
  NAND2_X1 U579 ( .A1(n516), .A2(n523), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n536), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U584 ( .A1(n516), .A2(n529), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NOR2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n521), .A2(n528), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n525) );
  NAND2_X1 U590 ( .A1(n528), .A2(n523), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n528), .A2(n536), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  INV_X1 U598 ( .A(KEYINPUT120), .ZN(n538) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n535) );
  INV_X1 U600 ( .A(KEYINPUT119), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n554) );
  NAND2_X1 U602 ( .A1(n554), .A2(n536), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n540) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n550) );
  NOR2_X1 U605 ( .A1(n550), .A2(n578), .ZN(n542) );
  XNOR2_X1 U606 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n543), .B(G113GAT), .ZN(G1340GAT) );
  XNOR2_X1 U609 ( .A(KEYINPUT123), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U611 ( .A(n546), .B(G120GAT), .Z(G1341GAT) );
  INV_X1 U612 ( .A(KEYINPUT50), .ZN(n548) );
  NOR2_X1 U613 ( .A1(n550), .A2(n585), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(G127GAT), .ZN(G1342GAT) );
  NOR2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n576), .ZN(n562) );
  NOR2_X1 U620 ( .A1(n578), .A2(n562), .ZN(n555) );
  XOR2_X1 U621 ( .A(G141GAT), .B(n555), .Z(G1344GAT) );
  NOR2_X1 U622 ( .A1(n507), .A2(n562), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT125), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(KEYINPUT124), .B(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NOR2_X1 U628 ( .A1(n585), .A2(n562), .ZN(n561) );
  XOR2_X1 U629 ( .A(G155GAT), .B(n561), .Z(G1346GAT) );
  INV_X1 U630 ( .A(n562), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT126), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  NOR2_X1 U634 ( .A1(n578), .A2(n572), .ZN(n567) );
  XOR2_X1 U635 ( .A(G169GAT), .B(n567), .Z(G1348GAT) );
  XNOR2_X1 U636 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(n571), .ZN(G1349GAT) );
  NOR2_X1 U639 ( .A1(n585), .A2(n572), .ZN(n573) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n573), .Z(G1350GAT) );
  AND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n587) );
  NOR2_X1 U643 ( .A1(n578), .A2(n587), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n587), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

