//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G101), .ZN(new_n189));
  INV_X1    g003(.A(G210), .ZN(new_n190));
  NOR3_X1   g004(.A1(new_n190), .A2(G237), .A3(G953), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT64), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n196), .B1(new_n201), .B2(new_n195), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n195), .A2(G143), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT67), .B1(new_n202), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n197), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  OAI21_X1  g022(.A(G128), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n210));
  AOI21_X1  g024(.A(G146), .B1(new_n198), .B2(new_n200), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n209), .B(new_n210), .C1(new_n211), .C2(new_n196), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(G143), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n207), .B1(new_n213), .B2(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT66), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n198), .A2(new_n200), .A3(G146), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n217), .A2(KEYINPUT66), .A3(new_n204), .A4(new_n215), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n206), .B(new_n212), .C1(new_n216), .C2(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT65), .A2(G137), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT65), .A2(G137), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n221), .A2(KEYINPUT11), .A3(G134), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT11), .B1(new_n224), .B2(G134), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(G134), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n221), .A2(new_n222), .ZN(new_n231));
  INV_X1    g045(.A(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n228), .B1(new_n233), .B2(new_n226), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n220), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n228), .B1(new_n223), .B2(new_n227), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n229), .ZN(new_n239));
  INV_X1    g053(.A(new_n196), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n213), .B2(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n241), .A2(new_n245), .B1(new_n214), .B2(new_n243), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n236), .A2(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n248), .A2(KEYINPUT74), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT68), .A2(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT68), .A2(G119), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(G116), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G116), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G119), .ZN(new_n255));
  INV_X1    g069(.A(G113), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT2), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G113), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n255), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n253), .B2(new_n255), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n250), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n253), .A2(new_n255), .ZN(new_n265));
  INV_X1    g079(.A(new_n260), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n261), .A3(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n248), .B2(KEYINPUT74), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT28), .B1(new_n249), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n236), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n220), .A2(KEYINPUT71), .A3(new_n235), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n230), .A2(new_n237), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n241), .A2(new_n245), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n214), .A2(new_n243), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT70), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n239), .A2(new_n246), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n275), .A2(new_n269), .A3(new_n276), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n248), .A2(new_n270), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n273), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n188), .B(new_n194), .C1(new_n272), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n194), .B1(new_n272), .B2(new_n287), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT75), .ZN(new_n290));
  INV_X1    g104(.A(new_n194), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT30), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n236), .A2(new_n294), .A3(new_n247), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n275), .A2(new_n276), .A3(new_n284), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(KEYINPUT30), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n293), .B1(new_n297), .B2(new_n269), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n236), .A2(new_n274), .B1(new_n281), .B2(new_n283), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n294), .B1(new_n299), .B2(new_n276), .ZN(new_n300));
  OAI211_X1 g114(.A(KEYINPUT72), .B(new_n270), .C1(new_n300), .C2(new_n295), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n292), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n288), .B(new_n290), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AOI211_X1 g118(.A(KEYINPUT31), .B(new_n292), .C1(new_n298), .C2(new_n301), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n187), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT76), .B(KEYINPUT32), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(KEYINPUT32), .B(new_n187), .C1(new_n304), .C2(new_n305), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n249), .A2(new_n271), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n273), .ZN(new_n312));
  INV_X1    g126(.A(new_n287), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n291), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n296), .A2(KEYINPUT30), .ZN(new_n317));
  INV_X1    g131(.A(new_n295), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT72), .B1(new_n319), .B2(new_n270), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n297), .A2(new_n293), .A3(new_n269), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n285), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n316), .B1(new_n322), .B2(new_n194), .ZN(new_n323));
  INV_X1    g137(.A(G902), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n296), .A2(new_n270), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n325), .A2(new_n285), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n312), .B1(new_n326), .B2(new_n273), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n291), .A2(KEYINPUT29), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G472), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n309), .A2(new_n310), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G214), .B1(G237), .B2(G902), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n334));
  INV_X1    g148(.A(G107), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G104), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g151(.A(G101), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n334), .A2(new_n339), .A3(new_n335), .A4(G104), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n335), .A2(G104), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n337), .A2(new_n338), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G104), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(G107), .ZN(new_n345));
  OAI21_X1  g159(.A(G101), .B1(new_n345), .B2(new_n341), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n251), .A2(new_n349), .A3(G116), .A4(new_n252), .ZN(new_n350));
  OAI211_X1 g164(.A(G113), .B(new_n350), .C1(new_n265), .C2(new_n349), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n261), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n341), .B1(new_n336), .B2(KEYINPUT3), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n340), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G101), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n343), .A2(KEYINPUT4), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n338), .B1(new_n353), .B2(new_n340), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n352), .B1(new_n269), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G110), .B(G122), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n352), .B(new_n361), .C1(new_n269), .C2(new_n359), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n217), .A2(new_n204), .A3(new_n215), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT66), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n218), .ZN(new_n369));
  INV_X1    g183(.A(G125), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n206), .A4(new_n212), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n280), .A2(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G953), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(G224), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(G224), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n371), .A2(new_n376), .A3(new_n372), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n360), .A2(new_n379), .A3(new_n362), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n365), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n361), .B(KEYINPUT8), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n253), .A2(KEYINPUT5), .A3(new_n255), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n350), .A2(G113), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n261), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(new_n347), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n351), .A2(new_n261), .B1(new_n343), .B2(new_n346), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n376), .A2(KEYINPUT7), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n371), .A2(new_n372), .A3(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n364), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n371), .A2(KEYINPUT85), .ZN(new_n393));
  INV_X1    g207(.A(new_n212), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n210), .B1(new_n241), .B2(new_n209), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n370), .A4(new_n369), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n393), .A2(new_n398), .A3(new_n372), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n389), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT86), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n392), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n246), .A2(new_n370), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n371), .B2(KEYINPUT85), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n390), .B1(new_n404), .B2(new_n398), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(KEYINPUT86), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n324), .B(new_n381), .C1(new_n402), .C2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G210), .B1(G237), .B2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n364), .A2(new_n388), .A3(new_n391), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n405), .B2(KEYINPUT86), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n400), .A2(new_n401), .ZN(new_n413));
  AOI21_X1  g227(.A(G902), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n408), .A3(new_n381), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n333), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT87), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G140), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n374), .A2(G227), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT80), .ZN(new_n421));
  AND4_X1   g235(.A1(new_n369), .A2(new_n206), .A3(new_n212), .A4(new_n347), .ZN(new_n422));
  INV_X1    g236(.A(new_n214), .ZN(new_n423));
  OAI21_X1  g237(.A(G128), .B1(new_n211), .B2(new_n208), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n347), .B1(new_n369), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(KEYINPUT12), .B(new_n239), .C1(new_n422), .C2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n396), .A2(new_n369), .A3(new_n347), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n369), .A2(new_n425), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n348), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(KEYINPUT82), .A3(KEYINPUT12), .A4(new_n239), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n239), .B1(new_n422), .B2(new_n426), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT12), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n429), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n426), .A2(KEYINPUT10), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n359), .A2(new_n280), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n348), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n277), .A4(new_n441), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n438), .A2(KEYINPUT83), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT83), .B1(new_n438), .B2(new_n442), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n421), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n420), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n239), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n445), .A2(G469), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n442), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n420), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n438), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n429), .A2(new_n434), .A3(new_n437), .A4(KEYINPUT84), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n447), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n453), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G469), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n324), .ZN(new_n460));
  NAND2_X1  g274(.A1(G469), .A2(G902), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n451), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT9), .B(G234), .ZN(new_n463));
  OAI21_X1  g277(.A(G221), .B1(new_n463), .B2(G902), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n464), .B(KEYINPUT79), .Z(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n417), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G217), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(G234), .B2(new_n324), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G140), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G125), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n370), .A2(G140), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT16), .ZN(new_n475));
  OR3_X1    g289(.A1(new_n370), .A2(KEYINPUT16), .A3(G140), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(G146), .ZN(new_n477));
  XNOR2_X1  g291(.A(G125), .B(G140), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n195), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n251), .A2(new_n252), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n203), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n482), .A2(KEYINPUT77), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n251), .A2(G128), .A3(new_n252), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT23), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(KEYINPUT77), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G110), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G119), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n484), .B1(new_n491), .B2(G128), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT24), .B(G110), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n480), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n488), .B1(new_n487), .B2(new_n489), .ZN(new_n496));
  INV_X1    g310(.A(new_n477), .ZN(new_n497));
  AOI21_X1  g311(.A(G146), .B1(new_n475), .B2(new_n476), .ZN(new_n498));
  OAI22_X1  g312(.A1(new_n497), .A2(new_n498), .B1(new_n492), .B2(new_n493), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT22), .B(G137), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n374), .A2(G221), .A3(G234), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n495), .B2(new_n500), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n324), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT25), .A4(new_n324), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n471), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n470), .A2(G902), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n505), .A2(new_n507), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT78), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n254), .A2(G122), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n254), .A2(G122), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G107), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n335), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n213), .A2(G128), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n197), .A2(G128), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n232), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n201), .A2(new_n203), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(new_n524), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT94), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n523), .B(new_n532), .C1(new_n524), .C2(new_n529), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT95), .B1(new_n523), .B2(new_n529), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n535));
  INV_X1    g349(.A(new_n529), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n528), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n531), .A2(new_n533), .A3(new_n534), .A4(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n527), .B1(new_n538), .B2(G134), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G134), .B1(new_n528), .B2(new_n524), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n541), .A2(new_n526), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n519), .A2(KEYINPUT14), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT14), .ZN(new_n544));
  OAI21_X1  g358(.A(G107), .B1(new_n518), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n521), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n463), .A2(new_n469), .A3(G953), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n540), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n549), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n539), .B2(new_n547), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT96), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n324), .ZN(new_n555));
  INV_X1    g369(.A(G478), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n557), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(KEYINPUT18), .A2(G131), .ZN(new_n561));
  INV_X1    g375(.A(G237), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n374), .A3(G214), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n563), .A2(new_n197), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n213), .A2(new_n563), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT89), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n561), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n561), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT89), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n473), .A2(new_n474), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G146), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n573), .A2(new_n479), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT88), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n574), .A2(KEYINPUT88), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT19), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n478), .A2(KEYINPUT19), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(KEYINPUT90), .B(new_n477), .C1(new_n581), .C2(G146), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT90), .ZN(new_n583));
  AOI21_X1  g397(.A(G146), .B1(new_n579), .B2(new_n580), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(new_n497), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n566), .A2(G131), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n564), .A2(new_n565), .A3(new_n228), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n582), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n577), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(G113), .B(G122), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n344), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n586), .A2(new_n595), .A3(new_n587), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n228), .B1(new_n564), .B2(new_n565), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n596), .A2(new_n597), .B1(KEYINPUT17), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n497), .B2(new_n498), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(new_n597), .A3(KEYINPUT17), .ZN(new_n602));
  INV_X1    g416(.A(new_n498), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(KEYINPUT91), .A3(new_n477), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n592), .B(new_n577), .C1(new_n599), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n594), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT20), .ZN(new_n608));
  NOR2_X1   g422(.A1(G475), .A2(G902), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n608), .B1(new_n607), .B2(new_n609), .ZN(new_n611));
  INV_X1    g425(.A(G475), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n577), .B1(new_n599), .B2(new_n605), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n593), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n614), .B2(new_n606), .ZN(new_n615));
  OAI22_X1  g429(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(G234), .A2(G237), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n617), .A2(G952), .A3(new_n374), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT21), .B(G898), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT97), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n617), .A2(G902), .A3(G953), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n560), .A2(new_n616), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n624), .A2(KEYINPUT98), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(KEYINPUT98), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n331), .A2(new_n468), .A3(new_n516), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  OAI21_X1  g443(.A(new_n324), .B1(new_n304), .B2(new_n305), .ZN(new_n630));
  INV_X1    g444(.A(new_n292), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n320), .B2(new_n321), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT31), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n302), .A2(new_n303), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n633), .A2(new_n634), .A3(new_n288), .A4(new_n290), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n630), .A2(G472), .B1(new_n635), .B2(new_n187), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n462), .A2(new_n516), .A3(new_n466), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n611), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n614), .A2(new_n606), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n324), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n639), .A2(new_n640), .B1(new_n642), .B2(G475), .ZN(new_n643));
  AOI21_X1  g457(.A(G478), .B1(new_n553), .B2(new_n324), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(KEYINPUT33), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(KEYINPUT33), .ZN(new_n648));
  INV_X1    g462(.A(new_n552), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n539), .A2(new_n547), .A3(new_n551), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n550), .A2(new_n552), .A3(KEYINPUT99), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n556), .A2(G902), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n644), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n643), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n623), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n416), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n638), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  NAND2_X1  g479(.A1(new_n642), .A2(G475), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n639), .A2(new_n640), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n642), .A2(KEYINPUT101), .A3(G475), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n560), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n661), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n638), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT35), .B(G107), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT102), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT103), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n674), .B(new_n677), .ZN(G9));
  NOR2_X1   g492(.A1(new_n506), .A2(KEYINPUT36), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n501), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n513), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n512), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n625), .B2(new_n626), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n468), .A2(new_n685), .A3(new_n636), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  NOR2_X1   g502(.A1(new_n407), .A2(new_n409), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n408), .B1(new_n414), .B2(new_n381), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n332), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT104), .B(G900), .Z(new_n692));
  AOI21_X1  g506(.A(new_n618), .B1(new_n692), .B2(new_n622), .ZN(new_n693));
  NOR4_X1   g507(.A1(new_n672), .A2(new_n691), .A3(new_n684), .A4(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n467), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n330), .A2(new_n310), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n307), .B1(new_n635), .B2(new_n187), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n694), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XOR2_X1   g513(.A(new_n693), .B(KEYINPUT39), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n309), .A2(new_n310), .ZN(new_n703));
  INV_X1    g517(.A(G472), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n326), .A2(new_n194), .ZN(new_n705));
  INV_X1    g519(.A(new_n285), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n298), .B2(new_n301), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n705), .B1(new_n707), .B2(new_n194), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n708), .A2(KEYINPUT106), .ZN(new_n709));
  AOI21_X1  g523(.A(G902), .B1(new_n708), .B2(KEYINPUT106), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n704), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n689), .A2(new_n690), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n684), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n560), .A2(new_n616), .ZN(new_n719));
  NOR4_X1   g533(.A1(new_n717), .A2(new_n333), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n702), .A2(new_n713), .A3(new_n714), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n201), .ZN(G45));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  INV_X1    g537(.A(new_n693), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n556), .B(G902), .C1(new_n651), .C2(new_n653), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n616), .B(new_n724), .C1(new_n725), .C2(new_n644), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n723), .B1(new_n691), .B2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n643), .A2(new_n656), .A3(new_n693), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n416), .A3(KEYINPUT107), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n684), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  NAND2_X1  g546(.A1(new_n458), .A2(new_n324), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G469), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(KEYINPUT108), .A3(new_n460), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n736), .A3(G469), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n465), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n331), .A2(new_n662), .A3(new_n516), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT109), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n739), .B(new_n741), .ZN(G15));
  INV_X1    g556(.A(new_n516), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n672), .A2(new_n743), .A3(new_n623), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n331), .A2(new_n744), .A3(new_n416), .A4(new_n738), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G116), .ZN(G18));
  NAND4_X1  g560(.A1(new_n331), .A2(new_n685), .A3(new_n416), .A4(new_n738), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT110), .B(G119), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G21));
  AOI21_X1  g563(.A(new_n273), .B1(new_n325), .B2(new_n285), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n194), .B1(new_n750), .B2(new_n272), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n302), .B2(new_n303), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT112), .B(new_n751), .C1(new_n302), .C2(new_n303), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n634), .A3(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n187), .B(KEYINPUT111), .Z(new_n757));
  AOI22_X1  g571(.A1(new_n756), .A2(new_n757), .B1(new_n630), .B2(G472), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n661), .A2(new_n719), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n516), .A3(new_n738), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  NOR2_X1   g575(.A1(new_n691), .A2(new_n726), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n758), .A2(new_n718), .A3(new_n738), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  AOI21_X1  g578(.A(KEYINPUT32), .B1(new_n635), .B2(new_n187), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n516), .B1(new_n696), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n715), .A2(new_n332), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n695), .A2(new_n728), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT42), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n467), .A2(new_n767), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n726), .A2(KEYINPUT42), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n331), .A2(new_n771), .A3(new_n516), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n228), .ZN(G33));
  NOR2_X1   g589(.A1(new_n672), .A2(new_n693), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n331), .A2(new_n771), .A3(new_n516), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(new_n636), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n656), .A2(new_n616), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT43), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n718), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n785), .A3(new_n767), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n445), .A2(new_n450), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT45), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(KEYINPUT45), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(G469), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT46), .B1(new_n790), .B2(new_n461), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n790), .A2(new_n461), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n794), .A2(KEYINPUT113), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n460), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n791), .B2(new_n792), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT113), .B1(new_n794), .B2(new_n795), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n793), .A2(new_n796), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n786), .A2(new_n466), .A3(new_n800), .A4(new_n700), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n466), .ZN(new_n803));
  NOR2_X1   g617(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n804));
  NAND2_X1  g618(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n800), .A2(new_n466), .A3(new_n805), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n331), .A2(new_n516), .A3(new_n726), .A4(new_n767), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n781), .A2(new_n618), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n758), .A3(new_n516), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n738), .A2(new_n333), .A3(new_n717), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n712), .A2(new_n516), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n618), .A2(new_n820), .A3(new_n738), .A4(new_n768), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n643), .A3(new_n656), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n816), .A2(new_n817), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n813), .A2(new_n738), .A3(new_n768), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n758), .A2(new_n718), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n818), .A2(new_n822), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n735), .A2(new_n737), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n807), .A2(new_n808), .B1(new_n465), .B2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n814), .A2(new_n767), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n738), .A2(new_n416), .ZN(new_n833));
  OAI211_X1 g647(.A(G952), .B(new_n374), .C1(new_n814), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n659), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(new_n821), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n824), .A2(new_n766), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT48), .Z(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n839), .A2(KEYINPUT119), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(KEYINPUT119), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n831), .A2(new_n832), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n763), .A2(new_n698), .A3(new_n731), .ZN(new_n843));
  INV_X1    g657(.A(new_n719), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n512), .A2(new_n683), .A3(new_n693), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n845), .A3(new_n416), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n467), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n703), .B2(new_n711), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n763), .A2(new_n848), .A3(new_n698), .A4(new_n731), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n467), .A2(new_n684), .A3(new_n767), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n671), .A2(new_n558), .A3(new_n559), .A4(new_n724), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n330), .A2(new_n310), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n309), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n756), .A2(new_n757), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n630), .A2(G472), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n860), .A2(new_n861), .A3(new_n728), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n856), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n770), .A3(new_n773), .A4(new_n777), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n657), .A2(KEYINPUT116), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n643), .B2(new_n656), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n560), .A2(new_n643), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n417), .A3(new_n623), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n636), .A3(new_n637), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n739), .A3(new_n760), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n628), .A2(new_n747), .A3(new_n745), .A4(new_n686), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n864), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n770), .A2(new_n773), .A3(new_n777), .ZN(new_n879));
  INV_X1    g693(.A(new_n874), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n872), .A2(new_n739), .A3(new_n760), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .A4(new_n863), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n850), .B(KEYINPUT52), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n876), .A2(new_n877), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n855), .A2(new_n875), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n878), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n882), .A2(new_n883), .A3(new_n878), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n885), .B1(KEYINPUT54), .B2(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n827), .B(KEYINPUT51), .C1(new_n829), .C2(new_n830), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n842), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(G952), .B2(G953), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n717), .A2(new_n332), .A3(new_n466), .A4(new_n780), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT49), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n828), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n820), .B(new_n896), .C1(new_n895), .C2(new_n828), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n897), .ZN(G75));
  NAND2_X1  g712(.A1(new_n876), .A2(new_n884), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT121), .B1(new_n899), .B2(G902), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n901), .B(new_n324), .C1(new_n876), .C2(new_n884), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n409), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n365), .A2(new_n380), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(new_n378), .Z(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n904), .A2(new_n905), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n324), .B1(new_n876), .B2(new_n884), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(G210), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT120), .B(new_n908), .C1(new_n912), .C2(KEYINPUT56), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT56), .B1(new_n911), .B2(G210), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n909), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n374), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n910), .A2(new_n917), .A3(new_n919), .ZN(G51));
  INV_X1    g734(.A(new_n790), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n461), .B(KEYINPUT57), .Z(new_n922));
  AOI21_X1  g736(.A(new_n877), .B1(new_n876), .B2(new_n884), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n885), .B2(new_n923), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n903), .A2(new_n921), .B1(new_n924), .B2(new_n458), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT122), .B1(new_n925), .B2(new_n918), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n924), .A2(new_n458), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n900), .A2(new_n902), .A3(new_n790), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n927), .B(new_n919), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n926), .A2(new_n930), .ZN(G54));
  AND2_X1   g745(.A1(KEYINPUT58), .A2(G475), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n903), .A2(new_n607), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n607), .B1(new_n903), .B2(new_n932), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n918), .ZN(G60));
  NOR2_X1   g749(.A1(new_n885), .A2(new_n923), .ZN(new_n936));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT59), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n654), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n919), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n653), .B(new_n651), .C1(new_n890), .C2(new_n938), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n941), .A2(new_n942), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT124), .Z(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n876), .B2(new_n884), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n919), .B1(new_n951), .B2(new_n515), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n681), .B2(new_n951), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g768(.A(new_n374), .B1(new_n620), .B2(G224), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n874), .A2(new_n873), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT125), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n957), .B2(new_n374), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n906), .B1(G898), .B2(new_n374), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT126), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G69));
  AOI21_X1  g775(.A(new_n374), .B1(G227), .B2(G900), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n319), .B(new_n581), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(G900), .B2(G953), .ZN(new_n964));
  INV_X1    g778(.A(new_n700), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n844), .A2(new_n416), .ZN(new_n966));
  OR4_X1    g780(.A1(new_n965), .A2(new_n803), .A3(new_n766), .A4(new_n966), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n801), .A2(new_n879), .A3(new_n843), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n810), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n969), .B2(G953), .ZN(new_n970));
  INV_X1    g784(.A(new_n963), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n721), .A2(new_n843), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  NOR3_X1   g787(.A1(new_n701), .A2(new_n767), .A3(new_n870), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n516), .A3(new_n331), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n801), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n810), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n971), .B1(new_n977), .B2(new_n374), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n970), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n962), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n978), .A2(new_n979), .ZN(new_n984));
  INV_X1    g798(.A(new_n962), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n981), .A3(new_n985), .A4(new_n970), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n969), .B2(new_n957), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(new_n194), .A3(new_n707), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n632), .B1(new_n291), .B2(new_n707), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n889), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n989), .B1(new_n977), .B2(new_n957), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n291), .A3(new_n322), .ZN(new_n995));
  AND4_X1   g809(.A1(new_n919), .A2(new_n991), .A3(new_n993), .A4(new_n995), .ZN(G57));
endmodule


