

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U326 ( .A(n384), .B(n344), .ZN(n345) );
  XOR2_X1 U327 ( .A(n333), .B(n332), .Z(n572) );
  XNOR2_X1 U328 ( .A(n555), .B(KEYINPUT79), .ZN(n540) );
  NOR2_X1 U329 ( .A1(n545), .A2(n416), .ZN(n570) );
  XNOR2_X1 U330 ( .A(KEYINPUT48), .B(KEYINPUT118), .ZN(n396) );
  XNOR2_X1 U331 ( .A(n346), .B(n345), .ZN(n351) );
  XNOR2_X1 U332 ( .A(n397), .B(n396), .ZN(n547) );
  AND2_X1 U333 ( .A1(n450), .A2(n529), .ZN(n565) );
  XNOR2_X1 U334 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n452) );
  XNOR2_X1 U335 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n295) );
  XNOR2_X1 U337 ( .A(G1GAT), .B(G57GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U339 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n297) );
  XNOR2_X1 U340 ( .A(KEYINPUT89), .B(KEYINPUT93), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U342 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U343 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n301) );
  NAND2_X1 U344 ( .A1(G225GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U346 ( .A(KEYINPUT5), .B(n302), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n311) );
  XOR2_X1 U348 ( .A(G148GAT), .B(G162GAT), .Z(n306) );
  XNOR2_X1 U349 ( .A(G120GAT), .B(G155GAT), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U351 ( .A(n307), .B(G85GAT), .Z(n309) );
  XOR2_X1 U352 ( .A(G134GAT), .B(KEYINPUT78), .Z(n337) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(n337), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U355 ( .A(n311), .B(n310), .Z(n316) );
  XOR2_X1 U356 ( .A(G127GAT), .B(KEYINPUT84), .Z(n313) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n445) );
  XNOR2_X1 U359 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U360 ( .A(n314), .B(KEYINPUT2), .ZN(n419) );
  XNOR2_X1 U361 ( .A(n445), .B(n419), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n545) );
  INV_X1 U363 ( .A(KEYINPUT54), .ZN(n415) );
  XOR2_X1 U364 ( .A(G197GAT), .B(G141GAT), .Z(n318) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(G22GAT), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n333) );
  XOR2_X1 U367 ( .A(KEYINPUT67), .B(KEYINPUT65), .Z(n320) );
  XNOR2_X1 U368 ( .A(KEYINPUT30), .B(KEYINPUT64), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U370 ( .A(G36GAT), .B(G50GAT), .Z(n322) );
  XOR2_X1 U371 ( .A(G15GAT), .B(G1GAT), .Z(n358) );
  XOR2_X1 U372 ( .A(G169GAT), .B(G8GAT), .Z(n399) );
  XNOR2_X1 U373 ( .A(n358), .B(n399), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U375 ( .A(n324), .B(n323), .Z(n326) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U378 ( .A(n327), .B(KEYINPUT29), .Z(n331) );
  XOR2_X1 U379 ( .A(G29GAT), .B(G43GAT), .Z(n329) );
  XNOR2_X1 U380 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n349) );
  XNOR2_X1 U382 ( .A(n349), .B(KEYINPUT66), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n335) );
  XNOR2_X1 U385 ( .A(KEYINPUT75), .B(KEYINPUT11), .ZN(n334) );
  XOR2_X1 U386 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U387 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U389 ( .A(G36GAT), .B(G190GAT), .Z(n403) );
  XNOR2_X1 U390 ( .A(n338), .B(n403), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n346) );
  XOR2_X1 U392 ( .A(KEYINPUT70), .B(G92GAT), .Z(n342) );
  XNOR2_X1 U393 ( .A(G99GAT), .B(G85GAT), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(n343), .ZN(n384) );
  NAND2_X1 U396 ( .A1(G232GAT), .A2(G233GAT), .ZN(n344) );
  XOR2_X1 U397 ( .A(G162GAT), .B(KEYINPUT74), .Z(n348) );
  XNOR2_X1 U398 ( .A(G50GAT), .B(G218GAT), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n420) );
  XNOR2_X1 U400 ( .A(n349), .B(n420), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n351), .B(n350), .ZN(n555) );
  XNOR2_X1 U402 ( .A(KEYINPUT36), .B(n540), .ZN(n583) );
  XOR2_X1 U403 ( .A(G57GAT), .B(KEYINPUT13), .Z(n370) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G155GAT), .Z(n426) );
  XOR2_X1 U405 ( .A(n370), .B(n426), .Z(n353) );
  XNOR2_X1 U406 ( .A(G127GAT), .B(G183GAT), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U408 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n355) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U411 ( .A(n357), .B(n356), .Z(n360) );
  XNOR2_X1 U412 ( .A(n358), .B(KEYINPUT12), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n360), .B(n359), .ZN(n368) );
  XOR2_X1 U414 ( .A(G64GAT), .B(G211GAT), .Z(n362) );
  XNOR2_X1 U415 ( .A(G71GAT), .B(G78GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U417 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n364) );
  XNOR2_X1 U418 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U420 ( .A(n366), .B(n365), .Z(n367) );
  XNOR2_X1 U421 ( .A(n368), .B(n367), .ZN(n536) );
  NOR2_X1 U422 ( .A1(n583), .A2(n536), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n369), .B(KEYINPUT45), .ZN(n386) );
  XOR2_X1 U424 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n372) );
  XOR2_X1 U425 ( .A(G176GAT), .B(G64GAT), .Z(n398) );
  XNOR2_X1 U426 ( .A(n370), .B(n398), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U428 ( .A(n373), .B(KEYINPUT72), .Z(n379) );
  XNOR2_X1 U429 ( .A(G78GAT), .B(KEYINPUT69), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n374), .B(G148GAT), .ZN(n417) );
  XOR2_X1 U431 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XOR2_X1 U432 ( .A(n417), .B(n435), .Z(n376) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U435 ( .A(G204GAT), .B(n377), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U437 ( .A(KEYINPUT68), .B(KEYINPUT73), .Z(n381) );
  XNOR2_X1 U438 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n575) );
  NAND2_X1 U442 ( .A1(n386), .A2(n575), .ZN(n387) );
  NOR2_X1 U443 ( .A1(n572), .A2(n387), .ZN(n388) );
  XOR2_X1 U444 ( .A(KEYINPUT117), .B(n388), .Z(n395) );
  XOR2_X1 U445 ( .A(KEYINPUT41), .B(n575), .Z(n533) );
  INV_X1 U446 ( .A(n533), .ZN(n562) );
  NAND2_X1 U447 ( .A1(n562), .A2(n572), .ZN(n390) );
  XNOR2_X1 U448 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n392) );
  INV_X1 U450 ( .A(n536), .ZN(n579) );
  NOR2_X1 U451 ( .A1(n579), .A2(n555), .ZN(n391) );
  AND2_X1 U452 ( .A1(n392), .A2(n391), .ZN(n393) );
  XOR2_X1 U453 ( .A(KEYINPUT47), .B(n393), .Z(n394) );
  NOR2_X1 U454 ( .A1(n395), .A2(n394), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n413) );
  XOR2_X1 U456 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n401) );
  XNOR2_X1 U457 ( .A(G218GAT), .B(G92GAT), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U459 ( .A(n403), .B(n402), .Z(n405) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n411) );
  XOR2_X1 U462 ( .A(G183GAT), .B(KEYINPUT17), .Z(n407) );
  XNOR2_X1 U463 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n444) );
  XOR2_X1 U465 ( .A(G204GAT), .B(G211GAT), .Z(n409) );
  XNOR2_X1 U466 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n418) );
  XOR2_X1 U468 ( .A(n444), .B(n418), .Z(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n477) );
  NOR2_X1 U471 ( .A1(n547), .A2(n477), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U473 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n430) );
  XOR2_X1 U476 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n424) );
  XNOR2_X1 U477 ( .A(G106GAT), .B(KEYINPUT23), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U479 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n465) );
  NAND2_X1 U483 ( .A1(n570), .A2(n465), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n431), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U485 ( .A(G190GAT), .B(G134GAT), .Z(n433) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(G99GAT), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U488 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U489 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n449) );
  XOR2_X1 U491 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n439) );
  XNOR2_X1 U492 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U494 ( .A(G176GAT), .B(KEYINPUT86), .Z(n441) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(G15GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U497 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n468) );
  INV_X1 U501 ( .A(n468), .ZN(n529) );
  INV_X1 U502 ( .A(n540), .ZN(n451) );
  NAND2_X1 U503 ( .A1(n565), .A2(n451), .ZN(n453) );
  NAND2_X1 U504 ( .A1(n540), .A2(n579), .ZN(n454) );
  XNOR2_X1 U505 ( .A(n454), .B(KEYINPUT16), .ZN(n455) );
  XNOR2_X1 U506 ( .A(KEYINPUT83), .B(n455), .ZN(n472) );
  NOR2_X1 U507 ( .A1(n529), .A2(n465), .ZN(n456) );
  XOR2_X1 U508 ( .A(KEYINPUT26), .B(n456), .Z(n569) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n457), .B(n477), .ZN(n466) );
  NOR2_X1 U511 ( .A1(n569), .A2(n466), .ZN(n544) );
  INV_X1 U512 ( .A(n465), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n468), .A2(n477), .ZN(n458) );
  NOR2_X1 U514 ( .A1(n459), .A2(n458), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n460) );
  XNOR2_X1 U516 ( .A(n461), .B(n460), .ZN(n462) );
  NOR2_X1 U517 ( .A1(n544), .A2(n462), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n545), .A2(n463), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(KEYINPUT99), .ZN(n471) );
  XOR2_X1 U520 ( .A(KEYINPUT28), .B(n465), .Z(n521) );
  NOR2_X1 U521 ( .A1(n466), .A2(n521), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n545), .A2(n467), .ZN(n527) );
  XNOR2_X1 U523 ( .A(KEYINPUT97), .B(n527), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n486) );
  NAND2_X1 U526 ( .A1(n472), .A2(n486), .ZN(n473) );
  XNOR2_X1 U527 ( .A(n473), .B(KEYINPUT100), .ZN(n504) );
  NAND2_X1 U528 ( .A1(n572), .A2(n575), .ZN(n490) );
  NOR2_X1 U529 ( .A1(n504), .A2(n490), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT101), .B(n474), .Z(n483) );
  NAND2_X1 U531 ( .A1(n483), .A2(n545), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n475), .B(KEYINPUT34), .ZN(n476) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  INV_X1 U534 ( .A(n477), .ZN(n518) );
  NAND2_X1 U535 ( .A1(n483), .A2(n518), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT102), .ZN(n479) );
  XNOR2_X1 U537 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n481) );
  NAND2_X1 U539 ( .A1(n483), .A2(n529), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U541 ( .A(G15GAT), .B(n482), .Z(G1326GAT) );
  NAND2_X1 U542 ( .A1(n521), .A2(n483), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(KEYINPUT104), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G22GAT), .B(n485), .ZN(G1327GAT) );
  XNOR2_X1 U545 ( .A(KEYINPUT105), .B(KEYINPUT39), .ZN(n497) );
  XOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT109), .Z(n495) );
  NAND2_X1 U547 ( .A1(n536), .A2(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(KEYINPUT106), .B(n487), .ZN(n488) );
  NOR2_X1 U549 ( .A1(n488), .A2(n583), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT37), .ZN(n515) );
  NOR2_X1 U551 ( .A1(n515), .A2(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT38), .B(KEYINPUT107), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U554 ( .A(KEYINPUT108), .B(n493), .Z(n501) );
  NAND2_X1 U555 ( .A1(n501), .A2(n545), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n518), .A2(n501), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n501), .A2(n529), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(KEYINPUT40), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NAND2_X1 U563 ( .A1(n521), .A2(n501), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n506) );
  INV_X1 U566 ( .A(n572), .ZN(n530) );
  NAND2_X1 U567 ( .A1(n530), .A2(n562), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(KEYINPUT110), .ZN(n516) );
  NOR2_X1 U569 ( .A1(n516), .A2(n504), .ZN(n510) );
  NAND2_X1 U570 ( .A1(n510), .A2(n545), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n518), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n529), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n509), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U578 ( .A1(n510), .A2(n521), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(n514) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT112), .Z(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n522) );
  NAND2_X1 U583 ( .A1(n522), .A2(n545), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n522), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n529), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(KEYINPUT115), .ZN(n526) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n524) );
  NAND2_X1 U591 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n547), .A2(n527), .ZN(n528) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n539) );
  NOR2_X1 U596 ( .A1(n530), .A2(n539), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(KEYINPUT119), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n539), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n539), .ZN(n537) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(n537), .Z(n538) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U606 ( .A(KEYINPUT120), .B(KEYINPUT51), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n543), .ZN(G1343GAT) );
  XOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT121), .Z(n549) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n556), .A2(n572), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U615 ( .A1(n556), .A2(n562), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n556), .A2(n579), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT122), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n572), .A2(n565), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT123), .B(n561), .Z(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n579), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n574) );
  INV_X1 U636 ( .A(n569), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n582) );
  INV_X1 U638 ( .A(n582), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n580), .A2(n572), .ZN(n573) );
  XOR2_X1 U640 ( .A(n574), .B(n573), .Z(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n577) );
  OR2_X1 U642 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

