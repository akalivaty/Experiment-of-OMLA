

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U324 ( .A(n421), .B(n292), .ZN(n422) );
  AND2_X1 U325 ( .A1(G231GAT), .A2(G233GAT), .ZN(n291) );
  AND2_X1 U326 ( .A1(G225GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U327 ( .A(G71GAT), .B(G211GAT), .Z(n293) );
  XOR2_X1 U328 ( .A(n411), .B(n410), .Z(n294) );
  XNOR2_X1 U329 ( .A(n435), .B(n291), .ZN(n437) );
  XNOR2_X1 U330 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U331 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n469) );
  XNOR2_X1 U332 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U333 ( .A(n442), .B(n293), .ZN(n443) );
  XNOR2_X1 U334 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U335 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n449) );
  XNOR2_X1 U336 ( .A(n450), .B(n449), .ZN(n509) );
  NOR2_X1 U337 ( .A1(n476), .A2(n475), .ZN(n562) );
  XNOR2_X1 U338 ( .A(n477), .B(G190GAT), .ZN(n478) );
  XNOR2_X1 U339 ( .A(n452), .B(G43GAT), .ZN(n453) );
  XNOR2_X1 U340 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT79), .B(G134GAT), .Z(n296) );
  XNOR2_X1 U343 ( .A(KEYINPUT0), .B(G113GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U345 ( .A(KEYINPUT80), .B(n297), .Z(n410) );
  XOR2_X1 U346 ( .A(KEYINPUT82), .B(G190GAT), .Z(n299) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G99GAT), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U349 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n301) );
  XNOR2_X1 U350 ( .A(G183GAT), .B(KEYINPUT20), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U352 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U353 ( .A(G127GAT), .B(G15GAT), .Z(n435) );
  XOR2_X1 U354 ( .A(G120GAT), .B(G71GAT), .Z(n316) );
  XOR2_X1 U355 ( .A(G176GAT), .B(n316), .Z(n305) );
  NAND2_X1 U356 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n435), .B(n306), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n410), .B(n309), .ZN(n313) );
  XOR2_X1 U361 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n311) );
  XNOR2_X1 U362 ( .A(KEYINPUT84), .B(G169GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U364 ( .A(KEYINPUT18), .B(n312), .Z(n400) );
  XNOR2_X1 U365 ( .A(n313), .B(n400), .ZN(n526) );
  XOR2_X1 U366 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n315) );
  XNOR2_X1 U367 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n320) );
  XOR2_X1 U369 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n318) );
  XOR2_X1 U370 ( .A(G85GAT), .B(G99GAT), .Z(n357) );
  XNOR2_X1 U371 ( .A(n357), .B(n316), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U373 ( .A(n320), .B(n319), .Z(n322) );
  NAND2_X1 U374 ( .A1(G230GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n324) );
  XNOR2_X1 U376 ( .A(G148GAT), .B(G106GAT), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n323), .B(G78GAT), .ZN(n382) );
  XOR2_X1 U378 ( .A(n324), .B(n382), .Z(n330) );
  XNOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n325), .B(KEYINPUT13), .ZN(n439) );
  XOR2_X1 U381 ( .A(KEYINPUT72), .B(G204GAT), .Z(n327) );
  XNOR2_X1 U382 ( .A(G92GAT), .B(G176GAT), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U384 ( .A(G64GAT), .B(n328), .Z(n393) );
  XNOR2_X1 U385 ( .A(n439), .B(n393), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n570) );
  XOR2_X1 U387 ( .A(KEYINPUT64), .B(KEYINPUT67), .Z(n332) );
  XNOR2_X1 U388 ( .A(KEYINPUT29), .B(KEYINPUT65), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n345) );
  XOR2_X1 U390 ( .A(G169GAT), .B(G15GAT), .Z(n334) );
  XNOR2_X1 U391 ( .A(G50GAT), .B(G36GAT), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U393 ( .A(G197GAT), .B(G8GAT), .Z(n336) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(G113GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U396 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U397 ( .A(G1GAT), .B(G22GAT), .Z(n442) );
  XOR2_X1 U398 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n340) );
  NAND2_X1 U399 ( .A1(G229GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n442), .B(n341), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U404 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n347) );
  XNOR2_X1 U405 ( .A(KEYINPUT7), .B(G43GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U407 ( .A(G29GAT), .B(n348), .ZN(n362) );
  XNOR2_X1 U408 ( .A(n349), .B(n362), .ZN(n566) );
  NAND2_X1 U409 ( .A1(n570), .A2(n566), .ZN(n483) );
  XOR2_X1 U410 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n351) );
  XNOR2_X1 U411 ( .A(KEYINPUT75), .B(KEYINPUT10), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n366) );
  XOR2_X1 U413 ( .A(G106GAT), .B(KEYINPUT11), .Z(n353) );
  XNOR2_X1 U414 ( .A(KEYINPUT76), .B(G92GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U416 ( .A(n354), .B(G218GAT), .Z(n356) );
  XOR2_X1 U417 ( .A(G190GAT), .B(G36GAT), .Z(n396) );
  XNOR2_X1 U418 ( .A(G134GAT), .B(n396), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n361) );
  XOR2_X1 U420 ( .A(n357), .B(KEYINPUT74), .Z(n359) );
  NAND2_X1 U421 ( .A1(G232GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U423 ( .A(n361), .B(n360), .Z(n364) );
  XOR2_X1 U424 ( .A(G162GAT), .B(G50GAT), .Z(n383) );
  XOR2_X1 U425 ( .A(n362), .B(n383), .Z(n363) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U427 ( .A(n366), .B(n365), .Z(n538) );
  XNOR2_X1 U428 ( .A(n538), .B(KEYINPUT102), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n367), .B(KEYINPUT36), .ZN(n580) );
  XOR2_X1 U430 ( .A(G197GAT), .B(KEYINPUT88), .Z(n369) );
  XNOR2_X1 U431 ( .A(KEYINPUT89), .B(KEYINPUT21), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U433 ( .A(n370), .B(KEYINPUT87), .Z(n372) );
  XNOR2_X1 U434 ( .A(G218GAT), .B(G211GAT), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n395) );
  XOR2_X1 U436 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n374) );
  XNOR2_X1 U437 ( .A(G22GAT), .B(KEYINPUT85), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U439 ( .A(KEYINPUT86), .B(KEYINPUT91), .Z(n376) );
  XNOR2_X1 U440 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U442 ( .A(n378), .B(n377), .Z(n388) );
  XOR2_X1 U443 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n380) );
  XNOR2_X1 U444 ( .A(G155GAT), .B(G141GAT), .ZN(n379) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U446 ( .A(KEYINPUT3), .B(n381), .Z(n425) );
  XOR2_X1 U447 ( .A(n383), .B(n382), .Z(n385) );
  NAND2_X1 U448 ( .A1(G228GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n425), .B(n386), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(n395), .B(n389), .Z(n473) );
  XNOR2_X1 U453 ( .A(G183GAT), .B(G8GAT), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n390), .B(KEYINPUT78), .ZN(n436) );
  XOR2_X1 U455 ( .A(KEYINPUT96), .B(n436), .Z(n392) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U458 ( .A(n394), .B(n393), .Z(n398) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n467) );
  INV_X1 U462 ( .A(n526), .ZN(n476) );
  NOR2_X1 U463 ( .A1(n467), .A2(n476), .ZN(n401) );
  NOR2_X1 U464 ( .A1(n473), .A2(n401), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n402), .B(KEYINPUT25), .ZN(n407) );
  AND2_X1 U466 ( .A1(n473), .A2(n476), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n403), .B(KEYINPUT100), .ZN(n404) );
  XOR2_X1 U468 ( .A(KEYINPUT26), .B(n404), .Z(n565) );
  INV_X1 U469 ( .A(n565), .ZN(n542) );
  XNOR2_X1 U470 ( .A(KEYINPUT97), .B(KEYINPUT27), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n405), .B(n467), .ZN(n427) );
  NAND2_X1 U472 ( .A1(n542), .A2(n427), .ZN(n406) );
  NAND2_X1 U473 ( .A1(n407), .A2(n406), .ZN(n426) );
  XOR2_X1 U474 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n409) );
  XNOR2_X1 U475 ( .A(KEYINPUT5), .B(KEYINPUT92), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U477 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n413) );
  XNOR2_X1 U478 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U480 ( .A(G148GAT), .B(G120GAT), .Z(n415) );
  XNOR2_X1 U481 ( .A(G29GAT), .B(G127GAT), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n294), .B(n418), .ZN(n423) );
  XOR2_X1 U485 ( .A(G85GAT), .B(G162GAT), .Z(n420) );
  XNOR2_X1 U486 ( .A(G57GAT), .B(G1GAT), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n471) );
  NAND2_X1 U489 ( .A1(n426), .A2(n471), .ZN(n432) );
  INV_X1 U490 ( .A(n471), .ZN(n510) );
  AND2_X1 U491 ( .A1(n510), .A2(n427), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n428), .B(KEYINPUT98), .ZN(n541) );
  XNOR2_X1 U493 ( .A(KEYINPUT28), .B(n473), .ZN(n519) );
  INV_X1 U494 ( .A(n519), .ZN(n429) );
  NAND2_X1 U495 ( .A1(n541), .A2(n429), .ZN(n524) );
  XNOR2_X1 U496 ( .A(n524), .B(KEYINPUT99), .ZN(n430) );
  NAND2_X1 U497 ( .A1(n430), .A2(n476), .ZN(n431) );
  NAND2_X1 U498 ( .A1(n432), .A2(n431), .ZN(n481) );
  XOR2_X1 U499 ( .A(KEYINPUT15), .B(G64GAT), .Z(n434) );
  XNOR2_X1 U500 ( .A(G155GAT), .B(G78GAT), .ZN(n433) );
  XNOR2_X1 U501 ( .A(n434), .B(n433), .ZN(n446) );
  XOR2_X1 U502 ( .A(n438), .B(KEYINPUT14), .Z(n441) );
  XNOR2_X1 U503 ( .A(n439), .B(KEYINPUT12), .ZN(n440) );
  XNOR2_X1 U504 ( .A(n441), .B(n440), .ZN(n444) );
  XOR2_X1 U505 ( .A(n446), .B(n445), .Z(n550) );
  NAND2_X1 U506 ( .A1(n481), .A2(n550), .ZN(n447) );
  XOR2_X1 U507 ( .A(n447), .B(KEYINPUT103), .Z(n448) );
  NOR2_X1 U508 ( .A1(n580), .A2(n448), .ZN(n450) );
  NOR2_X1 U509 ( .A1(n483), .A2(n509), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n451), .B(KEYINPUT38), .ZN(n495) );
  NAND2_X1 U511 ( .A1(n526), .A2(n495), .ZN(n454) );
  XOR2_X1 U512 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n452) );
  NOR2_X1 U513 ( .A1(n580), .A2(n550), .ZN(n455) );
  XNOR2_X1 U514 ( .A(KEYINPUT45), .B(n455), .ZN(n456) );
  NAND2_X1 U515 ( .A1(n456), .A2(n570), .ZN(n457) );
  NOR2_X1 U516 ( .A1(n566), .A2(n457), .ZN(n465) );
  INV_X1 U517 ( .A(KEYINPUT47), .ZN(n463) );
  XOR2_X1 U518 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n459) );
  XNOR2_X1 U519 ( .A(n570), .B(KEYINPUT41), .ZN(n558) );
  NAND2_X1 U520 ( .A1(n558), .A2(n566), .ZN(n458) );
  XNOR2_X1 U521 ( .A(n459), .B(n458), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n538), .A2(n550), .ZN(n460) );
  NOR2_X1 U523 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n463), .B(n462), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U526 ( .A(KEYINPUT48), .B(n466), .ZN(n544) );
  INV_X1 U527 ( .A(n467), .ZN(n514) );
  XNOR2_X1 U528 ( .A(KEYINPUT121), .B(n514), .ZN(n468) );
  NOR2_X1 U529 ( .A1(n544), .A2(n468), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n564) );
  NOR2_X1 U531 ( .A1(n473), .A2(n564), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT55), .ZN(n475) );
  INV_X1 U533 ( .A(n538), .ZN(n554) );
  NAND2_X1 U534 ( .A1(n562), .A2(n554), .ZN(n479) );
  XOR2_X1 U535 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n485) );
  NOR2_X1 U537 ( .A1(n550), .A2(n554), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT16), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n497) );
  NOR2_X1 U540 ( .A1(n483), .A2(n497), .ZN(n490) );
  NAND2_X1 U541 ( .A1(n490), .A2(n510), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U544 ( .A1(n490), .A2(n514), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U547 ( .A1(n490), .A2(n526), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  NAND2_X1 U549 ( .A1(n519), .A2(n490), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  NAND2_X1 U552 ( .A1(n510), .A2(n495), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n495), .A2(n514), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U556 ( .A1(n495), .A2(n519), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n500) );
  INV_X1 U559 ( .A(n566), .ZN(n527) );
  NAND2_X1 U560 ( .A1(n527), .A2(n558), .ZN(n508) );
  NOR2_X1 U561 ( .A1(n508), .A2(n497), .ZN(n498) );
  XNOR2_X1 U562 ( .A(KEYINPUT106), .B(n498), .ZN(n504) );
  NAND2_X1 U563 ( .A1(n510), .A2(n504), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n514), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n504), .A2(n526), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n503), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U571 ( .A1(n504), .A2(n519), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(n507), .ZN(G1335GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n512) );
  NOR2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n520) );
  NAND2_X1 U576 ( .A1(n520), .A2(n510), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n516) );
  NAND2_X1 U580 ( .A1(n520), .A2(n514), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n526), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n522) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n544), .ZN(n525) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n527), .A2(n537), .ZN(n528) );
  XOR2_X1 U592 ( .A(G113GAT), .B(n528), .Z(G1340GAT) );
  INV_X1 U593 ( .A(n558), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n537), .A2(n529), .ZN(n533) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n531) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT116), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n550), .A2(n537), .ZN(n535) );
  XNOR2_X1 U600 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n566), .A2(n553), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n545), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n547) );
  NAND2_X1 U612 ( .A1(n553), .A2(n558), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  XOR2_X1 U615 ( .A(G155GAT), .B(KEYINPUT119), .Z(n552) );
  INV_X1 U616 ( .A(n550), .ZN(n576) );
  NAND2_X1 U617 ( .A1(n553), .A2(n576), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT120), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n562), .A2(n566), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n562), .A2(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n576), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n575), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  INV_X1 U635 ( .A(n575), .ZN(n579) );
  NOR2_X1 U636 ( .A1(n579), .A2(n570), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT126), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

