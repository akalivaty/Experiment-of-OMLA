//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT65), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n191), .A3(G143), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n188), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n195), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n188), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n189), .A2(new_n191), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n198), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(G137), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n206), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n207), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n204), .A2(new_n205), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n205), .B1(new_n204), .B2(new_n217), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n212), .A2(new_n214), .A3(new_n207), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n216), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT65), .B(G146), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n199), .B1(new_n224), .B2(G143), .ZN(new_n225));
  XOR2_X1   g039(.A(KEYINPUT0), .B(G128), .Z(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n192), .A2(KEYINPUT0), .A3(G128), .A4(new_n194), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n223), .A2(new_n227), .A3(KEYINPUT66), .A4(new_n228), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n187), .B1(new_n220), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT68), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT2), .B(G113), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n237), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n239), .B1(KEYINPUT68), .B2(new_n235), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n204), .A2(new_n217), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT30), .A3(new_n229), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n234), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n241), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n229), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT26), .B(G101), .Z(new_n248));
  NOR2_X1   g062(.A1(G237), .A2(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G210), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n248), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n246), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT70), .B1(new_n256), .B2(KEYINPUT28), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n246), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n231), .B(new_n232), .C1(new_n218), .C2(new_n219), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n256), .B1(new_n262), .B2(new_n241), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n261), .B(new_n253), .C1(new_n259), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n255), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n245), .B1(new_n242), .B2(new_n229), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT28), .B1(new_n256), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n254), .A2(new_n265), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n257), .A2(new_n268), .A3(new_n260), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n270), .A2(KEYINPUT71), .A3(new_n271), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G472), .B1(new_n266), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n244), .A2(new_n253), .A3(new_n246), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT31), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n263), .A2(new_n259), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n257), .A2(new_n260), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n254), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n244), .A2(new_n283), .A3(new_n253), .A4(new_n246), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  NOR2_X1   g100(.A1(G472), .A2(G902), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n277), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G469), .ZN(new_n291));
  XNOR2_X1  g105(.A(G110), .B(G140), .ZN(new_n292));
  INV_X1    g106(.A(G953), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n293), .A2(G227), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n292), .B(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT82), .ZN(new_n297));
  INV_X1    g111(.A(new_n226), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n228), .B1(new_n203), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G104), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT3), .B1(new_n301), .B2(G107), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n303));
  INV_X1    g117(.A(G107), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(G104), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n301), .A2(G107), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(G101), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(G101), .ZN(new_n310));
  INV_X1    g124(.A(G101), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n302), .A2(new_n305), .A3(new_n311), .A4(new_n306), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n310), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n300), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n193), .B1(new_n224), .B2(G143), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n195), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n197), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n301), .A2(G107), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n304), .A2(G104), .ZN(new_n319));
  OAI21_X1  g133(.A(G101), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT10), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT81), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n312), .A2(new_n320), .A3(KEYINPUT10), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n204), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n326), .B1(new_n204), .B2(new_n327), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n314), .B(new_n325), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n297), .B1(new_n330), .B2(new_n223), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n313), .A2(new_n309), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n332), .A2(new_n300), .B1(new_n324), .B2(new_n323), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n204), .A2(new_n327), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT81), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n204), .A2(new_n326), .A3(new_n327), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n222), .A2(new_n216), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n333), .A2(new_n337), .A3(KEYINPUT82), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n330), .A2(new_n223), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n296), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n321), .B(new_n197), .C1(new_n198), .C2(new_n203), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n323), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT12), .B1(new_n344), .B2(new_n223), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT12), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n346), .B(new_n338), .C1(new_n323), .C2(new_n343), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI211_X1 g162(.A(new_n295), .B(new_n348), .C1(new_n331), .C2(new_n339), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n291), .B(new_n271), .C1(new_n342), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(G469), .A2(G902), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n340), .A2(new_n341), .A3(new_n296), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n348), .B1(new_n331), .B2(new_n339), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n352), .B(G469), .C1(new_n296), .C2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT9), .B(G234), .ZN(new_n356));
  OAI21_X1  g170(.A(G221), .B1(new_n356), .B2(G902), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT79), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G214), .B1(G237), .B2(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(G210), .B1(G237), .B2(G902), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n299), .A2(G125), .ZN(new_n364));
  INV_X1    g178(.A(G125), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(new_n197), .C1(new_n198), .C2(new_n203), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n293), .A2(G224), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n364), .A2(new_n366), .B1(KEYINPUT7), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT7), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n371), .B2(new_n367), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n364), .A2(new_n366), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G122), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT8), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n379));
  INV_X1    g193(.A(G119), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G116), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n379), .B(G113), .C1(KEYINPUT5), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n239), .A2(new_n235), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n322), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n322), .B1(new_n383), .B2(new_n382), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n378), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n313), .A2(new_n241), .A3(new_n309), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n384), .A3(new_n377), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n364), .A2(KEYINPUT86), .A3(new_n366), .A4(new_n373), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n376), .A2(new_n387), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n271), .B1(new_n370), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n384), .ZN(new_n393));
  INV_X1    g207(.A(new_n377), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(KEYINPUT83), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n389), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n364), .A2(new_n366), .ZN(new_n399));
  INV_X1    g213(.A(new_n367), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n393), .B(new_n394), .C1(KEYINPUT83), .C2(new_n396), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n363), .B1(new_n392), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n368), .B(KEYINPUT84), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n376), .A2(new_n390), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n405), .A2(new_n389), .A3(new_n387), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n407), .A2(new_n271), .A3(new_n362), .A4(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n361), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n355), .A2(new_n359), .A3(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n412));
  AOI21_X1  g226(.A(G140), .B1(KEYINPUT75), .B2(G125), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT16), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n365), .A2(G140), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT16), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n419), .B(KEYINPUT16), .C1(new_n412), .C2(new_n413), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(G146), .A3(new_n418), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT78), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT75), .A2(G125), .ZN(new_n423));
  INV_X1    g237(.A(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n417), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n427), .A2(new_n419), .B1(new_n417), .B2(new_n416), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT78), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n428), .A2(new_n429), .A3(G146), .A4(new_n415), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n249), .A2(G143), .A3(G214), .ZN(new_n431));
  AOI21_X1  g245(.A(G143), .B1(new_n249), .B2(G214), .ZN(new_n432));
  OAI21_X1  g246(.A(G131), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n249), .A2(G214), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n202), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n249), .A2(G143), .A3(G214), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n215), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G125), .B(G140), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT19), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n425), .A2(KEYINPUT19), .A3(new_n426), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(KEYINPUT87), .A3(new_n440), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n224), .A4(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n422), .A2(new_n430), .A3(new_n438), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n435), .A2(new_n436), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT18), .A3(G131), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n224), .A2(new_n439), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n425), .A2(new_n426), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n188), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(KEYINPUT18), .A2(G131), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n435), .A2(new_n436), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n447), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G113), .B(G122), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(new_n301), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n420), .A2(new_n418), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n419), .B1(new_n451), .B2(KEYINPUT16), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n188), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT17), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n433), .A2(new_n437), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n448), .A2(KEYINPUT17), .A3(G131), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n463), .A2(new_n465), .A3(new_n421), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n455), .A3(new_n458), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n460), .A2(KEYINPUT88), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(G475), .A2(G902), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n458), .B1(new_n447), .B2(new_n455), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n467), .A2(new_n455), .A3(new_n458), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT20), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n475), .B2(KEYINPUT20), .ZN(new_n478));
  NOR3_X1   g292(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n472), .B2(new_n473), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n458), .B1(new_n467), .B2(new_n455), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n271), .B1(new_n473), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G475), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G478), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT13), .B1(new_n195), .B2(G143), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n206), .ZN(new_n491));
  XNOR2_X1  g305(.A(G128), .B(G143), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G122), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G116), .ZN(new_n495));
  INV_X1    g309(.A(G116), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G122), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n495), .B2(new_n497), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n500), .A2(new_n304), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n501), .ZN(new_n503));
  AOI21_X1  g317(.A(G107), .B1(new_n503), .B2(new_n499), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n493), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n304), .B1(new_n500), .B2(new_n501), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n492), .B(new_n206), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n496), .A2(KEYINPUT14), .A3(G122), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n495), .A2(new_n497), .ZN(new_n509));
  OAI211_X1 g323(.A(G107), .B(new_n508), .C1(new_n509), .C2(KEYINPUT14), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G217), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n356), .A2(new_n512), .A3(G953), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT91), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n505), .A2(new_n511), .A3(new_n516), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n505), .A2(new_n511), .ZN(new_n518));
  INV_X1    g332(.A(new_n513), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n521), .A2(KEYINPUT93), .A3(new_n271), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT93), .B1(new_n521), .B2(new_n271), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n489), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n271), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT93), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n488), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n293), .A2(G952), .ZN(new_n529));
  NAND2_X1  g343(.A1(G234), .A2(G237), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n530), .A2(G902), .A3(G953), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT21), .B(G898), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR4_X1   g349(.A1(new_n482), .A2(new_n486), .A3(new_n528), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n512), .B1(G234), .B2(new_n271), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n380), .A2(G128), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n380), .A2(KEYINPUT72), .A3(G128), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n541), .B(new_n542), .C1(new_n380), .C2(G128), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT24), .B(G110), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT73), .B1(new_n380), .B2(G128), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT23), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT23), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT73), .B(new_n548), .C1(new_n380), .C2(G128), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n549), .A3(new_n539), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n545), .B1(G110), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n422), .A2(new_n551), .A3(new_n430), .A4(new_n450), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n543), .A2(new_n544), .ZN(new_n553));
  INV_X1    g367(.A(new_n550), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT74), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT74), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n556), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n553), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n463), .A2(new_n421), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n559), .A2(KEYINPUT77), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT77), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n552), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT22), .B(G137), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n293), .A2(G221), .A3(G234), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n552), .B(new_n566), .C1(new_n561), .C2(new_n562), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n271), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT25), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n568), .A2(KEYINPUT25), .A3(new_n271), .A4(new_n569), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n538), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n568), .A2(new_n569), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n537), .A2(G902), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n290), .A2(new_n411), .A3(new_n536), .A4(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(G101), .ZN(G3));
  AND3_X1   g394(.A1(new_n578), .A2(new_n355), .A3(new_n359), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n285), .A2(new_n271), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n582), .A2(G472), .B1(new_n287), .B2(new_n285), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI211_X1 g398(.A(new_n361), .B(new_n535), .C1(new_n404), .C2(new_n409), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n520), .A2(KEYINPUT33), .A3(new_n514), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n586), .A2(KEYINPUT94), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n521), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(KEYINPUT94), .ZN(new_n590));
  INV_X1    g404(.A(G478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(G902), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n587), .A2(new_n589), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n525), .A2(new_n591), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n585), .B(new_n596), .C1(new_n482), .C2(new_n486), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n584), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT34), .B(G104), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G6));
  INV_X1    g415(.A(new_n410), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n475), .A2(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT89), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT20), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n469), .A2(new_n474), .A3(new_n479), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n535), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n486), .B1(new_n524), .B2(new_n527), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n602), .B1(new_n610), .B2(KEYINPUT95), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n607), .A2(new_n612), .A3(new_n608), .A4(new_n609), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n611), .A2(KEYINPUT96), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT96), .B1(new_n611), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n584), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NAND2_X1  g432(.A1(new_n572), .A2(new_n573), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n537), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n563), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n576), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n411), .A2(new_n536), .A3(new_n583), .A4(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  INV_X1    g441(.A(G900), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n532), .B1(new_n533), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n607), .A2(new_n609), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n607), .A2(new_n633), .A3(new_n609), .A4(new_n630), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n410), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n355), .A2(new_n359), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n290), .A2(new_n638), .A3(new_n624), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n632), .A2(KEYINPUT98), .A3(new_n410), .A4(new_n634), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT99), .B(G128), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G30));
  XOR2_X1   g457(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n629), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT40), .Z(new_n647));
  INV_X1    g461(.A(new_n247), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n254), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n256), .A2(new_n267), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n650), .B2(new_n254), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n288), .B2(new_n289), .ZN(new_n654));
  INV_X1    g468(.A(new_n528), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n624), .A2(new_n361), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n604), .A2(new_n605), .A3(new_n480), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n485), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n404), .A2(new_n409), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT38), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n656), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n647), .A2(new_n654), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G143), .ZN(G45));
  AOI211_X1 g477(.A(new_n595), .B(new_n629), .C1(new_n657), .C2(new_n485), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n290), .A2(new_n411), .A3(new_n664), .A4(new_n624), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  OAI21_X1  g480(.A(new_n271), .B1(new_n342), .B2(new_n349), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n291), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  OAI221_X1 g484(.A(new_n271), .B1(new_n668), .B2(new_n291), .C1(new_n342), .C2(new_n349), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n670), .A2(new_n671), .A3(new_n357), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n598), .A2(new_n290), .A3(new_n578), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT41), .B(G113), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G15));
  NAND2_X1  g489(.A1(new_n290), .A2(new_n578), .ZN(new_n676));
  INV_X1    g490(.A(new_n672), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(new_n614), .B2(new_n615), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  AND4_X1   g494(.A1(new_n357), .A2(new_n670), .A3(new_n410), .A4(new_n671), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n290), .A2(new_n536), .A3(new_n681), .A4(new_n624), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G119), .ZN(G21));
  AND4_X1   g497(.A1(new_n357), .A2(new_n670), .A3(new_n608), .A4(new_n671), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n659), .A2(new_n528), .A3(new_n360), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n657), .B2(new_n485), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n261), .A2(new_n268), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n279), .B(new_n284), .C1(new_n253), .C2(new_n687), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n582), .A2(G472), .B1(new_n287), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n684), .A2(new_n686), .A3(new_n578), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  NAND4_X1  g505(.A1(new_n664), .A2(new_n681), .A3(new_n624), .A4(new_n689), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G125), .ZN(G27));
  INV_X1    g507(.A(new_n578), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n285), .A2(new_n287), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT32), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n694), .B1(new_n698), .B2(new_n277), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n659), .A2(new_n361), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n355), .A2(new_n357), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n699), .A2(KEYINPUT42), .A3(new_n664), .A4(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n290), .A2(new_n701), .A3(new_n664), .A4(new_n578), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G131), .ZN(G33));
  AND2_X1   g521(.A1(new_n632), .A2(new_n634), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n699), .A3(new_n709), .A4(new_n701), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n290), .A2(new_n701), .A3(new_n578), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n632), .A2(new_n634), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT102), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G134), .ZN(G36));
  OAI21_X1  g529(.A(new_n352), .B1(new_n296), .B2(new_n353), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n291), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n717), .B2(new_n716), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n351), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(KEYINPUT46), .A3(new_n351), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n350), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n357), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n645), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(KEYINPUT103), .A3(new_n645), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n732));
  OAI22_X1  g546(.A1(new_n658), .A2(new_n595), .B1(KEYINPUT104), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n482), .A2(new_n486), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n596), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n624), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n583), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n700), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n741), .B2(new_n740), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n731), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G137), .ZN(G39));
  XOR2_X1   g559(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n746));
  AND3_X1   g560(.A1(new_n724), .A2(new_n357), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n725), .B1(new_n749), .B2(KEYINPUT47), .ZN(new_n750));
  INV_X1    g564(.A(new_n664), .ZN(new_n751));
  INV_X1    g565(.A(new_n700), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n751), .A2(new_n290), .A3(new_n578), .A4(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n748), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  AND2_X1   g569(.A1(new_n737), .A2(new_n532), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n677), .A2(new_n752), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n676), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT48), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n761));
  INV_X1    g575(.A(new_n654), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n578), .A3(new_n532), .A4(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT113), .Z(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n658), .A3(new_n596), .ZN(new_n765));
  INV_X1    g579(.A(new_n689), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n694), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n756), .A2(new_n681), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n529), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n760), .B1(new_n761), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n758), .A2(new_n738), .A3(new_n766), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n658), .A2(new_n596), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n771), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n677), .A2(new_n360), .A3(new_n660), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n756), .A2(new_n767), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n670), .A2(new_n671), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n359), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n748), .B2(new_n750), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n756), .A2(new_n767), .A3(new_n700), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n773), .B(new_n778), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n783), .A2(KEYINPUT114), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT114), .B1(new_n783), .B2(new_n784), .ZN(new_n786));
  OAI221_X1 g600(.A(new_n770), .B1(new_n761), .B2(new_n769), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n783), .A2(new_n784), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT115), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n355), .A2(new_n357), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n620), .A2(new_n623), .A3(new_n630), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n654), .A2(new_n686), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n665), .A2(new_n794), .A3(new_n692), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n795), .A2(KEYINPUT108), .A3(new_n641), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT108), .B1(new_n795), .B2(new_n641), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n791), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n596), .B1(new_n482), .B2(new_n486), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT106), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT106), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n658), .A2(new_n801), .A3(new_n596), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n585), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT107), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT107), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n800), .A2(new_n805), .A3(new_n585), .A4(new_n802), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n584), .A3(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n673), .A2(new_n579), .A3(new_n625), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n658), .A2(new_n655), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n581), .A2(new_n585), .A3(new_n809), .A4(new_n583), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n810), .A2(new_n682), .A3(new_n690), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n808), .A3(new_n679), .A4(new_n811), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n485), .A2(new_n607), .A3(new_n655), .A4(new_n630), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n290), .A2(new_n638), .A3(new_n813), .A4(new_n624), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n664), .A2(new_n792), .A3(new_n624), .A4(new_n689), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n700), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n714), .A2(new_n706), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n665), .A2(new_n794), .A3(new_n692), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n795), .A2(new_n641), .A3(KEYINPUT108), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(KEYINPUT52), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n798), .A2(new_n819), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT110), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(new_n823), .B2(new_n824), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n791), .B1(new_n795), .B2(new_n641), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT109), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n831), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n798), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT53), .B1(new_n836), .B2(new_n819), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT54), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n819), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT111), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n826), .B2(new_n827), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n826), .A2(new_n841), .A3(new_n827), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n839), .B(new_n840), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n790), .A2(new_n838), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(G952), .B2(G953), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n779), .B(KEYINPUT49), .Z(new_n847));
  NAND3_X1  g661(.A1(new_n596), .A2(new_n359), .A3(new_n360), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n660), .A2(new_n694), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n734), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n846), .B1(new_n654), .B2(new_n850), .ZN(G75));
  NOR2_X1   g665(.A1(new_n293), .A2(G952), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n271), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT56), .B1(new_n856), .B2(G210), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n398), .A2(new_n402), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(new_n401), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT55), .Z(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n853), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n857), .B2(new_n861), .ZN(G51));
  NOR2_X1   g677(.A1(new_n843), .A2(new_n842), .ZN(new_n864));
  INV_X1    g678(.A(new_n819), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n827), .B(new_n865), .C1(new_n832), .C2(new_n835), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT54), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(KEYINPUT117), .A3(new_n844), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n854), .A2(new_n869), .A3(KEYINPUT54), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n351), .B(KEYINPUT57), .Z(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n342), .A2(new_n349), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n868), .A2(KEYINPUT118), .A3(new_n870), .A4(new_n871), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OR3_X1    g691(.A1(new_n855), .A2(new_n271), .A3(new_n719), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n852), .B1(new_n877), .B2(new_n878), .ZN(G54));
  NAND3_X1  g693(.A1(new_n856), .A2(KEYINPUT58), .A3(G475), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n469), .A2(new_n474), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(new_n852), .ZN(G60));
  XNOR2_X1  g698(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n591), .A2(new_n271), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n885), .B(new_n886), .Z(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n838), .B2(new_n844), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT119), .Z(new_n890));
  OAI21_X1  g704(.A(new_n853), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n868), .A2(new_n870), .ZN(new_n892));
  INV_X1    g706(.A(new_n887), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n891), .B1(new_n892), .B2(new_n894), .ZN(G63));
  NAND2_X1  g709(.A1(G217), .A2(G902), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT60), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n854), .A2(new_n622), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n855), .A2(new_n897), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n853), .B(new_n899), .C1(new_n900), .C2(new_n575), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n899), .A2(new_n902), .A3(new_n853), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT61), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n901), .B(new_n904), .ZN(G66));
  NAND2_X1  g719(.A1(new_n812), .A2(new_n293), .ZN(new_n906));
  INV_X1    g720(.A(G224), .ZN(new_n907));
  OAI21_X1  g721(.A(G953), .B1(new_n534), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(KEYINPUT122), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(KEYINPUT122), .B2(new_n906), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n858), .B1(G898), .B2(new_n293), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n910), .B(new_n911), .Z(G69));
  NAND2_X1  g726(.A1(new_n234), .A2(new_n243), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n628), .B2(new_n293), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n641), .A2(new_n665), .A3(new_n692), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n714), .A2(new_n706), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(KEYINPUT126), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n699), .A2(new_n686), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n731), .A2(KEYINPUT125), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT125), .B1(new_n731), .B2(new_n921), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n744), .B(new_n754), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n919), .B(new_n924), .C1(KEYINPUT126), .C2(new_n918), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n916), .B1(new_n925), .B2(new_n293), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n915), .B(KEYINPUT123), .Z(new_n927));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n917), .A2(new_n662), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n809), .B1(new_n800), .B2(new_n802), .ZN(new_n930));
  NOR4_X1   g744(.A1(new_n930), .A2(new_n676), .A3(new_n646), .A4(new_n752), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT124), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n744), .A2(new_n754), .A3(new_n929), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n928), .B1(new_n917), .B2(new_n662), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n927), .B1(new_n935), .B2(new_n293), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n926), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n927), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n293), .B1(G227), .B2(G900), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n937), .B(new_n941), .ZN(G72));
  NAND2_X1  g756(.A1(G472), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT63), .Z(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n935), .B2(new_n812), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n649), .ZN(new_n946));
  INV_X1    g760(.A(new_n944), .ZN(new_n947));
  INV_X1    g761(.A(new_n812), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n925), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n247), .A2(new_n253), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n853), .B(new_n946), .C1(new_n949), .C2(new_n951), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n829), .A2(new_n837), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n649), .A2(new_n950), .A3(new_n947), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(G57));
endmodule


