//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0007(.A(G97), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  AND2_X1   g0012(.A1(KEYINPUT65), .A2(G68), .ZN(new_n213));
  NOR2_X1   g0013(.A1(KEYINPUT65), .A2(G68), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  OAI21_X1  g0023(.A(new_n212), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n203), .A2(new_n205), .ZN(new_n227));
  INV_X1    g0027(.A(G50), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n212), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT0), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n233), .B(new_n236), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n226), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n201), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT68), .B(G50), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n252), .B(new_n253), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  OAI21_X1  g0055(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n231), .A2(G33), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n256), .B1(new_n257), .B2(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT70), .B1(new_n212), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT70), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n265), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n230), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n262), .A2(new_n267), .B1(new_n228), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n267), .A2(new_n270), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n272), .B(G50), .C1(G1), .C2(new_n231), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT9), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n280), .A3(G274), .ZN(new_n281));
  INV_X1    g0081(.A(G226), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G1698), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n289), .A2(G222), .B1(G77), .B2(new_n288), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n263), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G1698), .ZN(new_n295));
  XOR2_X1   g0095(.A(KEYINPUT69), .B(G223), .Z(new_n296));
  OAI21_X1  g0096(.A(new_n290), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n280), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n285), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(G190), .B2(new_n299), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n275), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT10), .B1(new_n302), .B2(KEYINPUT74), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n274), .B(new_n308), .C1(G169), .C2(new_n299), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT73), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT72), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n269), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n268), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n310), .B1(new_n315), .B2(new_n267), .ZN(new_n316));
  INV_X1    g0116(.A(new_n267), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(KEYINPUT73), .A3(new_n314), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n316), .A2(new_n318), .B1(new_n268), .B2(G20), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G77), .ZN(new_n320));
  INV_X1    g0120(.A(G77), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n261), .A2(new_n259), .B1(new_n231), .B2(new_n321), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n260), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n267), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT71), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n320), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G244), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n281), .B1(new_n330), .B2(new_n284), .ZN(new_n331));
  INV_X1    g0131(.A(G238), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G1698), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G232), .B2(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n294), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n280), .B1(new_n288), .B2(new_n209), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n300), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(G190), .B2(new_n337), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n329), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n337), .A2(G169), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n307), .B2(new_n337), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n328), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n305), .A2(new_n306), .A3(new_n309), .A4(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n216), .A2(new_n231), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n259), .A2(new_n228), .B1(new_n260), .B2(new_n321), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n267), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT11), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n319), .A2(G68), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT12), .B1(new_n270), .B2(new_n202), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n215), .A2(KEYINPUT12), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n315), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n357));
  INV_X1    g0157(.A(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n282), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n240), .A2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n286), .C2(new_n287), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT75), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(KEYINPUT75), .A3(new_n362), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(new_n298), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT13), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n281), .B1(new_n332), .B2(new_n284), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n368), .B1(new_n367), .B2(new_n370), .ZN(new_n372));
  OAI211_X1 g0172(.A(G169), .B(new_n357), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n361), .A2(KEYINPUT75), .A3(new_n362), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT75), .B1(new_n361), .B2(new_n362), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n374), .A2(new_n375), .A3(new_n280), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT13), .B1(new_n376), .B2(new_n369), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(G179), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n378), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n357), .B1(new_n381), .B2(G169), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n356), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n356), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(G200), .ZN(new_n385));
  INV_X1    g0185(.A(G190), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n384), .B(new_n385), .C1(new_n386), .C2(new_n381), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n261), .B1(new_n268), .B2(G20), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n272), .A2(new_n389), .B1(new_n270), .B2(new_n261), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(KEYINPUT65), .A2(G68), .ZN(new_n392));
  NAND2_X1  g0192(.A1(KEYINPUT65), .A2(G68), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n201), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n394), .B2(new_n227), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n259), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n292), .A2(new_n231), .A3(new_n293), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n231), .A4(new_n293), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n202), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n317), .B1(new_n405), .B2(KEYINPUT16), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n215), .B1(new_n402), .B2(new_n403), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n407), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n391), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G169), .ZN(new_n411));
  OR2_X1    g0211(.A1(G223), .A2(G1698), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n282), .A2(G1698), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n413), .C1(new_n286), .C2(new_n287), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n298), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n280), .A2(G232), .A3(new_n283), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n281), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n411), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n280), .B1(new_n414), .B2(new_n415), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n422), .A2(new_n419), .A3(new_n307), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT18), .B1(new_n410), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(G58), .B1(new_n213), .B2(new_n214), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(new_n205), .A3(new_n203), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n397), .B1(new_n427), .B2(G20), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n288), .B2(new_n231), .ZN(new_n429));
  INV_X1    g0229(.A(new_n403), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n431), .A3(KEYINPUT16), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n409), .A2(new_n432), .A3(new_n267), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n424), .B1(new_n433), .B2(new_n390), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n417), .A2(new_n420), .A3(new_n386), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n300), .B1(new_n422), .B2(new_n419), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n433), .A2(new_n390), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n433), .A2(KEYINPUT17), .A3(new_n390), .A4(new_n439), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n425), .A2(new_n436), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n347), .A2(new_n388), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(G116), .B1(new_n263), .B2(G1), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n316), .B2(new_n318), .ZN(new_n447));
  AOI21_X1  g0247(.A(G20), .B1(G33), .B2(G283), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n263), .A2(G97), .ZN(new_n449));
  INV_X1    g0249(.A(G116), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n448), .A2(new_n449), .B1(G20), .B2(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n267), .A2(KEYINPUT20), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT20), .B1(new_n267), .B2(new_n451), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n452), .A2(new_n453), .B1(G116), .B2(new_n314), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n294), .A2(G264), .A3(G1698), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n294), .A2(G257), .A3(new_n358), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n288), .A2(G303), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT82), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT82), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n456), .A2(new_n457), .A3(new_n461), .A4(new_n458), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n298), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT5), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT77), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(G41), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n276), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n277), .A2(G1), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n280), .A2(G274), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G270), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n280), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n411), .B1(new_n463), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT21), .B1(new_n455), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n280), .B1(new_n459), .B2(KEYINPUT82), .ZN(new_n479));
  AOI211_X1 g0279(.A(new_n386), .B(new_n475), .C1(new_n479), .C2(new_n462), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n300), .B1(new_n463), .B2(new_n476), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n455), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n475), .B1(new_n479), .B2(new_n462), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n477), .A2(KEYINPUT21), .B1(G179), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n455), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT83), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT83), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT21), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n483), .A2(new_n488), .A3(new_n411), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n307), .B(new_n475), .C1(new_n479), .C2(new_n462), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n487), .B(new_n455), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  AOI211_X1 g0291(.A(new_n478), .B(new_n482), .C1(new_n486), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n473), .A2(G257), .A3(new_n280), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n471), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G250), .A2(G1698), .ZN(new_n495));
  NAND2_X1  g0295(.A1(KEYINPUT4), .A2(G244), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(G1698), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n294), .A2(new_n497), .B1(G33), .B2(G283), .ZN(new_n498));
  OAI211_X1 g0298(.A(G244), .B(new_n358), .C1(new_n286), .C2(new_n287), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n298), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n386), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n280), .B1(new_n498), .B2(new_n501), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n471), .A2(new_n493), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n300), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT6), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n511), .A2(new_n208), .A3(G107), .ZN(new_n512));
  XNOR2_X1  g0312(.A(G97), .B(G107), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n514), .A2(new_n231), .B1(new_n321), .B2(new_n259), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n209), .B1(new_n402), .B2(new_n403), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n267), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n269), .A2(G97), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n263), .A2(G1), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n267), .A2(new_n270), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n518), .B1(new_n520), .B2(G97), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n510), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n494), .A2(new_n503), .A3(G179), .ZN(new_n525));
  OAI21_X1  g0325(.A(G169), .B1(new_n506), .B2(new_n507), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT78), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n522), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n527), .B2(new_n522), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n524), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT79), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n524), .B(KEYINPUT79), .C1(new_n530), .C2(new_n531), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n294), .A2(G257), .A3(G1698), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G294), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT86), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n289), .B2(G250), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n294), .A2(G250), .A3(new_n358), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n539), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n298), .ZN(new_n545));
  INV_X1    g0345(.A(new_n474), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G264), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n307), .A3(new_n471), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n289), .A2(new_n540), .A3(G250), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n538), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n471), .B(new_n547), .C1(new_n551), .C2(new_n280), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n411), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n231), .A2(G107), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT23), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT85), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT85), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n557), .B(KEYINPUT23), .C1(new_n231), .C2(G107), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n556), .A2(new_n558), .B1(new_n555), .B2(new_n554), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n560), .B(KEYINPUT84), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n231), .B(G87), .C1(new_n286), .C2(new_n287), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n563), .B(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT24), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n563), .B(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT24), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n561), .A4(new_n559), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n317), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n269), .A2(G107), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT25), .ZN(new_n572));
  INV_X1    g0372(.A(new_n520), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(new_n209), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n548), .B(new_n553), .C1(new_n570), .C2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n570), .A2(new_n574), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n552), .A2(new_n300), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n552), .A2(G190), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(G1698), .C1(new_n286), .C2(new_n287), .ZN(new_n580));
  OAI211_X1 g0380(.A(G238), .B(new_n358), .C1(new_n286), .C2(new_n287), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n263), .C2(new_n450), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n298), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n280), .A2(G274), .A3(new_n468), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n268), .A2(G45), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n280), .A2(G250), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT80), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n584), .A2(new_n586), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT80), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n583), .A2(new_n307), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT81), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n588), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n587), .B1(new_n584), .B2(new_n586), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(KEYINPUT81), .A3(new_n307), .A4(new_n583), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n583), .A2(new_n588), .A3(new_n590), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n411), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n294), .A2(new_n231), .A3(G68), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT19), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n231), .B1(new_n362), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G87), .B2(new_n210), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n260), .B2(new_n208), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n267), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n315), .A2(new_n324), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n573), .C2(new_n324), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n593), .A2(new_n597), .A3(new_n599), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n520), .A2(G87), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n610), .A2(new_n606), .A3(new_n607), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n596), .A2(G190), .A3(new_n583), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n583), .A2(new_n588), .A3(new_n590), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n611), .B(new_n612), .C1(new_n300), .C2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n535), .A2(new_n575), .A3(new_n579), .A4(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n445), .A2(new_n492), .A3(new_n534), .A4(new_n616), .ZN(G372));
  AND2_X1   g0417(.A1(new_n305), .A2(new_n306), .ZN(new_n618));
  AOI211_X1 g0418(.A(KEYINPUT18), .B(new_n424), .C1(new_n433), .C2(new_n390), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n433), .A2(new_n390), .ZN(new_n620));
  INV_X1    g0420(.A(new_n424), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n435), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n442), .A2(new_n443), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n387), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n383), .B2(new_n344), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n618), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(new_n309), .ZN(new_n629));
  INV_X1    g0429(.A(new_n445), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n527), .A2(new_n522), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT78), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(new_n529), .B1(new_n523), .B2(new_n510), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n455), .B1(new_n489), .B2(new_n490), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n455), .A2(new_n477), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n488), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n636), .A3(new_n575), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n611), .A2(new_n612), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n594), .B2(new_n595), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n590), .A2(KEYINPUT88), .A3(new_n588), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT87), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n582), .A2(new_n643), .A3(new_n298), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n583), .A2(KEYINPUT87), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G200), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n411), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n608), .A2(new_n591), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n638), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n633), .A2(new_n637), .A3(new_n579), .A4(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n632), .A2(new_n529), .A3(new_n614), .A4(new_n609), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n527), .A2(KEYINPUT89), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT89), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n525), .B2(new_n526), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n654), .A2(new_n523), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n647), .A2(new_n638), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n649), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n653), .A2(new_n661), .A3(new_n659), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n651), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n629), .B1(new_n630), .B2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n268), .A2(new_n231), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n570), .B2(new_n574), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n579), .A2(new_n575), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n672), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n548), .A2(new_n553), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT92), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n674), .A2(KEYINPUT92), .A3(new_n675), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n486), .A2(new_n491), .ZN(new_n680));
  INV_X1    g0480(.A(new_n482), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n455), .A2(new_n671), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n680), .A2(new_n636), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n477), .A2(KEYINPUT21), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n483), .A2(G179), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n455), .B(new_n671), .C1(new_n686), .C2(new_n478), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT90), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT91), .B1(new_n689), .B2(G330), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n688), .A2(KEYINPUT90), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT90), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n683), .B2(new_n687), .ZN(new_n693));
  OAI211_X1 g0493(.A(KEYINPUT91), .B(G330), .C1(new_n691), .C2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n679), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n671), .B1(new_n680), .B2(new_n636), .ZN(new_n697));
  INV_X1    g0497(.A(new_n575), .ZN(new_n698));
  INV_X1    g0498(.A(new_n671), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n679), .A2(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(new_n700), .ZN(G399));
  NAND3_X1  g0501(.A1(new_n234), .A2(KEYINPUT93), .A3(new_n276), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT93), .B1(new_n234), .B2(new_n276), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n210), .A2(G87), .A3(G116), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n229), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n706), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n616), .A2(new_n492), .A3(new_n534), .A4(new_n699), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n483), .A2(G179), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n646), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT94), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n552), .A2(new_n716), .A3(new_n504), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n552), .B2(new_n504), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n545), .A2(new_n613), .A3(new_n508), .A4(new_n547), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n685), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n544), .A2(new_n298), .B1(G264), .B2(new_n546), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n504), .A2(new_n598), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n490), .A2(KEYINPUT30), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(KEYINPUT31), .B(new_n671), .C1(new_n719), .C2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n552), .A2(new_n504), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT94), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n552), .A2(new_n716), .A3(new_n504), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n646), .A3(new_n731), .A4(new_n714), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n722), .A3(new_n725), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT31), .B1(new_n733), .B2(new_n671), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n712), .B1(new_n713), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n663), .A2(new_n699), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT29), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n487), .B1(new_n686), .B2(new_n455), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n484), .A2(KEYINPUT83), .A3(new_n485), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n636), .B(new_n575), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n650), .A2(new_n633), .A3(new_n579), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n660), .B1(new_n650), .B2(new_n657), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n659), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n671), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT29), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n736), .B1(new_n739), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n711), .B1(new_n750), .B2(G1), .ZN(G364));
  NOR2_X1   g0551(.A1(new_n689), .A2(G330), .ZN(new_n752));
  INV_X1    g0552(.A(G13), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n268), .B1(new_n754), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n705), .A2(new_n756), .ZN(new_n757));
  OR4_X1    g0557(.A1(new_n690), .A2(new_n752), .A3(new_n695), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n294), .A2(new_n234), .ZN(new_n759));
  INV_X1    g0559(.A(G355), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n759), .A2(new_n760), .B1(G116), .B2(new_n234), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n251), .A2(G45), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n288), .A2(new_n234), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT95), .Z(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n277), .B2(new_n229), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n761), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n230), .B1(G20), .B2(new_n411), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n773), .A2(new_n705), .A3(new_n756), .ZN(new_n774));
  INV_X1    g0574(.A(new_n770), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n231), .B1(new_n776), .B2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n208), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n231), .A2(G190), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n776), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G159), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n778), .B1(new_n782), .B2(KEYINPUT32), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(KEYINPUT32), .B2(new_n782), .ZN(new_n784));
  NAND3_X1  g0584(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n300), .A2(G179), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT97), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n779), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n294), .B1(new_n202), .B2(new_n787), .C1(new_n790), .C2(new_n209), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n231), .A2(new_n386), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n784), .B(new_n791), .C1(G87), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n307), .A2(G200), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n779), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G58), .A2(new_n798), .B1(new_n800), .B2(G77), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n785), .A2(new_n386), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n801), .B1(new_n228), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT96), .ZN(new_n805));
  INV_X1    g0605(.A(G303), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n793), .A2(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G311), .A2(new_n800), .B1(new_n781), .B2(G329), .ZN(new_n808));
  INV_X1    g0608(.A(G322), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n808), .B(new_n288), .C1(new_n809), .C2(new_n797), .ZN(new_n810));
  INV_X1    g0610(.A(new_n790), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n807), .B(new_n810), .C1(G283), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G294), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n777), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(KEYINPUT33), .A2(G317), .ZN(new_n815));
  NAND2_X1  g0615(.A1(KEYINPUT33), .A2(G317), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n787), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n814), .B(new_n817), .C1(G326), .C2(new_n802), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n795), .A2(new_n805), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n769), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n774), .B1(new_n775), .B2(new_n819), .C1(new_n689), .C2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n758), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  INV_X1    g0623(.A(KEYINPUT100), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n344), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n328), .A2(new_n671), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n328), .A2(KEYINPUT100), .A3(new_n343), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n825), .A2(new_n340), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n345), .A2(new_n671), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT101), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n737), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n825), .A2(new_n827), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n341), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n699), .B(new_n834), .C1(new_n651), .C2(new_n662), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n736), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n757), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n775), .A2(new_n768), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n757), .B1(G77), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT98), .Z(new_n842));
  AOI22_X1  g0642(.A1(G143), .A2(new_n798), .B1(new_n800), .B2(G159), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n803), .B2(new_n844), .C1(new_n257), .C2(new_n787), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT34), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n790), .A2(new_n202), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n793), .A2(new_n228), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n294), .B1(new_n777), .B2(new_n201), .C1(new_n850), .C2(new_n780), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n845), .A2(new_n846), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n803), .A2(new_n806), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n778), .B(new_n854), .C1(G283), .C2(new_n786), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n793), .A2(new_n209), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G116), .A2(new_n800), .B1(new_n781), .B2(G311), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n857), .B(new_n288), .C1(new_n813), .C2(new_n797), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n856), .B(new_n858), .C1(G87), .C2(new_n811), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n852), .A2(new_n853), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n842), .B1(new_n860), .B2(new_n775), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT99), .Z(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n768), .B2(new_n830), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n839), .A2(new_n863), .ZN(G384));
  NOR2_X1   g0664(.A1(new_n754), .A2(new_n268), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n669), .B1(new_n433), .B2(new_n390), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n867), .B2(KEYINPUT103), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n434), .ZN(new_n870));
  INV_X1    g0670(.A(new_n669), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n620), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n872), .A3(new_n440), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n433), .A2(new_n390), .A3(new_n439), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(new_n434), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n868), .B1(new_n876), .B2(new_n872), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n866), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n444), .A2(new_n867), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n869), .A2(new_n873), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n868), .A3(new_n872), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT104), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n407), .B1(new_n399), .B2(new_n404), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(new_n432), .A3(new_n267), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n669), .B1(new_n887), .B2(new_n390), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n444), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n870), .A2(new_n872), .A3(new_n890), .A4(new_n440), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n424), .B1(new_n887), .B2(new_n390), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n875), .A2(new_n892), .A3(new_n888), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n893), .B2(new_n890), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n356), .A2(new_n671), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n383), .A2(new_n387), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n383), .B2(new_n387), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n830), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n713), .B2(new_n735), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(KEYINPUT40), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n895), .A2(KEYINPUT102), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT102), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n889), .A2(new_n894), .A3(new_n906), .A4(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n887), .A2(new_n390), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n871), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n623), .B2(new_n625), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n621), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n909), .A2(new_n911), .A3(new_n440), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n912), .A2(KEYINPUT37), .B1(new_n876), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n884), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n905), .A2(new_n907), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n897), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n388), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n383), .A2(new_n387), .A3(new_n897), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n918), .A2(new_n919), .B1(new_n829), .B2(new_n828), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n579), .A2(new_n615), .A3(new_n575), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n921), .A2(new_n534), .A3(new_n535), .A4(new_n699), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n680), .A2(new_n636), .A3(new_n681), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n671), .B1(new_n719), .B2(new_n726), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT31), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n727), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n920), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n904), .B1(new_n916), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT105), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n905), .A2(new_n907), .A3(new_n915), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n901), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT105), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n934), .A3(new_n904), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n903), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT106), .Z(new_n937));
  NAND2_X1  g0737(.A1(new_n713), .A2(new_n735), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n445), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n939), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(G330), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n383), .A2(new_n671), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT39), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT38), .B1(new_n889), .B2(new_n894), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(KEYINPUT102), .B2(new_n895), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n947), .B2(new_n907), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n910), .A2(new_n914), .A3(new_n884), .ZN(new_n949));
  AOI211_X1 g0749(.A(KEYINPUT39), .B(new_n949), .C1(new_n883), .C2(new_n884), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n944), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n898), .A2(new_n899), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n671), .B1(new_n825), .B2(new_n827), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n952), .B1(new_n835), .B2(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n955), .A2(new_n932), .B1(new_n624), .B2(new_n669), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n739), .A2(new_n445), .A3(new_n749), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n629), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n957), .B(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n865), .B1(new_n942), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n960), .B2(new_n942), .ZN(new_n962));
  INV_X1    g0762(.A(new_n514), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT35), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT35), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n964), .A2(G116), .A3(new_n232), .A4(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT36), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n229), .A2(G77), .A3(new_n426), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(G50), .B2(new_n202), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(G1), .A3(new_n753), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(new_n967), .A3(new_n970), .ZN(G367));
  OAI221_X1 g0771(.A(new_n771), .B1(new_n234), .B2(new_n324), .C1(new_n764), .C2(new_n246), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n757), .ZN(new_n973));
  INV_X1    g0773(.A(new_n650), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n611), .A2(new_n699), .ZN(new_n975));
  MUX2_X1   g0775(.A(new_n974), .B(new_n659), .S(new_n975), .Z(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n797), .A2(new_n257), .B1(new_n799), .B2(new_n228), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n288), .B(new_n978), .C1(G137), .C2(new_n781), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n777), .A2(new_n202), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n787), .A2(new_n396), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(G143), .C2(new_n802), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n811), .A2(G77), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n794), .A2(G58), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n979), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n793), .A2(new_n450), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT46), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n811), .A2(G97), .ZN(new_n988));
  INV_X1    g0788(.A(G311), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n787), .A2(new_n813), .B1(new_n803), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n777), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n990), .B1(G107), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n294), .B1(new_n798), .B2(G303), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G283), .A2(new_n800), .B1(new_n781), .B2(G317), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n988), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n985), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT109), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  OAI221_X1 g0798(.A(new_n973), .B1(new_n977), .B2(new_n820), .C1(new_n775), .C2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT110), .Z(new_n1000));
  INV_X1    g0800(.A(new_n697), .ZN(new_n1001));
  OAI21_X1  g0801(.A(G330), .B1(new_n691), .B2(new_n693), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT91), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n679), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n1004), .A2(new_n694), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(new_n1004), .B2(new_n694), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n694), .A3(new_n1005), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n696), .A2(new_n697), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT45), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n698), .A2(new_n699), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n1005), .B2(new_n1001), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n633), .B1(new_n523), .B2(new_n699), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n657), .A2(new_n671), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1012), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n1017), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1014), .A2(KEYINPUT44), .A3(new_n1018), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT44), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n700), .B2(new_n1017), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n696), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n1007), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n750), .B1(new_n1011), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n705), .B(new_n1031), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n756), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1017), .A2(new_n698), .B1(new_n529), .B2(new_n632), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT107), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n671), .B1(new_n1035), .B2(KEYINPUT107), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n679), .A2(new_n697), .A3(new_n1017), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1036), .A2(new_n1037), .B1(new_n1038), .B2(KEYINPUT42), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(KEYINPUT42), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1039), .A2(new_n1040), .B1(KEYINPUT43), .B2(new_n977), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT43), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n976), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1041), .B(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1007), .A2(new_n1017), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1000), .B1(new_n1034), .B2(new_n1046), .ZN(G387));
  INV_X1    g0847(.A(new_n750), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1006), .A2(new_n1007), .A3(new_n1001), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n697), .B1(new_n696), .B2(new_n1009), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1008), .A2(new_n1010), .A3(new_n750), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n705), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1008), .A2(new_n1010), .A3(new_n756), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n759), .A2(new_n707), .B1(G107), .B2(new_n234), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n243), .A2(new_n277), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n261), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n228), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT50), .Z(new_n1059));
  INV_X1    g0859(.A(new_n707), .ZN(new_n1060));
  AOI211_X1 g0860(.A(G45), .B(new_n1060), .C1(G68), .C2(G77), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n764), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1055), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n757), .B1(new_n1063), .B2(new_n772), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n797), .A2(new_n228), .B1(new_n780), .B2(new_n257), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n288), .B(new_n1065), .C1(G68), .C2(new_n800), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n396), .A2(new_n803), .B1(new_n787), .B2(new_n261), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n777), .A2(new_n324), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n794), .A2(G77), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1066), .A2(new_n988), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n294), .B1(new_n781), .B2(G326), .ZN(new_n1072));
  INV_X1    g0872(.A(G283), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n793), .A2(new_n813), .B1(new_n1073), .B2(new_n777), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G317), .A2(new_n798), .B1(new_n800), .B2(G303), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n803), .B2(new_n809), .C1(new_n989), .C2(new_n787), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1072), .B1(new_n450), .B2(new_n790), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1071), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1064), .B1(new_n1083), .B2(new_n770), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n679), .B2(new_n820), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1054), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1053), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT111), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1053), .A2(new_n1086), .A3(KEYINPUT111), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(G393));
  INV_X1    g0891(.A(new_n1029), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n756), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n254), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n771), .B1(new_n208), .B2(new_n234), .C1(new_n1094), .C2(new_n764), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n757), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n288), .B1(new_n780), .B2(new_n809), .C1(new_n813), .C2(new_n799), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n798), .A2(G311), .B1(G317), .B2(new_n802), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1098), .B(new_n1099), .Z(new_n1100));
  OAI22_X1  g0900(.A1(new_n787), .A2(new_n806), .B1(new_n777), .B2(new_n450), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n209), .A2(new_n790), .B1(new_n793), .B2(new_n1073), .ZN(new_n1102));
  OR4_X1    g0902(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G87), .A2(new_n811), .B1(new_n794), .B2(new_n216), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n294), .B1(new_n799), .B2(new_n261), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n787), .A2(new_n228), .B1(new_n777), .B2(new_n321), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G143), .C2(new_n781), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n803), .A2(new_n257), .B1(new_n797), .B2(new_n396), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1109));
  XNOR2_X1  g0909(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1104), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1103), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1096), .B1(new_n1112), .B2(new_n770), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT114), .Z(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1017), .B2(new_n820), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1052), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(new_n1092), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n705), .B1(new_n1052), .B2(new_n1029), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1093), .B(new_n1115), .C1(new_n1117), .C2(new_n1118), .ZN(G390));
  NAND3_X1  g0919(.A1(new_n885), .A2(new_n945), .A3(new_n895), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n932), .A2(KEYINPUT39), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n767), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n757), .B1(new_n1057), .B2(new_n840), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n848), .B1(G294), .B2(new_n781), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT118), .Z(new_n1125));
  AOI21_X1  g0925(.A(new_n294), .B1(new_n794), .B2(G87), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT117), .Z(new_n1127));
  OAI22_X1  g0927(.A1(new_n797), .A2(new_n450), .B1(new_n799), .B2(new_n208), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n787), .A2(new_n209), .B1(new_n803), .B2(new_n1073), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(G77), .C2(new_n991), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1131), .A2(KEYINPUT119), .ZN(new_n1132));
  INV_X1    g0932(.A(G125), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n294), .B1(new_n780), .B2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n797), .A2(new_n850), .B1(new_n799), .B2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(new_n811), .C2(G50), .ZN(new_n1137));
  INV_X1    g0937(.A(G128), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n803), .A2(new_n1138), .B1(new_n777), .B2(new_n396), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G137), .B2(new_n786), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT53), .B1(new_n793), .B2(new_n257), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n793), .A2(KEYINPUT53), .A3(new_n257), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1137), .A2(new_n1140), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1131), .A2(KEYINPUT119), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1132), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1123), .B1(new_n1145), .B2(new_n770), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1122), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n953), .B1(new_n748), .B2(new_n834), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n943), .B(new_n896), .C1(new_n1148), .C2(new_n952), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1120), .B(new_n1121), .C1(new_n955), .C2(new_n944), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n952), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n938), .A2(G330), .A3(new_n830), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT115), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1149), .A2(new_n1150), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1147), .B1(new_n1157), .B2(new_n755), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT116), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n830), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n712), .B(new_n1160), .C1(new_n713), .C2(new_n735), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1159), .B1(new_n1161), .B2(new_n1151), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n736), .A2(new_n830), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1163), .A2(KEYINPUT116), .A3(new_n952), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1164), .A3(new_n1152), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n835), .A2(new_n954), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1152), .A2(new_n1148), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n831), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1151), .B1(new_n1169), .B2(new_n736), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n958), .B(new_n629), .C1(new_n630), .C2(new_n837), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n706), .B1(new_n1176), .B2(new_n1157), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1171), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(new_n1174), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n1156), .B2(new_n1155), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1158), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(G378));
  NAND2_X1  g0982(.A1(new_n618), .A2(new_n309), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n274), .A2(new_n871), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT120), .Z(new_n1185));
  XNOR2_X1  g0985(.A(new_n1183), .B(new_n1185), .ZN(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n957), .B1(new_n936), .B2(G330), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n934), .B1(new_n933), .B2(new_n904), .ZN(new_n1191));
  AOI211_X1 g0991(.A(KEYINPUT105), .B(KEYINPUT40), .C1(new_n901), .C2(new_n932), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G330), .B(new_n902), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n956), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n943), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1189), .B1(new_n1190), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n931), .A2(new_n935), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1200), .A2(new_n957), .A3(G330), .A4(new_n902), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1201), .A3(new_n1188), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1175), .B1(new_n1157), .B2(new_n1178), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1198), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT57), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n706), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1199), .A2(new_n1201), .A3(new_n1188), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1188), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT121), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(KEYINPUT57), .A4(new_n1203), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1198), .A2(new_n1203), .A3(KEYINPUT57), .A4(new_n1202), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT121), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1206), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n288), .A2(new_n276), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n797), .A2(new_n209), .B1(new_n799), .B2(new_n324), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G283), .C2(new_n781), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n803), .A2(new_n450), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n980), .B(new_n1218), .C1(G97), .C2(new_n786), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n811), .A2(G58), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1217), .A2(new_n1070), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G50), .B1(new_n263), .B2(new_n276), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1221), .A2(new_n1222), .B1(new_n1215), .B2(new_n1223), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n793), .A2(new_n1135), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n786), .A2(G132), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G128), .A2(new_n798), .B1(new_n800), .B2(G137), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n991), .A2(G150), .B1(G125), .B2(new_n802), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n811), .A2(G159), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G33), .B(G41), .C1(new_n781), .C2(G124), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1224), .B1(new_n1222), .B2(new_n1221), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n770), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1236), .B(new_n757), .C1(G50), .C2(new_n840), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1189), .B2(new_n767), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1209), .B2(new_n756), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1214), .A2(new_n1239), .ZN(G375));
  NAND2_X1  g1040(.A1(new_n1178), .A2(new_n1174), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1176), .A2(new_n1033), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n952), .A2(new_n767), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n757), .B1(G68), .B2(new_n840), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n802), .A2(G132), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT122), .Z(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n844), .B2(new_n797), .C1(new_n787), .C2(new_n1135), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT123), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n294), .B1(new_n780), .B2(new_n1138), .C1(new_n257), .C2(new_n799), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1220), .B1(new_n396), .B2(new_n793), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(G50), .C2(new_n991), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1068), .B1(new_n786), .B2(G116), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n813), .B2(new_n803), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n799), .A2(new_n209), .B1(new_n780), .B2(new_n806), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n294), .B(new_n1255), .C1(G283), .C2(new_n798), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n983), .C1(new_n208), .C2(new_n793), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1252), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1244), .B1(new_n1258), .B2(new_n770), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1243), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1178), .B2(new_n755), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1242), .A2(new_n1262), .ZN(G381));
  OR4_X1    g1063(.A1(G384), .A2(G378), .A3(G390), .A4(G381), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1089), .A2(new_n822), .A3(new_n1090), .ZN(new_n1265));
  OR4_X1    g1065(.A1(G387), .A2(new_n1264), .A3(G375), .A4(new_n1265), .ZN(G407));
  NAND2_X1  g1066(.A1(new_n670), .A2(G213), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1181), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G375), .C2(new_n1269), .ZN(G409));
  NAND2_X1  g1070(.A1(new_n1268), .A2(G2897), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1178), .A2(KEYINPUT60), .A3(new_n1174), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1272), .A2(new_n705), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1241), .B1(new_n1179), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G384), .B1(new_n1276), .B2(new_n1262), .ZN(new_n1277));
  INV_X1    g1077(.A(G384), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1278), .B(new_n1261), .C1(new_n1273), .C2(new_n1275), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1271), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1272), .A2(new_n705), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1176), .A2(KEYINPUT60), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n1241), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1278), .B1(new_n1283), .B2(new_n1261), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1276), .A2(G384), .A3(new_n1262), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1284), .A2(G2897), .A3(new_n1268), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT124), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1280), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1280), .B2(new_n1286), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1214), .A2(G378), .A3(new_n1239), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1239), .B1(new_n1032), .B2(new_n1204), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1181), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1268), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(G387), .B(G390), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1093), .A2(new_n1115), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT125), .B1(new_n1300), .B2(G387), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1053), .A2(KEYINPUT111), .A3(new_n1086), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT111), .B1(new_n1053), .B2(new_n1086), .ZN(new_n1304));
  OAI21_X1  g1104(.A(G396), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1305), .A2(new_n1265), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1297), .A2(new_n1302), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1300), .A2(G387), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G390), .B(new_n1000), .C1(new_n1034), .C2(new_n1046), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1265), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1310), .B1(new_n1311), .B2(new_n1301), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1307), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1294), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1315), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1296), .A2(new_n1314), .A3(new_n1318), .A4(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1294), .A2(new_n1321), .A3(new_n1315), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1280), .A2(new_n1286), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1313), .B1(new_n1294), .B2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1321), .B1(new_n1294), .B2(new_n1315), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1322), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1312), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1310), .A2(new_n1311), .A3(new_n1301), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1320), .B1(new_n1326), .B2(new_n1329), .ZN(G405));
  NAND3_X1  g1130(.A1(new_n1284), .A2(KEYINPUT126), .A3(new_n1285), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(KEYINPUT127), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1333), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G375), .A2(new_n1181), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1332), .A2(new_n1307), .A3(new_n1312), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1334), .A2(new_n1291), .A3(new_n1335), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1291), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1336), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1332), .B1(new_n1307), .B2(new_n1312), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1338), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1337), .A2(new_n1341), .ZN(G402));
endmodule


