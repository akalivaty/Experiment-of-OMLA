

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U547 ( .A1(G160), .A2(G40), .ZN(n588) );
  NOR2_X2 U548 ( .A1(G164), .A2(G1384), .ZN(n686) );
  INV_X1 U549 ( .A(n642), .ZN(n627) );
  XNOR2_X1 U550 ( .A(n526), .B(KEYINPUT23), .ZN(n527) );
  AND2_X2 U551 ( .A1(n531), .A2(G2104), .ZN(n866) );
  INV_X1 U552 ( .A(G2105), .ZN(n531) );
  NOR2_X2 U553 ( .A1(n535), .A2(n534), .ZN(G160) );
  NOR2_X1 U554 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U555 ( .A1(KEYINPUT33), .A2(n663), .ZN(n664) );
  NOR2_X1 U556 ( .A1(G543), .A2(G651), .ZN(n767) );
  NAND2_X1 U557 ( .A1(n642), .A2(G1341), .ZN(n512) );
  XOR2_X1 U558 ( .A(KEYINPUT27), .B(n616), .Z(n513) );
  AND2_X1 U559 ( .A1(n726), .A2(n719), .ZN(n514) );
  AND2_X1 U560 ( .A1(n716), .A2(n514), .ZN(n515) );
  AND2_X1 U561 ( .A1(n649), .A2(n648), .ZN(n650) );
  AND2_X1 U562 ( .A1(n717), .A2(n515), .ZN(n718) );
  NOR2_X1 U563 ( .A1(n570), .A2(G651), .ZN(n764) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n518), .Z(n763) );
  NAND2_X1 U565 ( .A1(G91), .A2(n767), .ZN(n517) );
  XOR2_X1 U566 ( .A(KEYINPUT0), .B(G543), .Z(n570) );
  NAND2_X1 U567 ( .A1(G53), .A2(n764), .ZN(n516) );
  NAND2_X1 U568 ( .A1(n517), .A2(n516), .ZN(n521) );
  INV_X1 U569 ( .A(G651), .ZN(n522) );
  NOR2_X1 U570 ( .A1(G543), .A2(n522), .ZN(n518) );
  NAND2_X1 U571 ( .A1(n763), .A2(G65), .ZN(n519) );
  XOR2_X1 U572 ( .A(KEYINPUT70), .B(n519), .Z(n520) );
  NOR2_X1 U573 ( .A1(n521), .A2(n520), .ZN(n525) );
  OR2_X1 U574 ( .A1(n522), .A2(n570), .ZN(n523) );
  XOR2_X1 U575 ( .A(KEYINPUT66), .B(n523), .Z(n768) );
  NAND2_X1 U576 ( .A1(G78), .A2(n768), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(G299) );
  NAND2_X1 U578 ( .A1(G101), .A2(n866), .ZN(n526) );
  XNOR2_X1 U579 ( .A(n527), .B(KEYINPUT65), .ZN(n530) );
  NOR2_X1 U580 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XOR2_X2 U581 ( .A(KEYINPUT17), .B(n528), .Z(n865) );
  NAND2_X1 U582 ( .A1(G137), .A2(n865), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n535) );
  NOR2_X1 U584 ( .A1(G2104), .A2(n531), .ZN(n861) );
  NAND2_X1 U585 ( .A1(G125), .A2(n861), .ZN(n533) );
  AND2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n862) );
  NAND2_X1 U587 ( .A1(G113), .A2(n862), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U589 ( .A1(G138), .A2(n865), .ZN(n537) );
  NAND2_X1 U590 ( .A1(G102), .A2(n866), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G126), .A2(n861), .ZN(n539) );
  NAND2_X1 U593 ( .A1(G114), .A2(n862), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U595 ( .A1(n541), .A2(n540), .ZN(G164) );
  NAND2_X1 U596 ( .A1(G64), .A2(n763), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G52), .A2(n764), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U599 ( .A(KEYINPUT69), .B(n544), .Z(n549) );
  NAND2_X1 U600 ( .A1(n767), .A2(G90), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G77), .A2(n768), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U603 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U604 ( .A1(n549), .A2(n548), .ZN(G171) );
  NAND2_X1 U605 ( .A1(n767), .A2(G89), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G76), .A2(n768), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n553), .B(KEYINPUT5), .ZN(n558) );
  NAND2_X1 U610 ( .A1(G63), .A2(n763), .ZN(n555) );
  NAND2_X1 U611 ( .A1(G51), .A2(n764), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U615 ( .A(n559), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(n767), .A2(G88), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G75), .A2(n768), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G62), .A2(n763), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G50), .A2(n764), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U623 ( .A1(n565), .A2(n564), .ZN(G166) );
  INV_X1 U624 ( .A(G166), .ZN(G303) );
  NAND2_X1 U625 ( .A1(G49), .A2(n764), .ZN(n567) );
  NAND2_X1 U626 ( .A1(G74), .A2(G651), .ZN(n566) );
  NAND2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U628 ( .A(KEYINPUT81), .B(n568), .Z(n569) );
  NOR2_X1 U629 ( .A1(n763), .A2(n569), .ZN(n572) );
  NAND2_X1 U630 ( .A1(n570), .A2(G87), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U632 ( .A1(G86), .A2(n767), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G48), .A2(n764), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n768), .A2(G73), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT2), .B(n575), .Z(n576) );
  NOR2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n763), .A2(G61), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n579), .A2(n578), .ZN(G305) );
  NAND2_X1 U640 ( .A1(G72), .A2(n768), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT67), .B(n580), .Z(n582) );
  NAND2_X1 U642 ( .A1(n767), .A2(G85), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT68), .B(n583), .Z(n587) );
  NAND2_X1 U645 ( .A1(G60), .A2(n763), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G47), .A2(n764), .ZN(n584) );
  AND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U648 ( .A1(n587), .A2(n586), .ZN(G290) );
  NAND2_X2 U649 ( .A1(n588), .A2(n686), .ZN(n642) );
  NAND2_X1 U650 ( .A1(G8), .A2(n642), .ZN(n679) );
  NAND2_X1 U651 ( .A1(n764), .A2(G54), .ZN(n590) );
  NAND2_X1 U652 ( .A1(G79), .A2(n768), .ZN(n589) );
  NAND2_X1 U653 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U654 ( .A1(G92), .A2(n767), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G66), .A2(n763), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U657 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U658 ( .A(n595), .B(KEYINPUT15), .ZN(n897) );
  NAND2_X1 U659 ( .A1(G1348), .A2(n642), .ZN(n597) );
  NAND2_X1 U660 ( .A1(G2067), .A2(n627), .ZN(n596) );
  NAND2_X1 U661 ( .A1(n597), .A2(n596), .ZN(n613) );
  NOR2_X1 U662 ( .A1(n897), .A2(n613), .ZN(n612) );
  XOR2_X1 U663 ( .A(G1996), .B(KEYINPUT97), .Z(n926) );
  NAND2_X1 U664 ( .A1(n627), .A2(n926), .ZN(n598) );
  XNOR2_X1 U665 ( .A(KEYINPUT26), .B(n598), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n599), .A2(n512), .ZN(n610) );
  XOR2_X1 U667 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n601) );
  NAND2_X1 U668 ( .A1(G56), .A2(n763), .ZN(n600) );
  XNOR2_X1 U669 ( .A(n601), .B(n600), .ZN(n607) );
  NAND2_X1 U670 ( .A1(n767), .A2(G81), .ZN(n602) );
  XNOR2_X1 U671 ( .A(n602), .B(KEYINPUT12), .ZN(n604) );
  NAND2_X1 U672 ( .A1(G68), .A2(n768), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U674 ( .A(KEYINPUT13), .B(n605), .Z(n606) );
  NOR2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n764), .A2(G43), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n907) );
  NOR2_X1 U678 ( .A1(n610), .A2(n907), .ZN(n611) );
  NOR2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n615) );
  AND2_X1 U680 ( .A1(n897), .A2(n613), .ZN(n614) );
  NOR2_X1 U681 ( .A1(n615), .A2(n614), .ZN(n620) );
  NAND2_X1 U682 ( .A1(n627), .A2(G2072), .ZN(n616) );
  NAND2_X1 U683 ( .A1(G1956), .A2(n642), .ZN(n617) );
  NAND2_X1 U684 ( .A1(n513), .A2(n617), .ZN(n621) );
  NOR2_X1 U685 ( .A1(G299), .A2(n621), .ZN(n618) );
  XNOR2_X1 U686 ( .A(n618), .B(KEYINPUT98), .ZN(n619) );
  NOR2_X1 U687 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U688 ( .A1(n621), .A2(G299), .ZN(n622) );
  XOR2_X1 U689 ( .A(n622), .B(KEYINPUT28), .Z(n623) );
  XNOR2_X1 U690 ( .A(n625), .B(KEYINPUT29), .ZN(n632) );
  XOR2_X1 U691 ( .A(G2078), .B(KEYINPUT95), .Z(n626) );
  XNOR2_X1 U692 ( .A(KEYINPUT25), .B(n626), .ZN(n927) );
  NAND2_X1 U693 ( .A1(n627), .A2(n927), .ZN(n628) );
  XNOR2_X1 U694 ( .A(n628), .B(KEYINPUT96), .ZN(n630) );
  INV_X1 U695 ( .A(G1961), .ZN(n945) );
  NAND2_X1 U696 ( .A1(n945), .A2(n642), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n630), .A2(n629), .ZN(n636) );
  NAND2_X1 U698 ( .A1(G171), .A2(n636), .ZN(n631) );
  NAND2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n641) );
  NOR2_X1 U700 ( .A1(G1966), .A2(n679), .ZN(n654) );
  NOR2_X1 U701 ( .A1(G2084), .A2(n642), .ZN(n651) );
  NOR2_X1 U702 ( .A1(n654), .A2(n651), .ZN(n633) );
  NAND2_X1 U703 ( .A1(G8), .A2(n633), .ZN(n634) );
  XNOR2_X1 U704 ( .A(KEYINPUT30), .B(n634), .ZN(n635) );
  NOR2_X1 U705 ( .A1(G168), .A2(n635), .ZN(n638) );
  NOR2_X1 U706 ( .A1(G171), .A2(n636), .ZN(n637) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U708 ( .A(KEYINPUT31), .B(n639), .Z(n640) );
  NAND2_X1 U709 ( .A1(n641), .A2(n640), .ZN(n652) );
  NAND2_X1 U710 ( .A1(n652), .A2(G286), .ZN(n649) );
  INV_X1 U711 ( .A(G8), .ZN(n647) );
  NOR2_X1 U712 ( .A1(G1971), .A2(n679), .ZN(n644) );
  NOR2_X1 U713 ( .A1(G2090), .A2(n642), .ZN(n643) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U715 ( .A1(n645), .A2(G303), .ZN(n646) );
  OR2_X1 U716 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n650), .B(KEYINPUT32), .ZN(n658) );
  NAND2_X1 U718 ( .A1(G8), .A2(n651), .ZN(n656) );
  INV_X1 U719 ( .A(n652), .ZN(n653) );
  NOR2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U721 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n658), .A2(n657), .ZN(n672) );
  NOR2_X1 U723 ( .A1(G1976), .A2(G288), .ZN(n665) );
  NOR2_X1 U724 ( .A1(G1971), .A2(G303), .ZN(n659) );
  NOR2_X1 U725 ( .A1(n665), .A2(n659), .ZN(n911) );
  NAND2_X1 U726 ( .A1(n672), .A2(n911), .ZN(n660) );
  NAND2_X1 U727 ( .A1(G1976), .A2(G288), .ZN(n900) );
  NAND2_X1 U728 ( .A1(n660), .A2(n900), .ZN(n661) );
  NOR2_X1 U729 ( .A1(n679), .A2(n661), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n662), .B(KEYINPUT64), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(KEYINPUT99), .ZN(n669) );
  XNOR2_X1 U732 ( .A(G1981), .B(G305), .ZN(n903) );
  NAND2_X1 U733 ( .A1(n665), .A2(KEYINPUT33), .ZN(n666) );
  NOR2_X1 U734 ( .A1(n679), .A2(n666), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n903), .A2(n667), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n684) );
  NOR2_X1 U737 ( .A1(G2090), .A2(G303), .ZN(n670) );
  NAND2_X1 U738 ( .A1(G8), .A2(n670), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n671), .B(KEYINPUT100), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U741 ( .A(KEYINPUT101), .B(n674), .Z(n675) );
  NAND2_X1 U742 ( .A1(n679), .A2(n675), .ZN(n676) );
  XOR2_X1 U743 ( .A(KEYINPUT102), .B(n676), .Z(n682) );
  NOR2_X1 U744 ( .A1(G1981), .A2(G305), .ZN(n677) );
  XOR2_X1 U745 ( .A(n677), .B(KEYINPUT24), .Z(n678) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n680), .B(KEYINPUT94), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n717) );
  NAND2_X1 U750 ( .A1(G160), .A2(G40), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n731) );
  XNOR2_X1 U752 ( .A(G1986), .B(G290), .ZN(n913) );
  NAND2_X1 U753 ( .A1(n731), .A2(n913), .ZN(n716) );
  NAND2_X1 U754 ( .A1(G140), .A2(n865), .ZN(n688) );
  NAND2_X1 U755 ( .A1(G104), .A2(n866), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n690) );
  XOR2_X1 U757 ( .A(KEYINPUT89), .B(KEYINPUT34), .Z(n689) );
  XNOR2_X1 U758 ( .A(n690), .B(n689), .ZN(n695) );
  NAND2_X1 U759 ( .A1(G128), .A2(n861), .ZN(n692) );
  NAND2_X1 U760 ( .A1(G116), .A2(n862), .ZN(n691) );
  NAND2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U762 ( .A(KEYINPUT35), .B(n693), .Z(n694) );
  NOR2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U764 ( .A(n696), .B(KEYINPUT36), .ZN(n697) );
  XNOR2_X1 U765 ( .A(n697), .B(KEYINPUT90), .ZN(n880) );
  XNOR2_X1 U766 ( .A(G2067), .B(KEYINPUT37), .ZN(n728) );
  NOR2_X1 U767 ( .A1(n880), .A2(n728), .ZN(n985) );
  NAND2_X1 U768 ( .A1(n731), .A2(n985), .ZN(n726) );
  NAND2_X1 U769 ( .A1(G131), .A2(n865), .ZN(n699) );
  NAND2_X1 U770 ( .A1(G119), .A2(n861), .ZN(n698) );
  NAND2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U772 ( .A1(G95), .A2(n866), .ZN(n701) );
  NAND2_X1 U773 ( .A1(G107), .A2(n862), .ZN(n700) );
  NAND2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n702) );
  OR2_X1 U775 ( .A1(n703), .A2(n702), .ZN(n879) );
  NAND2_X1 U776 ( .A1(G1991), .A2(n879), .ZN(n704) );
  XOR2_X1 U777 ( .A(KEYINPUT91), .B(n704), .Z(n714) );
  NAND2_X1 U778 ( .A1(G129), .A2(n861), .ZN(n706) );
  NAND2_X1 U779 ( .A1(G117), .A2(n862), .ZN(n705) );
  NAND2_X1 U780 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U781 ( .A1(n866), .A2(G105), .ZN(n707) );
  XOR2_X1 U782 ( .A(KEYINPUT38), .B(n707), .Z(n708) );
  NOR2_X1 U783 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U784 ( .A(n710), .B(KEYINPUT92), .ZN(n712) );
  NAND2_X1 U785 ( .A1(G141), .A2(n865), .ZN(n711) );
  NAND2_X1 U786 ( .A1(n712), .A2(n711), .ZN(n860) );
  NAND2_X1 U787 ( .A1(G1996), .A2(n860), .ZN(n713) );
  NAND2_X1 U788 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U789 ( .A(KEYINPUT93), .B(n715), .Z(n986) );
  NAND2_X1 U790 ( .A1(n731), .A2(n986), .ZN(n719) );
  XNOR2_X1 U791 ( .A(n718), .B(KEYINPUT103), .ZN(n733) );
  NOR2_X1 U792 ( .A1(G1996), .A2(n860), .ZN(n976) );
  INV_X1 U793 ( .A(n719), .ZN(n723) );
  NOR2_X1 U794 ( .A1(G1991), .A2(n879), .ZN(n984) );
  NOR2_X1 U795 ( .A1(G1986), .A2(G290), .ZN(n720) );
  XNOR2_X1 U796 ( .A(KEYINPUT104), .B(n720), .ZN(n721) );
  NOR2_X1 U797 ( .A1(n984), .A2(n721), .ZN(n722) );
  NOR2_X1 U798 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U799 ( .A1(n976), .A2(n724), .ZN(n725) );
  XNOR2_X1 U800 ( .A(KEYINPUT39), .B(n725), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U802 ( .A1(n880), .A2(n728), .ZN(n990) );
  NAND2_X1 U803 ( .A1(n729), .A2(n990), .ZN(n730) );
  NAND2_X1 U804 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U805 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U806 ( .A(n734), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U807 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U808 ( .A(G132), .ZN(G219) );
  INV_X1 U809 ( .A(G82), .ZN(G220) );
  INV_X1 U810 ( .A(G108), .ZN(G238) );
  NAND2_X1 U811 ( .A1(G7), .A2(G661), .ZN(n735) );
  XNOR2_X1 U812 ( .A(n735), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U813 ( .A(G223), .B(KEYINPUT71), .ZN(n814) );
  NAND2_X1 U814 ( .A1(n814), .A2(G567), .ZN(n736) );
  XOR2_X1 U815 ( .A(KEYINPUT11), .B(n736), .Z(G234) );
  XNOR2_X1 U816 ( .A(G860), .B(KEYINPUT73), .ZN(n744) );
  NOR2_X1 U817 ( .A1(n907), .A2(n744), .ZN(n737) );
  XOR2_X1 U818 ( .A(KEYINPUT74), .B(n737), .Z(G153) );
  NAND2_X1 U819 ( .A1(G868), .A2(G171), .ZN(n739) );
  INV_X1 U820 ( .A(n897), .ZN(n884) );
  INV_X1 U821 ( .A(G868), .ZN(n774) );
  NAND2_X1 U822 ( .A1(n884), .A2(n774), .ZN(n738) );
  NAND2_X1 U823 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U824 ( .A(n740), .B(KEYINPUT75), .ZN(G284) );
  XNOR2_X1 U825 ( .A(KEYINPUT76), .B(n774), .ZN(n741) );
  NOR2_X1 U826 ( .A1(G286), .A2(n741), .ZN(n743) );
  NOR2_X1 U827 ( .A1(G868), .A2(G299), .ZN(n742) );
  NOR2_X1 U828 ( .A1(n743), .A2(n742), .ZN(G297) );
  NAND2_X1 U829 ( .A1(G559), .A2(n744), .ZN(n745) );
  XOR2_X1 U830 ( .A(KEYINPUT77), .B(n745), .Z(n746) );
  NAND2_X1 U831 ( .A1(n746), .A2(n884), .ZN(n747) );
  XNOR2_X1 U832 ( .A(n747), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U833 ( .A1(G868), .A2(n907), .ZN(n748) );
  XNOR2_X1 U834 ( .A(KEYINPUT78), .B(n748), .ZN(n751) );
  NAND2_X1 U835 ( .A1(G868), .A2(n884), .ZN(n749) );
  NOR2_X1 U836 ( .A1(G559), .A2(n749), .ZN(n750) );
  NOR2_X1 U837 ( .A1(n751), .A2(n750), .ZN(G282) );
  NAND2_X1 U838 ( .A1(G123), .A2(n861), .ZN(n752) );
  XNOR2_X1 U839 ( .A(n752), .B(KEYINPUT18), .ZN(n759) );
  NAND2_X1 U840 ( .A1(G99), .A2(n866), .ZN(n754) );
  NAND2_X1 U841 ( .A1(G111), .A2(n862), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n757) );
  NAND2_X1 U843 ( .A1(G135), .A2(n865), .ZN(n755) );
  XNOR2_X1 U844 ( .A(KEYINPUT79), .B(n755), .ZN(n756) );
  NOR2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n981) );
  XNOR2_X1 U847 ( .A(G2096), .B(n981), .ZN(n760) );
  NOR2_X1 U848 ( .A1(G2100), .A2(n760), .ZN(n761) );
  XOR2_X1 U849 ( .A(KEYINPUT80), .B(n761), .Z(G156) );
  NAND2_X1 U850 ( .A1(n884), .A2(G559), .ZN(n783) );
  XNOR2_X1 U851 ( .A(n907), .B(n783), .ZN(n762) );
  NOR2_X1 U852 ( .A1(n762), .A2(G860), .ZN(n773) );
  NAND2_X1 U853 ( .A1(G67), .A2(n763), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G55), .A2(n764), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n767), .A2(G93), .ZN(n770) );
  NAND2_X1 U857 ( .A1(G80), .A2(n768), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n775) );
  XNOR2_X1 U860 ( .A(n773), .B(n775), .ZN(G145) );
  NAND2_X1 U861 ( .A1(n774), .A2(n775), .ZN(n786) );
  XNOR2_X1 U862 ( .A(n775), .B(G303), .ZN(n776) );
  XNOR2_X1 U863 ( .A(n776), .B(G299), .ZN(n777) );
  XNOR2_X1 U864 ( .A(KEYINPUT19), .B(n777), .ZN(n779) );
  XNOR2_X1 U865 ( .A(n907), .B(KEYINPUT82), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n779), .B(n778), .ZN(n780) );
  XOR2_X1 U867 ( .A(n780), .B(G305), .Z(n781) );
  XNOR2_X1 U868 ( .A(G288), .B(n781), .ZN(n782) );
  XNOR2_X1 U869 ( .A(G290), .B(n782), .ZN(n883) );
  XNOR2_X1 U870 ( .A(n883), .B(n783), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n784), .A2(G868), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U873 ( .A(n787), .B(KEYINPUT83), .ZN(G295) );
  NAND2_X1 U874 ( .A1(G2078), .A2(G2084), .ZN(n788) );
  XOR2_X1 U875 ( .A(KEYINPUT20), .B(n788), .Z(n789) );
  NAND2_X1 U876 ( .A1(G2090), .A2(n789), .ZN(n790) );
  XNOR2_X1 U877 ( .A(KEYINPUT21), .B(n790), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n791), .A2(G2072), .ZN(n792) );
  XNOR2_X1 U879 ( .A(KEYINPUT84), .B(n792), .ZN(G158) );
  XNOR2_X1 U880 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U881 ( .A1(G120), .A2(G69), .ZN(n793) );
  XNOR2_X1 U882 ( .A(KEYINPUT86), .B(n793), .ZN(n794) );
  NOR2_X1 U883 ( .A1(G238), .A2(n794), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G57), .A2(n795), .ZN(n818) );
  NAND2_X1 U885 ( .A1(n818), .A2(G567), .ZN(n801) );
  NOR2_X1 U886 ( .A1(G220), .A2(G219), .ZN(n796) );
  XNOR2_X1 U887 ( .A(KEYINPUT22), .B(n796), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n797), .A2(G96), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n798), .A2(G218), .ZN(n799) );
  XNOR2_X1 U890 ( .A(n799), .B(KEYINPUT85), .ZN(n819) );
  NAND2_X1 U891 ( .A1(n819), .A2(G2106), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n820) );
  NAND2_X1 U893 ( .A1(G661), .A2(G483), .ZN(n802) );
  XOR2_X1 U894 ( .A(KEYINPUT87), .B(n802), .Z(n803) );
  NOR2_X1 U895 ( .A1(n820), .A2(n803), .ZN(n817) );
  NAND2_X1 U896 ( .A1(G36), .A2(n817), .ZN(n804) );
  XNOR2_X1 U897 ( .A(n804), .B(KEYINPUT88), .ZN(G176) );
  XNOR2_X1 U898 ( .A(G1348), .B(G2454), .ZN(n805) );
  XNOR2_X1 U899 ( .A(n805), .B(G2430), .ZN(n806) );
  XNOR2_X1 U900 ( .A(n806), .B(G1341), .ZN(n812) );
  XOR2_X1 U901 ( .A(G2443), .B(G2427), .Z(n808) );
  XNOR2_X1 U902 ( .A(G2438), .B(G2446), .ZN(n807) );
  XNOR2_X1 U903 ( .A(n808), .B(n807), .ZN(n810) );
  XOR2_X1 U904 ( .A(G2451), .B(G2435), .Z(n809) );
  XNOR2_X1 U905 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U906 ( .A(n812), .B(n811), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n813), .A2(G14), .ZN(n889) );
  XNOR2_X1 U908 ( .A(KEYINPUT105), .B(n889), .ZN(G401) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n814), .ZN(G217) );
  AND2_X1 U910 ( .A1(G15), .A2(G2), .ZN(n815) );
  NAND2_X1 U911 ( .A1(G661), .A2(n815), .ZN(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(G188) );
  XOR2_X1 U914 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  INV_X1 U916 ( .A(G120), .ZN(G236) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  NOR2_X1 U918 ( .A1(n819), .A2(n818), .ZN(G325) );
  INV_X1 U919 ( .A(G325), .ZN(G261) );
  INV_X1 U920 ( .A(n820), .ZN(G319) );
  XNOR2_X1 U921 ( .A(G1991), .B(KEYINPUT41), .ZN(n830) );
  XOR2_X1 U922 ( .A(G1956), .B(G1981), .Z(n822) );
  XNOR2_X1 U923 ( .A(G1996), .B(G1986), .ZN(n821) );
  XNOR2_X1 U924 ( .A(n822), .B(n821), .ZN(n826) );
  XOR2_X1 U925 ( .A(G1961), .B(G1966), .Z(n824) );
  XNOR2_X1 U926 ( .A(G1976), .B(G1971), .ZN(n823) );
  XNOR2_X1 U927 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U928 ( .A(n826), .B(n825), .Z(n828) );
  XNOR2_X1 U929 ( .A(KEYINPUT110), .B(G2474), .ZN(n827) );
  XNOR2_X1 U930 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U931 ( .A(n830), .B(n829), .ZN(G229) );
  XNOR2_X1 U932 ( .A(G2084), .B(G2090), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n831), .B(KEYINPUT42), .ZN(n841) );
  XOR2_X1 U934 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n833) );
  XNOR2_X1 U935 ( .A(KEYINPUT108), .B(G2096), .ZN(n832) );
  XNOR2_X1 U936 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U937 ( .A(G2100), .B(G2072), .Z(n835) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2078), .ZN(n834) );
  XNOR2_X1 U939 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U940 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U941 ( .A(KEYINPUT109), .B(G2678), .ZN(n838) );
  XNOR2_X1 U942 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(G227) );
  NAND2_X1 U944 ( .A1(G124), .A2(n861), .ZN(n842) );
  XOR2_X1 U945 ( .A(KEYINPUT111), .B(n842), .Z(n843) );
  XNOR2_X1 U946 ( .A(n843), .B(KEYINPUT44), .ZN(n845) );
  NAND2_X1 U947 ( .A1(G100), .A2(n866), .ZN(n844) );
  NAND2_X1 U948 ( .A1(n845), .A2(n844), .ZN(n849) );
  NAND2_X1 U949 ( .A1(G136), .A2(n865), .ZN(n847) );
  NAND2_X1 U950 ( .A1(G112), .A2(n862), .ZN(n846) );
  NAND2_X1 U951 ( .A1(n847), .A2(n846), .ZN(n848) );
  NOR2_X1 U952 ( .A1(n849), .A2(n848), .ZN(G162) );
  XNOR2_X1 U953 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n981), .B(KEYINPUT48), .ZN(n850) );
  XNOR2_X1 U955 ( .A(n851), .B(n850), .ZN(n877) );
  NAND2_X1 U956 ( .A1(G139), .A2(n865), .ZN(n853) );
  NAND2_X1 U957 ( .A1(G103), .A2(n866), .ZN(n852) );
  NAND2_X1 U958 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G127), .A2(n861), .ZN(n855) );
  NAND2_X1 U960 ( .A1(G115), .A2(n862), .ZN(n854) );
  NAND2_X1 U961 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U962 ( .A(KEYINPUT47), .B(n856), .Z(n857) );
  NOR2_X1 U963 ( .A1(n858), .A2(n857), .ZN(n969) );
  XOR2_X1 U964 ( .A(n969), .B(G162), .Z(n859) );
  XNOR2_X1 U965 ( .A(n860), .B(n859), .ZN(n873) );
  NAND2_X1 U966 ( .A1(G130), .A2(n861), .ZN(n864) );
  NAND2_X1 U967 ( .A1(G118), .A2(n862), .ZN(n863) );
  NAND2_X1 U968 ( .A1(n864), .A2(n863), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G142), .A2(n865), .ZN(n868) );
  NAND2_X1 U970 ( .A1(G106), .A2(n866), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U972 ( .A(KEYINPUT45), .B(n869), .Z(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(n873), .B(n872), .Z(n875) );
  XNOR2_X1 U975 ( .A(G164), .B(G160), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(n877), .B(n876), .Z(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n881), .B(n880), .ZN(n882) );
  NOR2_X1 U980 ( .A1(G37), .A2(n882), .ZN(G395) );
  INV_X1 U981 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U982 ( .A(n883), .B(KEYINPUT113), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n884), .B(G286), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(G301), .ZN(n888) );
  NOR2_X1 U986 ( .A1(G37), .A2(n888), .ZN(G397) );
  NAND2_X1 U987 ( .A1(G319), .A2(n889), .ZN(n892) );
  NOR2_X1 U988 ( .A1(G229), .A2(G227), .ZN(n890) );
  XNOR2_X1 U989 ( .A(KEYINPUT49), .B(n890), .ZN(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n894) );
  NOR2_X1 U991 ( .A1(G395), .A2(G397), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(G225) );
  INV_X1 U993 ( .A(G225), .ZN(G308) );
  INV_X1 U994 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U995 ( .A(KEYINPUT56), .B(G16), .ZN(n917) );
  XNOR2_X1 U996 ( .A(G1961), .B(G171), .ZN(n896) );
  NAND2_X1 U997 ( .A1(G1971), .A2(G303), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n899) );
  XNOR2_X1 U999 ( .A(G1348), .B(n897), .ZN(n898) );
  NOR2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n906) );
  XOR2_X1 U1002 ( .A(G1966), .B(G168), .Z(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n904), .B(KEYINPUT57), .ZN(n905) );
  NOR2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(n915) );
  XNOR2_X1 U1006 ( .A(n907), .B(G1341), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(G299), .B(G1956), .ZN(n908) );
  NOR2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n1003) );
  XNOR2_X1 U1013 ( .A(G2084), .B(G34), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n918), .B(KEYINPUT54), .ZN(n938) );
  XNOR2_X1 U1015 ( .A(G2090), .B(G35), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n919), .B(KEYINPUT118), .ZN(n935) );
  XOR2_X1 U1017 ( .A(G1991), .B(G25), .Z(n920) );
  NAND2_X1 U1018 ( .A1(G28), .A2(n920), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n921), .B(KEYINPUT119), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(G2067), .B(G26), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(G2072), .B(G33), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n932) );
  XOR2_X1 U1024 ( .A(n926), .B(G32), .Z(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT120), .B(n927), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(G27), .B(n928), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(n933), .B(KEYINPUT53), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(n936), .B(KEYINPUT121), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1033 ( .A(n939), .B(KEYINPUT55), .Z(n940) );
  XNOR2_X1 U1034 ( .A(KEYINPUT122), .B(n940), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(G29), .A2(n941), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT123), .B(n942), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n943), .A2(G11), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n944), .B(KEYINPUT124), .ZN(n1001) );
  XNOR2_X1 U1039 ( .A(G5), .B(n945), .ZN(n958) );
  XNOR2_X1 U1040 ( .A(G1348), .B(KEYINPUT59), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(n946), .B(G4), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G1981), .B(G6), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G19), .B(G1341), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1046 ( .A(KEYINPUT125), .B(G1956), .Z(n951) );
  XNOR2_X1 U1047 ( .A(G20), .B(n951), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1049 ( .A(KEYINPUT60), .B(n954), .Z(n956) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n965) );
  XNOR2_X1 U1053 ( .A(G1976), .B(G23), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n962) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n963), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1060 ( .A(KEYINPUT61), .B(n966), .Z(n967) );
  NOR2_X1 U1061 ( .A1(G16), .A2(n967), .ZN(n968) );
  XOR2_X1 U1062 ( .A(KEYINPUT126), .B(n968), .Z(n999) );
  XNOR2_X1 U1063 ( .A(G2072), .B(n969), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G164), .B(G2078), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n970), .B(KEYINPUT116), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(KEYINPUT50), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(KEYINPUT117), .B(n974), .ZN(n979) );
  XOR2_X1 U1069 ( .A(G2090), .B(G162), .Z(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1071 ( .A(KEYINPUT51), .B(n977), .Z(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n993) );
  XNOR2_X1 U1073 ( .A(G160), .B(G2084), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n980), .B(KEYINPUT114), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(KEYINPUT115), .B(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(KEYINPUT52), .B(n994), .ZN(n996) );
  INV_X1 U1083 ( .A(KEYINPUT55), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1085 ( .A1(n997), .A2(G29), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(n1004), .B(KEYINPUT127), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(KEYINPUT62), .B(n1005), .ZN(G311) );
  INV_X1 U1091 ( .A(G311), .ZN(G150) );
endmodule

