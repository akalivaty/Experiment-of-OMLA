//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT35), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT83), .ZN(new_n204));
  XOR2_X1   g003(.A(G78gat), .B(G106gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT31), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(G50gat), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(KEYINPUT74), .B(KEYINPUT22), .Z(new_n209));
  NAND2_X1  g008(.A1(G211gat), .A2(G218gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G197gat), .B(G204gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G211gat), .ZN(new_n214));
  INV_X1    g013(.A(G218gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n210), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n210), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n211), .A2(new_n218), .A3(new_n212), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n217), .A2(KEYINPUT75), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT75), .B1(new_n217), .B2(new_n219), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G155gat), .ZN(new_n223));
  INV_X1    g022(.A(G162gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G141gat), .ZN(new_n230));
  INV_X1    g029(.A(G141gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G148gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n227), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n228), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G141gat), .B(G148gat), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT79), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n226), .B1(new_n225), .B2(KEYINPUT2), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT79), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n233), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n234), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(KEYINPUT81), .A3(new_n246), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n222), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n217), .A2(new_n219), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n246), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n243), .B1(new_n253), .B2(new_n244), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G228gat), .ZN(new_n256));
  INV_X1    g055(.A(G233gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n251), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n252), .B1(new_n246), .B2(new_n245), .ZN(new_n260));
  OAI22_X1  g059(.A1(new_n254), .A2(new_n260), .B1(new_n256), .B2(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n208), .B1(new_n262), .B2(G22gat), .ZN(new_n263));
  XOR2_X1   g062(.A(KEYINPUT82), .B(G22gat), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n259), .A2(new_n265), .A3(new_n261), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n204), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n264), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n207), .B1(new_n269), .B2(new_n266), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n263), .A2(new_n204), .A3(new_n266), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G15gat), .B(G43gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT69), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(G71gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G99gat), .ZN(new_n277));
  INV_X1    g076(.A(G71gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n275), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G99gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n284));
  OAI21_X1  g083(.A(G120gat), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G120gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(KEYINPUT68), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G127gat), .B(G134gat), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n285), .A2(new_n288), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G113gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n287), .B2(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n292), .A2(new_n295), .B1(new_n299), .B2(new_n290), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n301));
  NAND2_X1  g100(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OR2_X1    g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT24), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n306), .A2(new_n307), .A3(new_n309), .A4(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT64), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n308), .B2(KEYINPUT23), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n315), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n303), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n316), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n307), .B1(new_n305), .B2(KEYINPUT24), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n315), .A2(G169gat), .A3(G176gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n319), .A2(new_n322), .A3(new_n302), .A4(new_n306), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n301), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n308), .A2(KEYINPUT66), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT26), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT26), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n308), .A2(KEYINPUT66), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n307), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT27), .B(G183gat), .ZN(new_n330));
  INV_X1    g129(.A(G190gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(KEYINPUT28), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT28), .B1(new_n330), .B2(new_n331), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n305), .B(new_n329), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n300), .B1(new_n324), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n301), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n309), .A2(new_n307), .A3(new_n311), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n305), .A2(KEYINPUT24), .ZN(new_n340));
  NOR2_X1   g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n302), .B1(new_n343), .B2(new_n319), .ZN(new_n344));
  AND4_X1   g143(.A1(new_n302), .A2(new_n319), .A3(new_n322), .A4(new_n306), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OR2_X1    g145(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n297), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n294), .B1(new_n349), .B2(new_n287), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n350), .A2(new_n296), .A3(new_n291), .A4(new_n289), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n299), .A2(new_n290), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n346), .A2(new_n353), .A3(new_n335), .ZN(new_n354));
  AND2_X1   g153(.A1(G227gat), .A2(G233gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT33), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n282), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(KEYINPUT32), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n358), .B2(new_n360), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n277), .A2(new_n281), .A3(KEYINPUT33), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(KEYINPUT32), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT71), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT34), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n355), .B1(new_n337), .B2(new_n354), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n358), .A2(new_n360), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT70), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT34), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT71), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n365), .B(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n367), .A2(new_n369), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n369), .B1(new_n367), .B2(new_n377), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n203), .B(new_n273), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n239), .A2(new_n242), .ZN(new_n383));
  INV_X1    g182(.A(new_n234), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n353), .A3(new_n245), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(new_n300), .B2(new_n243), .ZN(new_n389));
  AND4_X1   g188(.A1(new_n388), .A2(new_n351), .A3(new_n243), .A4(new_n352), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n382), .B(new_n387), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n382), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n300), .A2(new_n243), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n353), .A2(new_n385), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n381), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT4), .B1(new_n353), .B2(new_n385), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n300), .A2(new_n388), .A3(new_n243), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n352), .A2(new_n351), .B1(new_n243), .B2(new_n244), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n397), .A2(new_n398), .B1(new_n399), .B2(new_n386), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT5), .B1(new_n400), .B2(new_n382), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT0), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G57gat), .ZN(new_n405));
  INV_X1    g204(.A(G85gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(KEYINPUT6), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n381), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n391), .A2(new_n395), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n408), .B(new_n412), .C1(new_n413), .C2(new_n381), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n407), .B1(new_n396), .B2(new_n401), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n409), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n411), .B1(KEYINPUT84), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n324), .A2(new_n336), .ZN(new_n420));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT77), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n246), .B1(new_n324), .B2(new_n336), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n421), .B(KEYINPUT76), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n346), .A2(new_n335), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT77), .ZN(new_n427));
  INV_X1    g226(.A(new_n421), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n222), .ZN(new_n431));
  INV_X1    g230(.A(new_n424), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n423), .A2(new_n421), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n252), .ZN(new_n434));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435));
  INV_X1    g234(.A(G64gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G92gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n431), .A2(new_n434), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT78), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT30), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n431), .A2(new_n434), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n439), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(KEYINPUT78), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n419), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n202), .B1(new_n380), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n273), .B1(new_n378), .B2(new_n379), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT80), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n417), .A2(new_n409), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n441), .A2(KEYINPUT78), .A3(new_n446), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n446), .B1(new_n441), .B2(KEYINPUT78), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(KEYINPUT80), .A3(new_n418), .A4(new_n445), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT35), .B1(new_n451), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n263), .A2(new_n204), .A3(new_n266), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n461), .A2(new_n267), .A3(new_n270), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n363), .A2(KEYINPUT34), .A3(new_n366), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n374), .B1(new_n373), .B2(new_n376), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n463), .A2(new_n464), .B1(KEYINPUT72), .B2(new_n368), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n367), .A2(new_n369), .A3(new_n377), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n419), .A2(new_n448), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT85), .A4(new_n203), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n460), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n431), .A2(new_n434), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n440), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n472), .B2(new_n471), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT38), .ZN(new_n475));
  OAI22_X1  g274(.A1(new_n430), .A2(new_n222), .B1(new_n252), .B2(new_n433), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT38), .B1(new_n476), .B2(KEYINPUT37), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n419), .A2(new_n475), .A3(new_n441), .A4(new_n478), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n400), .A2(new_n382), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n393), .A2(new_n394), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n480), .B(KEYINPUT39), .C1(new_n392), .C2(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n482), .B(new_n407), .C1(KEYINPUT39), .C2(new_n480), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT40), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n414), .A3(new_n448), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n479), .A2(new_n485), .A3(new_n273), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT73), .ZN(new_n487));
  OAI22_X1  g286(.A1(new_n378), .A2(new_n379), .B1(new_n487), .B2(KEYINPUT36), .ZN(new_n488));
  XOR2_X1   g287(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n489));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n466), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n459), .A2(new_n462), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n486), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n470), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G57gat), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n436), .B1(new_n495), .B2(KEYINPUT94), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(G57gat), .A3(G64gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT9), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n499), .A2(G71gat), .A3(G78gat), .ZN(new_n500));
  INV_X1    g299(.A(G78gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n278), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n496), .B(new_n498), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504));
  OAI22_X1  g303(.A1(new_n504), .A2(new_n499), .B1(new_n278), .B2(new_n501), .ZN(new_n505));
  NOR2_X1   g304(.A1(G71gat), .A2(G78gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT93), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT95), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n510), .B(new_n503), .C1(new_n505), .C2(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(KEYINPUT21), .ZN(new_n514));
  XOR2_X1   g313(.A(G127gat), .B(G155gat), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G183gat), .B(G211gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n518), .B(new_n519), .Z(new_n520));
  INV_X1    g319(.A(KEYINPUT97), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n509), .A2(KEYINPUT97), .A3(new_n511), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT21), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(G1gat), .B2(new_n525), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G8gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n520), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(G43gat), .B(G50gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n539), .B1(KEYINPUT87), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n540), .A2(KEYINPUT87), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n544));
  NAND2_X1  g343(.A1(G29gat), .A2(G36gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT14), .ZN(new_n546));
  INV_X1    g345(.A(G29gat), .ZN(new_n547));
  INV_X1    g346(.A(G36gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT88), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n551), .A2(KEYINPUT86), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT86), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n545), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(KEYINPUT15), .B(new_n538), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n553), .A2(new_n541), .A3(new_n545), .A4(new_n542), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT89), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT100), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT101), .ZN(new_n565));
  NAND3_X1  g364(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT7), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n406), .B2(new_n438), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n564), .A2(KEYINPUT7), .A3(new_n566), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT101), .B1(new_n562), .B2(KEYINPUT7), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n567), .B(new_n569), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n564), .A2(KEYINPUT7), .A3(new_n566), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n575), .B(KEYINPUT101), .C1(KEYINPUT7), .C2(new_n562), .ZN(new_n576));
  INV_X1    g375(.A(new_n573), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n576), .A2(new_n577), .A3(new_n567), .A4(new_n569), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n578), .A3(KEYINPUT102), .ZN(new_n579));
  OR3_X1    g378(.A1(new_n572), .A2(KEYINPUT102), .A3(new_n573), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n561), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n554), .A2(KEYINPUT17), .A3(new_n558), .A4(new_n560), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n537), .B(new_n582), .C1(new_n586), .C2(new_n581), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT103), .B(G190gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n215), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n590), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n591), .A2(new_n592), .A3(new_n593), .A4(new_n597), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n536), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n494), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n584), .A2(new_n530), .A3(new_n585), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT90), .B1(new_n561), .B2(new_n529), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n561), .A2(KEYINPUT90), .A3(new_n529), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT18), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G197gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT11), .ZN(new_n615));
  INV_X1    g414(.A(G169gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n607), .A2(new_n606), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n620), .A2(KEYINPUT18), .A3(new_n605), .A4(new_n604), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n605), .B(KEYINPUT13), .Z(new_n622));
  NOR2_X1   g421(.A1(new_n561), .A2(new_n529), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT91), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT91), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n561), .B2(new_n529), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n607), .A2(new_n606), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n622), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n621), .A2(new_n610), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n619), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n621), .A2(new_n610), .A3(new_n629), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n632), .A2(new_n612), .A3(new_n618), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n581), .A2(new_n522), .A3(KEYINPUT10), .A4(new_n523), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n505), .A2(new_n507), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n574), .A2(new_n578), .A3(new_n503), .A4(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n581), .B2(new_n513), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n636), .B1(new_n639), .B2(KEYINPUT10), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  INV_X1    g445(.A(G176gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(G204gat), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n649), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n642), .A2(new_n644), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n635), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n603), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n453), .B(KEYINPUT104), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g459(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n661));
  INV_X1    g460(.A(new_n448), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n665), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n663), .A2(KEYINPUT106), .A3(KEYINPUT42), .A4(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(G8gat), .B1(new_n655), .B2(new_n662), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n666), .B(new_n668), .C1(new_n671), .C2(new_n672), .ZN(G1325gat));
  INV_X1    g472(.A(new_n491), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n656), .A2(G15gat), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n378), .A2(new_n379), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(G15gat), .B1(new_n656), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n675), .A2(new_n678), .ZN(G1326gat));
  NOR2_X1   g478(.A1(new_n655), .A2(new_n273), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT43), .B(G22gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n494), .A2(new_n683), .A3(new_n601), .ZN(new_n684));
  INV_X1    g483(.A(new_n601), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT110), .B(new_n685), .C1(new_n470), .C2(new_n493), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n684), .C1(new_n686), .C2(new_n683), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n494), .A2(new_n601), .ZN(new_n689));
  OAI211_X1 g488(.A(KEYINPUT109), .B(new_n688), .C1(new_n689), .C2(KEYINPUT110), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT111), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n654), .A2(new_n536), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT108), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n691), .A2(new_n692), .A3(new_n658), .A4(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n687), .A2(new_n658), .A3(new_n690), .A4(new_n694), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT111), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(G29gat), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n685), .B1(new_n470), .B2(new_n493), .ZN(new_n699));
  INV_X1    g498(.A(new_n693), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n699), .A2(new_n547), .A3(new_n658), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT107), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n703), .ZN(G1328gat));
  NAND4_X1  g503(.A1(new_n691), .A2(KEYINPUT113), .A3(new_n448), .A4(new_n694), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n687), .A2(new_n448), .A3(new_n690), .A4(new_n694), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT113), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(G36gat), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n689), .A2(new_n693), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n548), .A3(new_n448), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(KEYINPUT46), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n712), .A2(KEYINPUT46), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n709), .A2(new_n715), .ZN(G1329gat));
  NAND4_X1  g515(.A1(new_n687), .A2(new_n674), .A3(new_n690), .A4(new_n694), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n710), .A2(new_n719), .A3(new_n677), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n718), .A2(KEYINPUT47), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1330gat));
  NOR4_X1   g524(.A1(new_n689), .A2(G50gat), .A3(new_n273), .A4(new_n693), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n687), .A2(new_n462), .A3(new_n690), .A4(new_n694), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(G50gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI211_X1 g529(.A(KEYINPUT48), .B(new_n726), .C1(new_n727), .C2(G50gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  INV_X1    g531(.A(new_n653), .ZN(new_n733));
  NOR4_X1   g532(.A1(new_n536), .A2(new_n733), .A3(new_n634), .A4(new_n601), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n494), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n657), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n495), .ZN(G1332gat));
  AOI211_X1 g536(.A(new_n662), .B(new_n735), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1333gat));
  NOR3_X1   g539(.A1(new_n735), .A2(G71gat), .A3(new_n676), .ZN(new_n741));
  INV_X1    g540(.A(new_n735), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n674), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(G71gat), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g544(.A1(new_n735), .A2(new_n273), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(new_n501), .ZN(G1335gat));
  INV_X1    g546(.A(new_n536), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n634), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n699), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n749), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n733), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n658), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n748), .A2(new_n733), .A3(new_n634), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT114), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n691), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n657), .A2(new_n406), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(G1336gat));
  NAND4_X1  g559(.A1(new_n687), .A2(new_n448), .A3(new_n690), .A4(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n752), .A2(new_n753), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n448), .A2(new_n438), .A3(new_n653), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT115), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT52), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n762), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1337gat));
  AOI21_X1  g570(.A(G99gat), .B1(new_n754), .B2(new_n677), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n491), .A2(new_n280), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n758), .B2(new_n773), .ZN(G1338gat));
  AOI21_X1  g573(.A(G106gat), .B1(new_n754), .B2(new_n462), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n462), .A2(G106gat), .ZN(new_n777));
  AND4_X1   g576(.A1(new_n687), .A2(new_n690), .A3(new_n757), .A4(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n779), .A3(KEYINPUT53), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n775), .B2(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1339gat));
  OAI211_X1 g582(.A(new_n636), .B(new_n643), .C1(new_n639), .C2(KEYINPUT10), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n651), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n642), .A2(KEYINPUT54), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n642), .A2(KEYINPUT116), .A3(KEYINPUT54), .A4(new_n784), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n652), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT117), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(new_n796), .A3(new_n652), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n792), .A2(new_n634), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n618), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n630), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n620), .A2(new_n626), .A3(new_n624), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n584), .A2(new_n585), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n628), .B1(new_n530), .B2(new_n802), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n622), .A2(new_n801), .B1(new_n803), .B2(new_n605), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n617), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n653), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n601), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n601), .A3(new_n795), .A4(new_n797), .ZN(new_n809));
  INV_X1    g608(.A(new_n806), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n536), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n602), .A2(new_n733), .A3(new_n635), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n657), .A2(new_n448), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n467), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n634), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G113gat), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n283), .A2(new_n284), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n819), .ZN(G1340gat));
  NOR2_X1   g621(.A1(new_n817), .A2(new_n733), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(new_n297), .ZN(G1341gat));
  NOR2_X1   g623(.A1(new_n817), .A2(new_n536), .ZN(new_n825));
  NOR2_X1   g624(.A1(KEYINPUT118), .A2(G127gat), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT119), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n825), .B(new_n827), .ZN(G1342gat));
  NAND2_X1  g627(.A1(new_n818), .A2(new_n601), .ZN(new_n829));
  NOR2_X1   g628(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n830));
  AND2_X1   g629(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n829), .B2(new_n830), .ZN(G1343gat));
  NOR4_X1   g632(.A1(new_n536), .A2(new_n653), .A3(new_n634), .A4(new_n601), .ZN(new_n834));
  INV_X1    g633(.A(new_n791), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n631), .A2(new_n633), .B1(new_n794), .B2(new_n793), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n835), .A2(new_n836), .B1(new_n806), .B2(new_n653), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n837), .A2(new_n601), .B1(new_n810), .B2(new_n809), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n834), .B1(new_n838), .B2(new_n536), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT57), .B1(new_n839), .B2(new_n273), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n814), .A2(new_n841), .A3(new_n462), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n491), .A2(new_n815), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT120), .Z(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G141gat), .B1(new_n845), .B2(new_n635), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n814), .A2(new_n462), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n843), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n231), .A3(new_n634), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n229), .A3(new_n653), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT121), .ZN(new_n853));
  INV_X1    g652(.A(new_n845), .ZN(new_n854));
  AOI211_X1 g653(.A(KEYINPUT59), .B(new_n229), .C1(new_n854), .C2(new_n653), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n273), .A2(KEYINPUT57), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n809), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n809), .A2(new_n859), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n806), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n837), .A2(new_n601), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n748), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n858), .B1(new_n864), .B2(new_n834), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n857), .A2(new_n865), .A3(new_n653), .A4(new_n844), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n856), .B1(new_n866), .B2(G148gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n853), .B1(new_n855), .B2(new_n867), .ZN(G1345gat));
  AOI21_X1  g667(.A(G155gat), .B1(new_n848), .B2(new_n748), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n536), .A2(new_n223), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n854), .B2(new_n870), .ZN(G1346gat));
  AOI21_X1  g670(.A(G162gat), .B1(new_n848), .B2(new_n601), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n685), .A2(new_n224), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n854), .B2(new_n873), .ZN(G1347gat));
  AOI21_X1  g673(.A(new_n658), .B1(new_n812), .B2(new_n813), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n875), .A2(new_n448), .A3(new_n467), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n616), .A3(new_n634), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n657), .A2(new_n448), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n676), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT123), .Z(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n814), .A3(new_n273), .ZN(new_n881));
  OAI21_X1  g680(.A(G169gat), .B1(new_n881), .B2(new_n635), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n877), .A2(new_n882), .ZN(G1348gat));
  NOR3_X1   g682(.A1(new_n881), .A2(new_n647), .A3(new_n733), .ZN(new_n884));
  AOI21_X1  g683(.A(G176gat), .B1(new_n876), .B2(new_n653), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(KEYINPUT124), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(KEYINPUT124), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(G1349gat));
  NAND3_X1  g687(.A1(new_n876), .A2(new_n748), .A3(new_n330), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT60), .ZN(new_n891));
  OAI21_X1  g690(.A(G183gat), .B1(new_n881), .B2(new_n536), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n890), .A2(KEYINPUT60), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n881), .B2(new_n685), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT61), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n331), .A3(new_n601), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1351gat));
  XNOR2_X1  g698(.A(KEYINPUT126), .B(G197gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n674), .A2(new_n878), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n857), .A2(new_n865), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n902), .B2(new_n635), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n273), .A2(new_n662), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n875), .A2(new_n491), .A3(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n635), .A2(new_n900), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(G1352gat));
  INV_X1    g706(.A(KEYINPUT127), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n857), .A2(new_n865), .A3(new_n653), .A4(new_n901), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(G204gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n733), .A2(G204gat), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n875), .A2(new_n491), .A3(new_n904), .A4(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT62), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n908), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n913), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n909), .A2(G204gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT127), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n917), .ZN(G1353gat));
  INV_X1    g717(.A(new_n905), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n214), .A3(new_n748), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n857), .A2(new_n865), .A3(new_n748), .A4(new_n901), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1354gat));
  NOR3_X1   g723(.A1(new_n902), .A2(new_n215), .A3(new_n685), .ZN(new_n925));
  AOI21_X1  g724(.A(G218gat), .B1(new_n919), .B2(new_n601), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(G1355gat));
endmodule


