//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT28), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n202), .A2(new_n214), .A3(new_n203), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n206), .A2(new_n207), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n207), .A2(KEYINPUT24), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n208), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(new_n203), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT24), .A3(new_n207), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n212), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT25), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n221), .A2(new_n227), .A3(new_n212), .A4(new_n224), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n216), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT71), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232));
  NAND2_X1  g031(.A1(G226gat), .A2(G233gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G197gat), .B(G204gat), .Z(new_n235));
  AOI21_X1  g034(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT70), .Z(new_n240));
  OR2_X1    g039(.A1(new_n229), .A2(new_n233), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n233), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n231), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n232), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n233), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT72), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT72), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n248), .A3(new_n233), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n244), .A2(new_n239), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(G64gat), .B(G92gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(KEYINPUT30), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n255), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n250), .A3(new_n256), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT73), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT30), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n259), .B2(new_n261), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n257), .B(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT74), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n271));
  INV_X1    g070(.A(G155gat), .ZN(new_n272));
  INV_X1    g071(.A(G162gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n271), .B1(new_n274), .B2(new_n267), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(KEYINPUT2), .ZN(new_n277));
  INV_X1    g076(.A(G148gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(G141gat), .ZN(new_n279));
  INV_X1    g078(.A(G141gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(G148gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n277), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n267), .B1(new_n274), .B2(KEYINPUT2), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(KEYINPUT75), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G148gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n280), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT76), .B(new_n284), .C1(new_n288), .C2(new_n279), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n279), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT75), .B(G148gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n280), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT76), .B1(new_n293), .B2(new_n284), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n283), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G113gat), .B(G120gat), .Z(new_n297));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n299), .B(new_n300), .Z(new_n303));
  INV_X1    g102(.A(KEYINPUT77), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(KEYINPUT77), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n302), .B1(new_n307), .B2(new_n296), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n266), .B1(new_n309), .B2(KEYINPUT5), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT4), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n285), .A2(new_n287), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n279), .B1(new_n314), .B2(G141gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n277), .B1(new_n268), .B2(new_n269), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI221_X4 g116(.A(new_n312), .B1(new_n282), .B2(new_n276), .C1(new_n317), .C2(new_n289), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n289), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT80), .B1(new_n319), .B2(new_n283), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n311), .B(new_n301), .C1(new_n318), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT82), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n302), .A2(KEYINPUT4), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n295), .A2(new_n312), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(KEYINPUT80), .A3(new_n283), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT82), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n326), .A2(new_n327), .A3(new_n311), .A4(new_n301), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n322), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT79), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n295), .A2(KEYINPUT3), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n305), .A3(new_n306), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n295), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n334), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n301), .B(new_n304), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT79), .A4(new_n331), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n329), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT5), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n310), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT4), .B1(new_n296), .B2(new_n301), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n303), .B1(new_n324), .B2(new_n325), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(KEYINPUT4), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n339), .A2(KEYINPUT5), .A3(new_n266), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n348));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT6), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n340), .A2(new_n341), .ZN(new_n355));
  INV_X1    g154(.A(new_n310), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(new_n352), .A3(new_n346), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n347), .A2(new_n360), .A3(new_n353), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n265), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n232), .B1(new_n295), .B2(new_n333), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n240), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G228gat), .ZN(new_n365));
  INV_X1    g164(.A(G233gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n295), .A2(new_n232), .A3(new_n239), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n364), .A2(new_n331), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n239), .A2(new_n232), .ZN(new_n370));
  INV_X1    g169(.A(new_n333), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(new_n324), .A3(new_n325), .ZN(new_n373));
  INV_X1    g172(.A(new_n239), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n367), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT83), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n378));
  AOI211_X1 g177(.A(new_n378), .B(new_n367), .C1(new_n373), .C2(new_n375), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n369), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT31), .B(G50gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(G22gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n381), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n369), .C1(new_n377), .C2(new_n379), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n382), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(new_n382), .B2(new_n386), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n362), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G15gat), .B(G43gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n229), .A2(new_n303), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n301), .A2(new_n216), .A3(new_n226), .A4(new_n228), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n398), .B(KEYINPUT64), .Z(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT32), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n394), .B1(new_n401), .B2(KEYINPUT66), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT67), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT33), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT66), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n400), .A2(new_n406), .A3(KEYINPUT32), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n402), .A2(new_n403), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n399), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n395), .B2(new_n396), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT32), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT66), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n407), .A2(new_n405), .A3(new_n412), .A4(new_n393), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT67), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n401), .B1(KEYINPUT33), .B2(new_n393), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT34), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n397), .B2(new_n399), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n395), .A2(KEYINPUT34), .A3(new_n409), .A4(new_n396), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n418), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT36), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n420), .A2(KEYINPUT68), .A3(new_n421), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n415), .B2(new_n417), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n416), .B(new_n427), .C1(new_n408), .C2(new_n414), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT36), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT69), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n429), .A2(new_n431), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT69), .A3(KEYINPUT36), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n390), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n357), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n342), .A2(KEYINPUT86), .A3(new_n352), .A4(new_n346), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n266), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n340), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n309), .A2(new_n266), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(KEYINPUT39), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n266), .B1(new_n329), .B2(new_n339), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n352), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(KEYINPUT40), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n443), .A2(new_n264), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n340), .A2(new_n449), .A3(new_n444), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n353), .ZN(new_n455));
  INV_X1    g254(.A(new_n446), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n448), .A2(new_n449), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n453), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT40), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n447), .A2(KEYINPUT84), .A3(new_n450), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT85), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n458), .A2(KEYINPUT85), .A3(new_n459), .A4(new_n460), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n452), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n361), .B1(new_n443), .B2(new_n354), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n255), .B1(new_n251), .B2(KEYINPUT37), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n247), .A2(new_n249), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n239), .B1(new_n470), .B2(new_n244), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n240), .B1(new_n234), .B2(new_n241), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n251), .A2(KEYINPUT37), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT38), .B1(new_n475), .B2(new_n467), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n474), .A2(new_n476), .A3(new_n259), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n389), .B1(new_n466), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n465), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT87), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n439), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  INV_X1    g283(.A(new_n436), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n484), .B1(new_n485), .B2(new_n389), .ZN(new_n486));
  INV_X1    g285(.A(new_n361), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n264), .B1(new_n358), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n387), .A2(new_n388), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(KEYINPUT88), .A3(new_n436), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n418), .B(new_n422), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n489), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n493), .A2(KEYINPUT35), .A3(new_n466), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n491), .A2(KEYINPUT35), .B1(new_n494), .B2(new_n265), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT89), .B1(new_n483), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT69), .B1(new_n436), .B2(KEYINPUT36), .ZN(new_n497));
  NOR4_X1   g296(.A1(new_n429), .A2(new_n431), .A3(new_n434), .A4(new_n425), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n499), .A2(new_n426), .B1(new_n362), .B2(new_n389), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n465), .A2(new_n478), .A3(new_n481), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n481), .B1(new_n465), .B2(new_n478), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n494), .A2(new_n265), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n496), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G8gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(G1gat), .B2(new_n511), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n515), .B(new_n516), .Z(new_n517));
  NAND2_X1  g316(.A1(KEYINPUT96), .A2(G57gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G64gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(G71gat), .A2(G78gat), .ZN(new_n520));
  OR2_X1    g319(.A1(G71gat), .A2(G78gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G57gat), .A2(G64gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT9), .ZN(new_n526));
  NOR2_X1   g325(.A1(G57gat), .A2(G64gat), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n520), .B(new_n521), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT21), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n517), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(new_n222), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n529), .A2(KEYINPUT21), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G231gat), .A2(G233gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G211gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n536), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  INV_X1    g340(.A(G29gat), .ZN(new_n542));
  INV_X1    g341(.A(G36gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT14), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n544), .B(new_n546), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  XOR2_X1   g346(.A(G43gat), .B(G50gat), .Z(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(KEYINPUT90), .B2(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n547), .A2(new_n548), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT15), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT7), .ZN(new_n557));
  INV_X1    g356(.A(G99gat), .ZN(new_n558));
  INV_X1    g357(.A(G106gat), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT8), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n557), .B(new_n560), .C1(G85gat), .C2(G92gat), .ZN(new_n561));
  XOR2_X1   g360(.A(G99gat), .B(G106gat), .Z(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n555), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n567), .B(new_n568), .C1(new_n566), .C2(new_n553), .ZN(new_n569));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n570), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n578), .A2(KEYINPUT97), .ZN(new_n579));
  OR3_X1    g378(.A1(new_n569), .A2(new_n573), .A3(new_n570), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(KEYINPUT97), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n575), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n572), .A2(new_n578), .A3(new_n574), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n564), .A2(KEYINPUT10), .A3(new_n529), .A4(new_n565), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT100), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(KEYINPUT100), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n529), .B1(new_n563), .B2(KEYINPUT99), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n566), .B(new_n589), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n587), .B(new_n588), .C1(new_n591), .C2(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n593), .B2(new_n590), .ZN(new_n595));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT101), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n598), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n541), .A2(new_n585), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT102), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n555), .A2(new_n517), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT92), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT92), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n555), .A2(new_n608), .A3(new_n517), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n607), .B(new_n609), .C1(new_n517), .C2(new_n553), .ZN(new_n610));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT18), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G113gat), .B(G141gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(G197gat), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT11), .B(G169gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  XOR2_X1   g421(.A(new_n517), .B(new_n553), .Z(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n611), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n617), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n617), .A2(KEYINPUT95), .A3(new_n622), .A4(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n627), .ZN(new_n633));
  INV_X1    g432(.A(new_n622), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n509), .A2(new_n605), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n359), .A2(new_n361), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g440(.A1(new_n637), .A2(new_n265), .ZN(new_n642));
  NAND2_X1  g441(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n512), .A2(new_n510), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT42), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n510), .B2(new_n642), .ZN(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n637), .A2(new_n648), .A3(new_n438), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n637), .A2(new_n424), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n648), .B2(new_n650), .ZN(G1326gat));
  NOR2_X1   g450(.A1(new_n637), .A2(new_n489), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G22gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NAND3_X1  g454(.A1(new_n496), .A2(new_n584), .A3(new_n508), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT44), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n503), .A2(KEYINPUT105), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n659), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n507), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n584), .B(KEYINPUT106), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n630), .A2(new_n631), .B1(new_n634), .B2(new_n633), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n666), .A2(new_n541), .A3(new_n602), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n638), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(G29gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n509), .A2(new_n584), .A3(new_n667), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(G29gat), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n672), .B2(new_n639), .ZN(new_n673));
  OR4_X1    g472(.A1(KEYINPUT104), .A2(new_n671), .A3(G29gat), .A4(new_n639), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n673), .B2(new_n674), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n670), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(KEYINPUT107), .B(new_n670), .C1(new_n676), .C2(new_n677), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1328gat));
  NOR2_X1   g481(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n671), .A2(G36gat), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n264), .ZN(new_n685));
  NAND2_X1  g484(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n668), .A2(new_n264), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n543), .B2(new_n688), .ZN(G1329gat));
  INV_X1    g488(.A(G43gat), .ZN(new_n690));
  INV_X1    g489(.A(new_n438), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n668), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n671), .A2(G43gat), .A3(new_n424), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT110), .B1(new_n692), .B2(new_n695), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n692), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n702), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n698), .A3(new_n697), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1330gat));
  NOR3_X1   g505(.A1(new_n671), .A2(G50gat), .A3(new_n489), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n668), .A2(new_n389), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(G50gat), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1331gat));
  NAND2_X1  g512(.A1(new_n661), .A2(new_n666), .ZN(new_n714));
  INV_X1    g513(.A(new_n541), .ZN(new_n715));
  NOR4_X1   g514(.A1(new_n714), .A2(new_n715), .A3(new_n584), .A4(new_n603), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n638), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n716), .A2(new_n264), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT112), .ZN(new_n721));
  NOR2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1333gat));
  NAND3_X1  g522(.A1(new_n716), .A2(G71gat), .A3(new_n691), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n716), .A2(new_n492), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(G71gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n716), .A2(new_n389), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g528(.A1(new_n636), .A2(new_n541), .A3(new_n585), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n661), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT51), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n661), .A2(new_n733), .A3(new_n730), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n732), .A2(new_n602), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n638), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n715), .A2(new_n602), .A3(new_n666), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n657), .B2(new_n664), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n638), .A2(G85gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(G1336gat));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n732), .A2(new_n602), .A3(new_n264), .A4(new_n734), .ZN(new_n744));
  INV_X1    g543(.A(G92gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n265), .A2(new_n745), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n743), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n744), .A2(new_n745), .B1(new_n740), .B2(new_n747), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n753));
  AND4_X1   g552(.A1(KEYINPUT114), .A2(new_n746), .A3(KEYINPUT52), .A4(new_n748), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT114), .B1(new_n752), .B2(KEYINPUT52), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n751), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n749), .B2(new_n750), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n752), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n762), .B(KEYINPUT116), .C1(new_n751), .C2(new_n753), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n758), .A2(new_n763), .ZN(G1337gat));
  INV_X1    g563(.A(new_n740), .ZN(new_n765));
  OAI21_X1  g564(.A(G99gat), .B1(new_n765), .B2(new_n438), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n735), .A2(new_n558), .A3(new_n492), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(G1338gat));
  OAI21_X1  g567(.A(G106gat), .B1(new_n765), .B2(new_n489), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT53), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n735), .A2(new_n559), .A3(new_n389), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n771), .B(new_n773), .Z(G1339gat));
  INV_X1    g573(.A(new_n663), .ZN(new_n775));
  INV_X1    g574(.A(new_n598), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n592), .A2(new_n593), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(KEYINPUT54), .A3(new_n594), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI221_X1 g579(.A(new_n780), .B1(new_n779), .B2(new_n778), .C1(KEYINPUT54), .C2(new_n594), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n600), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n666), .A2(new_n785), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n610), .A2(new_n612), .B1(new_n623), .B2(new_n626), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n787), .A2(new_n621), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n632), .A2(new_n602), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n775), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n632), .A2(new_n788), .ZN(new_n791));
  INV_X1    g590(.A(new_n785), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n663), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n541), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n604), .A2(new_n636), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n639), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n486), .A2(new_n490), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n264), .ZN(new_n800));
  INV_X1    g599(.A(G113gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n801), .A3(new_n636), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n796), .A2(new_n493), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n639), .A2(new_n264), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G113gat), .B1(new_n805), .B2(new_n666), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n802), .A2(new_n806), .ZN(G1340gat));
  INV_X1    g606(.A(G120gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n800), .A2(new_n808), .A3(new_n602), .ZN(new_n809));
  OAI21_X1  g608(.A(G120gat), .B1(new_n805), .B2(new_n603), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1341gat));
  INV_X1    g610(.A(G127gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n805), .A2(new_n812), .A3(new_n715), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n800), .A2(new_n541), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n812), .ZN(G1342gat));
  NOR4_X1   g614(.A1(new_n799), .A2(G134gat), .A3(new_n585), .A4(new_n264), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT56), .ZN(new_n817));
  OAI21_X1  g616(.A(G134gat), .B1(new_n805), .B2(new_n585), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1343gat));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(new_n389), .C1(new_n794), .C2(new_n795), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n438), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n789), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n781), .A2(KEYINPUT119), .A3(new_n782), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n781), .A2(KEYINPUT119), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT55), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n636), .A2(new_n600), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n584), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n793), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n715), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n795), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n489), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n821), .B(new_n823), .C1(new_n833), .C2(new_n820), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(KEYINPUT121), .A3(new_n636), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n834), .B2(new_n666), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(G141gat), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n797), .A2(new_n389), .A3(new_n438), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n666), .A2(G141gat), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n797), .A2(KEYINPUT120), .A3(new_n389), .A4(new_n438), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n843), .A2(new_n265), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n839), .A2(new_n840), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n280), .B1(new_n835), .B2(new_n636), .ZN(new_n848));
  NOR4_X1   g647(.A1(new_n841), .A2(G141gat), .A3(new_n264), .A4(new_n666), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT58), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n843), .A2(new_n845), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n853), .A2(new_n314), .A3(new_n602), .A4(new_n265), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n314), .B1(new_n835), .B2(new_n602), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n855), .A2(KEYINPUT59), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n791), .A2(new_n584), .A3(new_n792), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n715), .B1(new_n829), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n605), .A2(new_n666), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n820), .A3(new_n389), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT57), .B1(new_n796), .B2(new_n489), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n823), .A2(new_n602), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT59), .B(G148gat), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n854), .A2(new_n856), .A3(new_n865), .ZN(G1345gat));
  NOR3_X1   g665(.A1(new_n834), .A2(new_n272), .A3(new_n715), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n853), .A2(new_n541), .A3(new_n265), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n272), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n834), .B2(new_n775), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n584), .A2(new_n273), .A3(new_n265), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n852), .B2(new_n871), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n638), .A2(new_n265), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n803), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G169gat), .B1(new_n874), .B2(new_n666), .ZN(new_n875));
  INV_X1    g674(.A(new_n796), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n798), .A3(new_n873), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n666), .A2(G169gat), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(G1348gat));
  INV_X1    g678(.A(G176gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n877), .B2(new_n603), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT122), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n874), .A2(new_n880), .A3(new_n603), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(G1349gat));
  INV_X1    g683(.A(new_n877), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n541), .A3(new_n202), .ZN(new_n886));
  OAI21_X1  g685(.A(G183gat), .B1(new_n874), .B2(new_n715), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(G1350gat));
  NOR3_X1   g689(.A1(new_n877), .A2(G190gat), .A3(new_n775), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT124), .ZN(new_n892));
  OAI21_X1  g691(.A(G190gat), .B1(new_n874), .B2(new_n585), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(G1351gat));
  AND2_X1   g696(.A1(new_n873), .A2(new_n438), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT126), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n863), .A2(new_n666), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(KEYINPUT125), .B(G197gat), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n876), .A2(new_n389), .A3(new_n898), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n636), .A2(new_n903), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n901), .A2(new_n903), .B1(new_n904), .B2(new_n905), .ZN(G1352gat));
  INV_X1    g705(.A(new_n863), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n602), .A3(new_n899), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n907), .A2(KEYINPUT127), .A3(new_n602), .A4(new_n899), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(G204gat), .A3(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n904), .A2(G204gat), .A3(new_n603), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT62), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1353gat));
  OR3_X1    g714(.A1(new_n904), .A2(G211gat), .A3(new_n715), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n907), .A2(new_n541), .A3(new_n899), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n917), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT63), .B1(new_n917), .B2(G211gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(G1354gat));
  NOR3_X1   g719(.A1(new_n863), .A2(new_n585), .A3(new_n900), .ZN(new_n921));
  INV_X1    g720(.A(G218gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n663), .A2(new_n922), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n921), .A2(new_n922), .B1(new_n904), .B2(new_n923), .ZN(G1355gat));
endmodule


