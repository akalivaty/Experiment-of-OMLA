//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n215), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n209), .B1(new_n213), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G68), .Z(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n210), .ZN(new_n251));
  AND2_X1   g0051(.A1(G58), .A2(G68), .ZN(new_n252));
  OAI21_X1  g0052(.A(G20), .B1(new_n252), .B2(new_n201), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G159), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n253), .A2(KEYINPUT77), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT77), .B1(new_n253), .B2(new_n255), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT7), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n260), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT76), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT76), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n263), .A2(new_n269), .A3(new_n264), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n270), .A3(new_n211), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n265), .B1(new_n271), .B2(new_n259), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n258), .B(KEYINPUT16), .C1(new_n272), .C2(new_n215), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n253), .A2(new_n255), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT77), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n253), .A2(KEYINPUT77), .A3(new_n255), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT67), .B1(new_n266), .B2(new_n267), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n263), .A2(new_n280), .A3(new_n264), .ZN(new_n281));
  AOI21_X1  g0081(.A(G20), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT78), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n266), .A2(new_n267), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(new_n260), .ZN(new_n285));
  AND4_X1   g0085(.A1(new_n283), .A2(new_n260), .A3(new_n263), .A4(new_n264), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n282), .A2(KEYINPUT7), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n278), .B1(new_n287), .B2(G68), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n251), .B(new_n273), .C1(new_n288), .C2(KEYINPUT16), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT69), .A2(G58), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT8), .ZN(new_n291));
  INV_X1    g0091(.A(G1), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n251), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(G1), .B2(new_n211), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(new_n297), .B2(new_n291), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G41), .ZN(new_n300));
  OAI211_X1 g0100(.A(G1), .B(G13), .C1(new_n262), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G226), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G1698), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n303), .B1(G223), .B2(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G87), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G45), .ZN(new_n307));
  AOI21_X1  g0107(.A(G1), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n301), .A2(G274), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n292), .B1(G41), .B2(G45), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n311), .B2(new_n237), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(G200), .B2(new_n313), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n289), .A2(new_n299), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT17), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT18), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n273), .A2(new_n251), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT16), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT67), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n280), .B1(new_n263), .B2(new_n264), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n211), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n259), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n284), .A2(new_n260), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n265), .A2(new_n283), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n215), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n322), .B1(new_n331), .B2(new_n278), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n298), .B1(new_n321), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  INV_X1    g0134(.A(new_n306), .ZN(new_n335));
  INV_X1    g0135(.A(new_n312), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n306), .A2(new_n312), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n320), .B1(new_n333), .B2(new_n340), .ZN(new_n341));
  AOI211_X1 g0141(.A(new_n320), .B(new_n340), .C1(new_n289), .C2(new_n299), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(KEYINPUT79), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n289), .A2(new_n299), .ZN(new_n344));
  INV_X1    g0144(.A(new_n340), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT79), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n320), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n319), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n279), .A2(new_n281), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G77), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n279), .A2(new_n281), .A3(G223), .A4(G1698), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G1698), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n354), .A2(G222), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n279), .A2(new_n281), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT68), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT68), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n279), .A2(new_n281), .A3(new_n358), .A4(new_n355), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n301), .B1(new_n353), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n309), .B1(new_n311), .B2(new_n302), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n334), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n362), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n351), .A2(new_n352), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n359), .B2(new_n357), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n338), .B(new_n364), .C1(new_n366), .C2(new_n301), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n291), .A2(new_n211), .A3(G33), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n254), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n296), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n293), .A2(G50), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n251), .B1(new_n292), .B2(G20), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n372), .B1(new_n373), .B2(G50), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n363), .A2(new_n367), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n294), .A2(new_n224), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n297), .B2(new_n224), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G20), .A2(G77), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n211), .A2(G33), .ZN(new_n381));
  INV_X1    g0181(.A(new_n254), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT8), .B(G58), .ZN(new_n383));
  OAI221_X1 g0183(.A(new_n379), .B1(new_n380), .B2(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n378), .B1(new_n251), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n309), .B1(new_n311), .B2(new_n225), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n323), .A2(new_n324), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n219), .A2(G1698), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G232), .B2(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT70), .B(G107), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n301), .B1(new_n350), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n386), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G200), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n385), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT71), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT71), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n385), .B(new_n397), .C1(new_n393), .C2(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(G190), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n385), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n393), .A2(new_n338), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n401), .B(new_n402), .C1(G169), .C2(new_n393), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(G200), .B1(new_n361), .B2(new_n362), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT10), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT9), .ZN(new_n408));
  INV_X1    g0208(.A(new_n374), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(new_n370), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n371), .A2(KEYINPUT9), .A3(new_n374), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n405), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(G190), .B(new_n364), .C1(new_n366), .C2(new_n301), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n405), .A2(new_n413), .A3(new_n410), .A4(new_n411), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(KEYINPUT10), .A3(new_n406), .ZN(new_n416));
  AOI211_X1 g0216(.A(new_n376), .B(new_n404), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n382), .A2(new_n202), .B1(new_n211), .B2(G68), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n381), .A2(new_n224), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n251), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT11), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT73), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n422), .ZN(new_n424));
  OR3_X1    g0224(.A1(new_n293), .A2(KEYINPUT12), .A3(G68), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT12), .B1(new_n293), .B2(G68), .ZN(new_n426));
  AOI22_X1  g0226(.A1(G68), .A2(new_n373), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n302), .A2(new_n354), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n237), .A2(G1698), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n279), .A2(new_n281), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G97), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n262), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n309), .B1(new_n311), .B2(new_n219), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT13), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n301), .B1(new_n432), .B2(new_n435), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT13), .B1(new_n443), .B2(new_n439), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n429), .B1(new_n445), .B2(G169), .ZN(new_n446));
  AOI211_X1 g0246(.A(KEYINPUT14), .B(new_n334), .C1(new_n442), .C2(new_n444), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT74), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n445), .B2(new_n338), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n442), .A2(new_n444), .A3(KEYINPUT74), .A4(G179), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n448), .A2(KEYINPUT75), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT75), .B1(new_n448), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n428), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n445), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n428), .B1(new_n456), .B2(G190), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n445), .A2(G200), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AND4_X1   g0260(.A1(new_n349), .A2(new_n417), .A3(new_n455), .A4(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT81), .B1(new_n262), .B2(G1), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n462), .A2(new_n293), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT81), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n292), .A3(G33), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n463), .A2(KEYINPUT82), .A3(new_n296), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT82), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(new_n465), .A3(new_n293), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(new_n251), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(G107), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n226), .A2(G20), .ZN(new_n471));
  INV_X1    g0271(.A(G13), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n471), .A2(G1), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT25), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT89), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n211), .A2(G87), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT22), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT87), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(new_n279), .A3(new_n281), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n211), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  OAI22_X1  g0288(.A1(KEYINPUT23), .A2(new_n471), .B1(new_n381), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n391), .A2(G20), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(KEYINPUT23), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n487), .A2(new_n491), .A3(new_n493), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n477), .B1(new_n497), .B2(new_n251), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n487), .A2(new_n491), .A3(new_n493), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n493), .B1(new_n487), .B2(new_n491), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n477), .B(new_n251), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n476), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G250), .A2(G1698), .ZN(new_n504));
  INV_X1    g0304(.A(G257), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(G1698), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n263), .A2(new_n264), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G294), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT90), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n437), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n307), .A2(G1), .ZN(new_n513));
  OR2_X1    g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n437), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n301), .A2(G274), .ZN(new_n518));
  INV_X1    g0318(.A(new_n515), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n513), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n517), .A2(G264), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n506), .A2(new_n507), .B1(G33), .B2(G294), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT90), .B1(new_n524), .B2(new_n301), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n512), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G169), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n518), .A2(new_n522), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n521), .A2(G264), .A3(new_n301), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(new_n524), .C2(new_n301), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n338), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n503), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G303), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n279), .B2(new_n281), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n227), .A2(G1698), .ZN(new_n535));
  OAI221_X1 g0335(.A(new_n535), .B1(G257), .B2(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n437), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n517), .A2(G270), .B1(new_n518), .B2(new_n522), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n463), .A2(G116), .A3(new_n296), .A4(new_n465), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n294), .A2(new_n488), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n250), .A2(new_n210), .B1(G20), .B2(new_n488), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G283), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n211), .C1(G33), .C2(new_n433), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n544), .A2(KEYINPUT20), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT20), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n542), .B(new_n543), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n538), .A2(new_n539), .A3(G190), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n541), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n540), .A2(G169), .A3(new_n549), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT21), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n549), .A2(G179), .A3(new_n538), .A4(new_n539), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n334), .B1(new_n538), .B2(new_n539), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(KEYINPUT21), .A3(new_n549), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n552), .A2(new_n555), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n219), .A2(new_n354), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n225), .A2(G1698), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(new_n266), .C2(new_n267), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT85), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G116), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n437), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n513), .A2(new_n221), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n518), .A2(new_n513), .B1(new_n301), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n334), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT86), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(KEYINPUT19), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(KEYINPUT86), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n434), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(G87), .A2(G97), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(new_n211), .B1(new_n577), .B2(new_n391), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n574), .A2(KEYINPUT86), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n572), .A2(KEYINPUT19), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n579), .B(new_n580), .C1(new_n381), .C2(new_n433), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n211), .B(G68), .C1(new_n266), .C2(new_n267), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n251), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n380), .A2(new_n294), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n466), .A2(new_n469), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n380), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n567), .A2(new_n338), .A3(new_n569), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n571), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n466), .A2(G87), .A3(new_n469), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n584), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n562), .A2(new_n564), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT85), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n301), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n569), .ZN(new_n596));
  OAI21_X1  g0396(.A(G200), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n567), .A2(G190), .A3(new_n569), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n591), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n589), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n559), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n512), .A2(new_n523), .A3(new_n525), .A4(new_n314), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n530), .A2(new_n394), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n605), .B(new_n476), .C1(new_n498), .C2(new_n502), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n532), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n294), .A2(G97), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n586), .B2(G97), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT80), .ZN(new_n611));
  INV_X1    g0411(.A(new_n391), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n287), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT6), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n614), .A2(new_n433), .A3(G107), .ZN(new_n615));
  XNOR2_X1  g0415(.A(G97), .B(G107), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n617), .A2(new_n211), .B1(new_n224), .B2(new_n382), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n611), .B1(new_n620), .B2(new_n251), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n287), .B2(new_n612), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n622), .A2(KEYINPUT80), .A3(new_n296), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n610), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT84), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n301), .A2(G274), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(new_n521), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT83), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n517), .A2(new_n628), .A3(G257), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n521), .A2(new_n301), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT83), .B1(new_n630), .B2(new_n505), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n627), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n279), .A2(new_n281), .A3(G250), .A4(G1698), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n354), .A2(G244), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT4), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n279), .A2(new_n281), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n635), .B1(new_n284), .B2(new_n634), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n633), .A2(new_n637), .A3(new_n545), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n437), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n632), .A2(new_n640), .A3(G179), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n334), .B1(new_n632), .B2(new_n640), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n624), .A2(new_n625), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT80), .B1(new_n622), .B2(new_n296), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n391), .B1(new_n326), .B2(new_n330), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n611), .B(new_n251), .C1(new_n646), .C2(new_n618), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n609), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n641), .A2(new_n642), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT84), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n632), .A2(new_n640), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G200), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n632), .A2(new_n640), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G190), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n648), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n644), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n607), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n461), .A2(new_n657), .ZN(G372));
  XNOR2_X1  g0458(.A(new_n317), .B(KEYINPUT17), .ZN(new_n659));
  INV_X1    g0459(.A(new_n428), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT75), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n450), .A2(new_n451), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n441), .B1(new_n438), .B2(new_n440), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n443), .A2(KEYINPUT13), .A3(new_n439), .ZN(new_n664));
  OAI21_X1  g0464(.A(G169), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT14), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n445), .A2(new_n429), .A3(G169), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n661), .B1(new_n662), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n448), .A2(KEYINPUT75), .A3(new_n452), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n660), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n403), .B1(new_n457), .B2(new_n458), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n659), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT18), .B1(new_n344), .B2(new_n345), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n342), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n414), .A2(new_n416), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n376), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n461), .ZN(new_n680));
  INV_X1    g0480(.A(new_n589), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n503), .B2(new_n531), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT91), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n591), .A2(new_n597), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n394), .B1(new_n567), .B2(new_n569), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n584), .A2(new_n585), .A3(new_n590), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT91), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(new_n688), .A3(new_n598), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n606), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n644), .A2(new_n650), .A3(new_n655), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n681), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n624), .A2(new_n689), .A3(new_n643), .A4(new_n589), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT26), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n600), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n625), .B1(new_n624), .B2(new_n643), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT84), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n696), .B1(new_n700), .B2(new_n695), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n679), .B1(new_n680), .B2(new_n703), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT92), .Z(G369));
  NOR3_X1   g0505(.A1(new_n472), .A2(G1), .A3(G20), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT93), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT27), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(G213), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G343), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n550), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n559), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT94), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n682), .A2(new_n714), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n716), .B1(new_n715), .B2(new_n717), .ZN(new_n719));
  INV_X1    g0519(.A(G330), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n251), .B1(new_n499), .B2(new_n500), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT89), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n475), .B1(new_n724), .B2(new_n501), .ZN(new_n725));
  INV_X1    g0525(.A(new_n531), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n475), .B(new_n604), .C1(new_n724), .C2(new_n501), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n713), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n503), .A2(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n729), .A2(new_n731), .B1(new_n727), .B2(new_n730), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n722), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n682), .A2(new_n713), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n532), .A2(new_n735), .A3(new_n606), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n727), .A2(new_n713), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(new_n738), .ZN(G399));
  INV_X1    g0539(.A(new_n207), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G41), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G1), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n391), .A2(new_n488), .A3(new_n577), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n744), .B1(new_n217), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n694), .A2(new_n695), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n700), .B2(new_n695), .ZN(new_n748));
  INV_X1    g0548(.A(new_n598), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n591), .A2(new_n597), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(new_n750), .B2(KEYINPUT91), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n725), .A2(new_n605), .B1(new_n751), .B2(new_n685), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n558), .A2(new_n556), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT21), .B1(new_n557), .B2(new_n549), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n725), .B2(new_n726), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n589), .B1(new_n757), .B2(new_n656), .ZN(new_n758));
  OAI211_X1 g0558(.A(KEYINPUT29), .B(new_n713), .C1(new_n748), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n730), .B1(new_n693), .B2(new_n701), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n761));
  OAI21_X1  g0561(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n692), .A2(new_n729), .A3(new_n601), .A4(new_n713), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n529), .B1(new_n524), .B2(new_n301), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT95), .B1(new_n570), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n540), .A2(new_n338), .ZN(new_n766));
  INV_X1    g0566(.A(new_n764), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT95), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n767), .A2(new_n567), .A3(new_n768), .A4(new_n569), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n765), .A2(new_n653), .A3(new_n766), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT30), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n651), .A2(new_n338), .A3(new_n540), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n773), .A2(KEYINPUT30), .A3(new_n769), .A4(new_n765), .ZN(new_n774));
  AOI21_X1  g0574(.A(G179), .B1(new_n767), .B2(new_n528), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n775), .A2(new_n651), .A3(new_n540), .A4(new_n570), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n772), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n730), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT31), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(KEYINPUT31), .A3(new_n730), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n763), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G330), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n762), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n746), .B1(new_n785), .B2(G1), .ZN(G364));
  NOR2_X1   g0586(.A1(new_n718), .A2(new_n719), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G330), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n472), .A2(G20), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n292), .B1(new_n790), .B2(G45), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n741), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n721), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(G1), .B(G13), .C1(new_n211), .C2(G169), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT98), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT98), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n211), .A2(new_n394), .A3(G179), .A4(G190), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT101), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n226), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(G20), .A2(G179), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT100), .Z(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G190), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G200), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(G190), .A3(G200), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n804), .B1(new_n809), .B2(new_n214), .C1(new_n202), .C2(new_n810), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n806), .A2(new_n314), .A3(G200), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT102), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n812), .A2(KEYINPUT102), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n215), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G179), .A2(G200), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n211), .B1(new_n818), .B2(G190), .ZN(new_n819));
  NOR4_X1   g0619(.A1(new_n211), .A2(new_n314), .A3(new_n394), .A4(G179), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n387), .B1(new_n433), .B2(new_n819), .C1(new_n821), .C2(new_n220), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n818), .A2(G20), .A3(new_n314), .ZN(new_n823));
  INV_X1    g0623(.A(G159), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT32), .ZN(new_n826));
  NOR2_X1   g0626(.A1(G190), .A2(G200), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n806), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n826), .B1(new_n224), .B2(new_n828), .ZN(new_n829));
  OR4_X1    g0629(.A1(new_n811), .A2(new_n817), .A3(new_n822), .A4(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  INV_X1    g0631(.A(G326), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n802), .A2(new_n831), .B1(new_n832), .B2(new_n810), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G322), .B2(new_n808), .ZN(new_n834));
  INV_X1    g0634(.A(G329), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n350), .B1(new_n835), .B2(new_n823), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n821), .A2(new_n533), .B1(new_n837), .B2(new_n819), .ZN(new_n838));
  INV_X1    g0638(.A(new_n828), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n836), .B(new_n838), .C1(G311), .C2(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(KEYINPUT33), .B(G317), .Z(new_n841));
  OAI211_X1 g0641(.A(new_n834), .B(new_n840), .C1(new_n816), .C2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n799), .B1(new_n830), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(G13), .A2(G33), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(G20), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n798), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT99), .Z(new_n848));
  NAND2_X1  g0648(.A1(new_n268), .A2(new_n270), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n740), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(G45), .B2(new_n217), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n851), .A2(KEYINPUT97), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(KEYINPUT97), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(new_n307), .C2(new_n248), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n350), .A2(new_n740), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n855), .A2(G355), .B1(new_n488), .B2(new_n740), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n848), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NOR4_X1   g0657(.A1(new_n843), .A2(new_n741), .A3(new_n857), .A4(new_n792), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n715), .A2(new_n717), .A3(new_n846), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n789), .A2(new_n794), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G396));
  NOR2_X1   g0661(.A1(new_n403), .A2(new_n713), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT104), .Z(new_n863));
  OAI211_X1 g0663(.A(new_n400), .B(new_n403), .C1(new_n385), .C2(new_n713), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n760), .B(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n793), .B1(new_n866), .B2(new_n783), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n783), .B2(new_n866), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n799), .A2(new_n845), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT103), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n793), .B1(new_n870), .B2(G77), .ZN(new_n871));
  INV_X1    g0671(.A(G137), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n810), .A2(new_n872), .B1(new_n828), .B2(new_n824), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G143), .B2(new_n808), .ZN(new_n874));
  INV_X1    g0674(.A(G150), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n816), .B2(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT34), .Z(new_n877));
  NOR2_X1   g0677(.A1(new_n802), .A2(new_n215), .ZN(new_n878));
  INV_X1    g0678(.A(G132), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n849), .B1(new_n879), .B2(new_n823), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n821), .A2(new_n202), .B1(new_n214), .B2(new_n819), .ZN(new_n881));
  OR3_X1    g0681(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n802), .A2(new_n220), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n884), .B1(new_n809), .B2(new_n837), .C1(new_n533), .C2(new_n810), .ZN(new_n885));
  INV_X1    g0685(.A(G311), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n350), .B1(new_n886), .B2(new_n823), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n821), .A2(new_n226), .B1(new_n433), .B2(new_n819), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n887), .B(new_n888), .C1(G116), .C2(new_n839), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n816), .B2(new_n831), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n877), .A2(new_n882), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n871), .B1(new_n891), .B2(new_n798), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n845), .B2(new_n865), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n868), .A2(new_n893), .ZN(G384));
  INV_X1    g0694(.A(new_n617), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n897));
  NOR4_X1   g0697(.A1(new_n896), .A2(new_n897), .A3(new_n488), .A4(new_n213), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT36), .Z(new_n899));
  OAI21_X1  g0699(.A(G77), .B1(new_n214), .B2(new_n215), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n217), .A2(new_n900), .B1(G50), .B2(new_n215), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(G1), .A3(new_n472), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT105), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n344), .A2(KEYINPUT18), .A3(new_n345), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n674), .B1(new_n347), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n348), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n659), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n271), .A2(new_n259), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n215), .B1(new_n909), .B2(new_n327), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n322), .B1(new_n910), .B2(new_n278), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n298), .B1(new_n321), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n912), .A2(new_n711), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n289), .A2(new_n299), .A3(new_n316), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n911), .A2(new_n251), .A3(new_n273), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n340), .B1(new_n917), .B2(new_n299), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT106), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT106), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(new_n317), .C1(new_n912), .C2(new_n340), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n921), .A3(new_n913), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n344), .A2(new_n712), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n346), .A2(new_n924), .A3(new_n317), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(KEYINPUT37), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n915), .A2(new_n928), .A3(KEYINPUT38), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT107), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n319), .A2(new_n675), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n925), .A2(KEYINPUT37), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n931), .A2(new_n924), .B1(new_n932), .B2(new_n926), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT38), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT107), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n915), .A2(new_n928), .A3(new_n936), .A4(KEYINPUT38), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n863), .A2(new_n864), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n428), .A2(new_n730), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n455), .A2(new_n460), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n669), .A2(new_n670), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n428), .B(new_n730), .C1(new_n942), .C2(new_n459), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n939), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n778), .A2(KEYINPUT108), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT108), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n777), .A2(new_n946), .A3(new_n730), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n779), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n781), .A3(new_n763), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n944), .A2(KEYINPUT40), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n938), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT40), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n343), .A2(new_n348), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n913), .B1(new_n953), .B2(new_n659), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n926), .B1(KEYINPUT37), .B2(new_n922), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n954), .A2(new_n955), .A3(new_n934), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT38), .B1(new_n915), .B2(new_n928), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n944), .A2(new_n949), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n951), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n461), .A2(new_n949), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n963), .A2(new_n964), .A3(new_n720), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT109), .Z(new_n966));
  NOR2_X1   g0766(.A1(new_n455), .A2(new_n730), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT39), .B1(new_n933), .B2(new_n934), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n930), .A2(new_n937), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n934), .B1(new_n954), .B2(new_n955), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n929), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT39), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n968), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n681), .B1(new_n751), .B2(new_n685), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n648), .A2(new_n649), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT26), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n600), .B1(new_n644), .B2(new_n650), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n977), .B1(KEYINPUT26), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n713), .B(new_n865), .C1(new_n979), .C2(new_n758), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n730), .A2(new_n403), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n941), .A2(new_n943), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n984), .A2(new_n958), .B1(new_n676), .B2(new_n712), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n974), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n759), .B(new_n461), .C1(new_n760), .C2(new_n761), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n679), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n986), .B(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n966), .A2(new_n990), .B1(new_n292), .B2(new_n790), .ZN(new_n991));
  INV_X1    g0791(.A(new_n966), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n989), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n904), .B1(new_n991), .B2(new_n993), .ZN(G367));
  OAI21_X1  g0794(.A(new_n847), .B1(new_n207), .B2(new_n380), .ZN(new_n995));
  INV_X1    g0795(.A(new_n850), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n234), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n793), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n821), .B2(new_n488), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n820), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n831), .C2(new_n828), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n800), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n1003), .A2(new_n433), .B1(new_n391), .B2(new_n819), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n823), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n849), .B(new_n1004), .C1(G317), .C2(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n533), .B2(new_n809), .C1(new_n886), .C2(new_n810), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n816), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1002), .B(new_n1007), .C1(G294), .C2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT112), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n810), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(G143), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n819), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(G68), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1012), .B(new_n1014), .C1(new_n809), .C2(new_n875), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT113), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1008), .A2(G159), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n821), .A2(new_n214), .B1(new_n1003), .B2(new_n224), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n387), .B1(new_n872), .B2(new_n823), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(G50), .C2(new_n839), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1010), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT47), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n799), .B1(new_n1025), .B2(KEYINPUT47), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n998), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n846), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n975), .B1(new_n591), .B2(new_n713), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n681), .A2(new_n687), .A3(new_n730), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1028), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n736), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n732), .B2(new_n734), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(new_n721), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n784), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT45), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n624), .A2(new_n730), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n644), .A2(new_n650), .A3(new_n1039), .A4(new_n655), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT110), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n976), .B2(new_n730), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT110), .A4(new_n713), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n736), .A2(new_n737), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1038), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n738), .A2(new_n1044), .A3(KEYINPUT45), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT44), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n738), .B2(new_n1044), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1051), .A2(new_n1046), .A3(KEYINPUT44), .A4(new_n1040), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1047), .A2(new_n1048), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n733), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n722), .A2(new_n732), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(KEYINPUT111), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT111), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1053), .B2(new_n733), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1037), .A2(new_n1054), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n785), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n741), .B(KEYINPUT41), .Z(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n792), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1044), .A2(new_n1034), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT42), .Z(new_n1068));
  NOR2_X1   g0868(.A1(new_n1045), .A2(new_n532), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n644), .A2(new_n650), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n713), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1032), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT43), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1032), .A2(KEYINPUT43), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1072), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1068), .A2(new_n1074), .A3(new_n1073), .A4(new_n1071), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n733), .A2(new_n1045), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1077), .A2(new_n1080), .A3(new_n1078), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1033), .B1(new_n1066), .B2(new_n1084), .ZN(G387));
  INV_X1    g0885(.A(new_n1036), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n732), .A2(new_n846), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n855), .A2(new_n744), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(G107), .B2(new_n207), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n240), .A2(G45), .ZN(new_n1090));
  AOI211_X1 g0890(.A(G45), .B(new_n744), .C1(G68), .C2(G77), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n383), .A2(G50), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT50), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n996), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1089), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n793), .B1(new_n1095), .B2(new_n848), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n802), .A2(new_n433), .B1(new_n824), .B2(new_n810), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G50), .B2(new_n808), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1008), .A2(new_n291), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n849), .B1(new_n875), .B2(new_n823), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n820), .A2(G77), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n380), .B2(new_n819), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G68), .C2(new_n839), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1098), .A2(new_n1099), .A3(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n821), .A2(new_n837), .B1(new_n831), .B2(new_n819), .ZN(new_n1105));
  INV_X1    g0905(.A(G322), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n810), .A2(new_n1106), .B1(new_n828), .B2(new_n533), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G317), .B2(new_n808), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n816), .B2(new_n886), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT48), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n1110), .B2(new_n1109), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT49), .Z(new_n1113));
  INV_X1    g0913(.A(new_n849), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n832), .B2(new_n823), .C1(new_n488), .C2(new_n1003), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1104), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1096), .B1(new_n1116), .B2(new_n798), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1086), .A2(new_n792), .B1(new_n1087), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n785), .A2(new_n1086), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n741), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n785), .A2(new_n1086), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(G393));
  OAI21_X1  g0922(.A(new_n847), .B1(new_n433), .B2(new_n207), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n996), .A2(new_n244), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n793), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G311), .A2(new_n808), .B1(new_n1011), .B2(G317), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT52), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1008), .A2(G303), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n839), .A2(G294), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n821), .A2(new_n831), .B1(new_n488), .B2(new_n819), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n387), .B(new_n1130), .C1(G322), .C2(new_n1005), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1128), .A2(new_n804), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1008), .A2(G50), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n828), .A2(new_n383), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n821), .A2(new_n215), .B1(new_n224), .B2(new_n819), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1114), .B(new_n1135), .C1(G143), .C2(new_n1005), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1133), .A2(new_n884), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G159), .A2(new_n808), .B1(new_n1011), .B2(G150), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT51), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1127), .A2(new_n1132), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1125), .B1(new_n1140), .B2(new_n798), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1044), .B2(new_n1029), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1054), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n1144), .B2(new_n791), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n742), .B1(new_n1119), .B2(new_n1144), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n1062), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(G390));
  OAI211_X1 g0948(.A(new_n713), .B(new_n865), .C1(new_n748), .C2(new_n758), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n981), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n967), .B1(new_n1150), .B2(new_n983), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n938), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n970), .A2(new_n973), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n980), .A2(new_n981), .B1(new_n941), .B2(new_n943), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(new_n967), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1152), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n781), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n657), .B2(new_n713), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n720), .B1(new_n1158), .B2(new_n948), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n944), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1156), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n970), .B(new_n973), .C1(new_n967), .C2(new_n1154), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n983), .A2(new_n782), .A3(G330), .A4(new_n865), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1152), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n782), .A2(G330), .A3(new_n865), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n983), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1160), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n982), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1167), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1150), .B1(new_n1172), .B2(new_n983), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n983), .B1(new_n1159), .B2(new_n865), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n461), .A2(new_n949), .A3(G330), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT114), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n987), .A2(new_n679), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n987), .A2(new_n679), .A3(new_n1178), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT114), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1177), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n742), .B1(new_n1166), .B2(new_n1183), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1163), .A2(new_n1152), .A3(new_n1164), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1160), .B1(new_n1163), .B2(new_n1152), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n1180), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1175), .A2(new_n1173), .B1(new_n1170), .B2(new_n982), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1184), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1162), .A2(new_n792), .A3(new_n1165), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n793), .B1(new_n870), .B2(new_n291), .ZN(new_n1194));
  OR3_X1    g0994(.A1(new_n821), .A2(KEYINPUT53), .A3(new_n875), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT53), .B1(new_n821), .B2(new_n875), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT54), .B(G143), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1196), .C1(new_n828), .C2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1008), .B2(G137), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n1003), .A2(new_n202), .B1(new_n824), .B2(new_n819), .ZN(new_n1200));
  INV_X1    g1000(.A(G125), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n387), .B1(new_n1201), .B2(new_n823), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G128), .C2(new_n1011), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1199), .B(new_n1203), .C1(new_n879), .C2(new_n809), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n878), .B1(G116), .B2(new_n808), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n831), .B2(new_n810), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n350), .B1(new_n837), .B2(new_n823), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n821), .A2(new_n220), .B1(new_n224), .B2(new_n819), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(G97), .C2(new_n839), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n816), .B2(new_n391), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1204), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1194), .B1(new_n1211), .B2(new_n798), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT115), .Z(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1153), .B2(new_n845), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1193), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1192), .A2(new_n1216), .ZN(G378));
  INV_X1    g1017(.A(new_n376), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n678), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n712), .A2(new_n375), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT55), .Z(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1219), .B(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1224));
  XNOR2_X1  g1024(.A(new_n1223), .B(new_n1224), .ZN(new_n1225));
  AND4_X1   g1025(.A1(G330), .A2(new_n951), .A3(new_n960), .A4(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n944), .B(new_n949), .C1(new_n956), .C2(new_n957), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n720), .B1(new_n1227), .B2(new_n952), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1225), .B1(new_n1228), .B2(new_n951), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n986), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n951), .A2(new_n960), .A3(G330), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1225), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n974), .A2(new_n985), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1228), .A2(new_n951), .A3(new_n1225), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1230), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1225), .A2(new_n844), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n793), .B1(new_n870), .B2(G50), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n828), .A2(new_n380), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n800), .A2(G58), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1005), .A2(G283), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1101), .A2(new_n1014), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1114), .A2(new_n300), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1240), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G107), .A2(new_n808), .B1(new_n1011), .B2(G116), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n816), .C2(new_n433), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT58), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G50), .B1(new_n262), .B2(new_n300), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1247), .A2(new_n1248), .B1(new_n1244), .B2(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n839), .A2(G137), .B1(G150), .B2(new_n1013), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1201), .B2(new_n810), .ZN(new_n1252));
  INV_X1    g1052(.A(G128), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n809), .A2(new_n1253), .B1(new_n821), .B2(new_n1197), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT116), .Z(new_n1255));
  AOI211_X1 g1055(.A(new_n1252), .B(new_n1255), .C1(G132), .C2(new_n1008), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT59), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n800), .A2(G159), .ZN(new_n1259));
  AOI211_X1 g1059(.A(G33), .B(G41), .C1(new_n1005), .C2(G124), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1257), .A2(KEYINPUT59), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1250), .B1(new_n1248), .B2(new_n1247), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1239), .B1(new_n1263), .B2(new_n798), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1237), .A2(new_n792), .B1(new_n1238), .B2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1180), .B(new_n1182), .C1(new_n1166), .C2(new_n1189), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT57), .B1(new_n1266), .B2(new_n1237), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1188), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1230), .A2(new_n1236), .A3(KEYINPUT57), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n741), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1265), .B1(new_n1267), .B2(new_n1270), .ZN(G375));
  NAND2_X1  g1071(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1183), .A2(new_n1065), .A3(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT118), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1168), .A2(new_n844), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n793), .B1(new_n870), .B2(G68), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n809), .A2(new_n831), .B1(new_n837), .B2(new_n810), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(G77), .B2(new_n801), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n350), .B1(new_n533), .B2(new_n823), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n821), .A2(new_n433), .B1(new_n380), .B2(new_n819), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n1279), .B(new_n1280), .C1(new_n612), .C2(new_n839), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1278), .B(new_n1281), .C1(new_n488), .C2(new_n816), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n849), .B1(new_n1253), .B2(new_n823), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n1241), .B1(new_n202), .B2(new_n819), .C1(new_n821), .C2(new_n824), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(G150), .C2(new_n839), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G137), .A2(new_n808), .B1(new_n1011), .B2(G132), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1285), .B(new_n1286), .C1(new_n816), .C2(new_n1197), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1276), .B1(new_n1288), .B2(new_n798), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1275), .A2(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n791), .B(KEYINPUT119), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1189), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1274), .A2(new_n1293), .ZN(G381));
  NOR3_X1   g1094(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(KEYINPUT120), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1033), .B(new_n1147), .C1(new_n1066), .C2(new_n1084), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(G381), .A2(new_n1296), .A3(G378), .A4(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1298), .B(new_n1265), .C1(new_n1267), .C2(new_n1270), .ZN(G407));
  AOI21_X1  g1099(.A(new_n1215), .B1(new_n1184), .B2(new_n1191), .ZN(new_n1300));
  INV_X1    g1100(.A(G213), .ZN(new_n1301));
  OR3_X1    g1101(.A1(new_n1301), .A2(KEYINPUT121), .A3(G343), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT121), .B1(new_n1301), .B2(G343), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1300), .A2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G407), .B(G213), .C1(G375), .C2(new_n1306), .ZN(G409));
  NAND3_X1  g1107(.A1(new_n1230), .A2(new_n1236), .A3(new_n1065), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1268), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1291), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1230), .A2(new_n1236), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1264), .A2(new_n1238), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1300), .B1(new_n1309), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT122), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G378), .B(new_n1265), .C1(new_n1267), .C2(new_n1270), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT122), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1300), .B(new_n1317), .C1(new_n1309), .C2(new_n1313), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1315), .A2(new_n1316), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1304), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1305), .A2(G2897), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1188), .A2(new_n1189), .A3(KEYINPUT60), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1322), .A2(new_n741), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT60), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1272), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(G384), .B1(new_n1326), .B2(new_n1293), .ZN(new_n1327));
  INV_X1    g1127(.A(G384), .ZN(new_n1328));
  AOI211_X1 g1128(.A(new_n1328), .B(new_n1292), .C1(new_n1323), .C2(new_n1325), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1305), .A2(KEYINPUT124), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1321), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1324), .A2(new_n1272), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1322), .A2(new_n741), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1293), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1328), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1326), .A2(G384), .A3(new_n1293), .ZN(new_n1337));
  AND4_X1   g1137(.A1(new_n1336), .A2(new_n1337), .A3(new_n1321), .A4(new_n1331), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1332), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1319), .A2(new_n1341), .A3(new_n1304), .A4(new_n1330), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1319), .A2(new_n1304), .A3(new_n1330), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(KEYINPUT62), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1340), .A2(new_n1342), .A3(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT126), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(G393), .B(new_n860), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1297), .A2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1064), .B1(new_n1062), .B2(new_n785), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1083), .B(new_n1082), .C1(new_n1349), .C2(new_n792), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1147), .B1(new_n1350), .B2(new_n1033), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1346), .B1(new_n1348), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G387), .A2(G390), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1353), .A2(KEYINPUT126), .A3(new_n1297), .A4(new_n1347), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1352), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT127), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G387), .A2(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1347), .B1(new_n1357), .B2(G390), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(G387), .A2(new_n1356), .A3(new_n1147), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1355), .A2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1345), .A2(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(KEYINPUT125), .B1(new_n1332), .B2(new_n1338), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1336), .A2(new_n1337), .A3(new_n1331), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1365), .A2(G2897), .A3(new_n1305), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT125), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1330), .A2(new_n1321), .A3(new_n1331), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1366), .A2(new_n1367), .A3(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1364), .A2(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1320), .A2(KEYINPUT123), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT123), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1319), .A2(new_n1372), .A3(new_n1304), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1370), .A2(new_n1371), .A3(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT63), .ZN(new_n1375));
  OR2_X1    g1175(.A1(new_n1343), .A2(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT61), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1361), .A2(new_n1377), .ZN(new_n1378));
  AOI21_X1  g1178(.A(new_n1378), .B1(new_n1375), .B2(new_n1343), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1374), .A2(new_n1376), .A3(new_n1379), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1363), .A2(new_n1380), .ZN(G405));
  NAND2_X1  g1181(.A1(G375), .A2(new_n1300), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1382), .A2(new_n1316), .ZN(new_n1383));
  OR2_X1    g1183(.A1(new_n1383), .A2(new_n1330), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1383), .A2(new_n1330), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1384), .A2(new_n1385), .ZN(new_n1386));
  XNOR2_X1  g1186(.A(new_n1386), .B(new_n1362), .ZN(G402));
endmodule


