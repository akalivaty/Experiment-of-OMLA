//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n458), .B1(new_n448), .B2(new_n454), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT66), .B(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT67), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n464), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  OAI21_X1  g049(.A(G137), .B1(new_n462), .B2(new_n463), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT66), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n474), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n467), .A2(new_n469), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n482), .A2(new_n461), .A3(KEYINPUT68), .A4(G137), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n466), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G101), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n473), .A2(new_n486), .ZN(G160));
  NOR2_X1   g062(.A1(new_n462), .A2(new_n463), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(new_n461), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n461), .C2(G112), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n488), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n464), .A2(new_n470), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n461), .A2(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT4), .A4(G138), .ZN(new_n499));
  NAND2_X1  g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(new_n482), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT69), .A2(G114), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT69), .A2(G114), .ZN(new_n504));
  OAI21_X1  g079(.A(G2105), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n476), .A2(G102), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G2104), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n498), .A2(new_n502), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT70), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT70), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT71), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT6), .B1(new_n517), .B2(new_n518), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n523), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n514), .B1(new_n524), .B2(new_n526), .ZN(new_n528));
  AOI22_X1  g103(.A1(G50), .A2(new_n527), .B1(new_n528), .B2(G88), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n522), .A2(new_n529), .ZN(G166));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  OR3_X1    g106(.A1(new_n514), .A2(KEYINPUT72), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  OAI21_X1  g109(.A(KEYINPUT72), .B1(new_n514), .B2(new_n531), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(G89), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  INV_X1    g113(.A(new_n527), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(G168));
  OR2_X1    g116(.A1(KEYINPUT5), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(KEYINPUT5), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n519), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n527), .A2(G52), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n528), .A2(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  AOI22_X1  g125(.A1(new_n544), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n519), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n527), .A2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n528), .A2(G81), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  INV_X1    g138(.A(G78), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n514), .A2(new_n563), .B1(new_n564), .B2(new_n523), .ZN(new_n565));
  AOI22_X1  g140(.A1(G91), .A2(new_n528), .B1(new_n565), .B2(G651), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT6), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT70), .ZN(new_n568));
  INV_X1    g143(.A(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(KEYINPUT70), .A2(G651), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g147(.A(G53), .B(G543), .C1(new_n572), .C2(new_n525), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n527), .B2(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n566), .B1(new_n574), .B2(new_n576), .ZN(G299));
  XNOR2_X1  g152(.A(new_n540), .B(KEYINPUT73), .ZN(G286));
  NAND2_X1  g153(.A1(new_n522), .A2(new_n529), .ZN(G303));
  NAND2_X1  g154(.A1(new_n528), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n527), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n544), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n544), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n519), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n514), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n589), .A2(KEYINPUT74), .A3(new_n520), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(G48), .A2(new_n527), .B1(new_n528), .B2(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n528), .A2(G85), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n544), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(KEYINPUT75), .B(G47), .ZN(new_n596));
  OAI221_X1 g171(.A(new_n594), .B1(new_n519), .B2(new_n595), .C1(new_n539), .C2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n528), .A2(G92), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT10), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n544), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n569), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n605));
  OAI21_X1  g180(.A(G54), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT77), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n598), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n598), .B1(new_n608), .B2(G868), .ZN(G321));
  AOI21_X1  g185(.A(new_n563), .B1(new_n542), .B2(new_n543), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n564), .A2(new_n523), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n544), .B1(new_n572), .B2(new_n525), .ZN(new_n614));
  INV_X1    g189(.A(G91), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n527), .A2(new_n575), .A3(G53), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT78), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G868), .B2(G286), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT79), .ZN(G297));
  XNOR2_X1  g198(.A(new_n622), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n608), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n608), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n556), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(KEYINPUT81), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(KEYINPUT81), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g207(.A1(new_n464), .A2(new_n470), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(new_n484), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n489), .A2(G123), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n643), .B(new_n644), .C1(new_n461), .C2(G111), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n492), .A2(G135), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n640), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n638), .A2(new_n639), .A3(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2430), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(KEYINPUT85), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(KEYINPUT85), .ZN(new_n659));
  OAI22_X1  g234(.A1(new_n658), .A2(new_n659), .B1(new_n654), .B2(new_n655), .ZN(new_n660));
  XOR2_X1   g235(.A(G2443), .B(G2446), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2451), .B(G2454), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT84), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT86), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  INV_X1    g254(.A(new_n675), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n676), .B1(new_n682), .B2(new_n673), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n674), .B2(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n674), .A2(new_n677), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n680), .B1(new_n685), .B2(KEYINPUT17), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n679), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(new_n650), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2100), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(new_n693), .ZN(new_n699));
  INV_X1    g274(.A(new_n694), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n691), .B2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(new_n701), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n696), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT88), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT89), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1981), .B(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n707), .B(new_n711), .ZN(G229));
  XOR2_X1   g287(.A(KEYINPUT31), .B(G11), .Z(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G28), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(KEYINPUT96), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n715), .B2(G28), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(KEYINPUT96), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n713), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT90), .B(G29), .Z(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n649), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G1966), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(G21), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n540), .B2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n722), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  NOR2_X1   g303(.A1(G171), .A2(new_n724), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G5), .B2(new_n724), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n727), .B1(new_n728), .B2(new_n730), .C1(new_n723), .C2(new_n726), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT97), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n633), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n461), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n734), .B2(new_n733), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n492), .A2(G139), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT25), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G33), .B(new_n742), .S(G29), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2072), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n714), .A2(G32), .ZN(new_n745));
  AOI22_X1  g320(.A1(G129), .A2(new_n489), .B1(new_n492), .B2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT26), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n749), .A2(new_n750), .B1(G105), .B2(new_n484), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n745), .B1(new_n753), .B2(new_n714), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n721), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(G27), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n757), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n756), .B1(G2078), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n759), .ZN(new_n761));
  INV_X1    g336(.A(G2078), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT24), .B(G34), .Z(new_n763));
  NOR2_X1   g338(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G160), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n761), .A2(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n730), .A2(new_n728), .B1(new_n765), .B2(G2084), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n760), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n744), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n732), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(KEYINPUT98), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n732), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n724), .A2(G4), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n608), .B2(new_n724), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1348), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n724), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G1956), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n721), .A2(G26), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT28), .Z(new_n785));
  AOI22_X1  g360(.A1(G128), .A2(new_n489), .B1(new_n492), .B2(G140), .ZN(new_n786));
  OAI221_X1 g361(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n461), .C2(G116), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n785), .B1(new_n788), .B2(G29), .ZN(new_n789));
  INV_X1    g364(.A(G2067), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n757), .A2(G35), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n757), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G2090), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G16), .A2(G19), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n556), .B2(G16), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT94), .B(G1341), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n797), .B(new_n801), .C1(new_n796), .C2(new_n795), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n778), .A2(new_n783), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n773), .A2(new_n775), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT93), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(KEYINPUT36), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n721), .A2(G25), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT91), .Z(new_n808));
  AOI22_X1  g383(.A1(G119), .A2(new_n489), .B1(new_n492), .B2(G131), .ZN(new_n809));
  OAI221_X1 g384(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n461), .C2(G107), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n808), .B1(new_n811), .B2(new_n757), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(G16), .A2(G24), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G290), .B2(new_n724), .ZN(new_n816));
  INV_X1    g391(.A(G1986), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n814), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(G16), .A2(G22), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G166), .B2(G16), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(G1971), .Z(new_n824));
  MUX2_X1   g399(.A(G6), .B(G305), .S(G16), .Z(new_n825));
  XOR2_X1   g400(.A(KEYINPUT32), .B(G1981), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n724), .A2(G23), .ZN(new_n828));
  INV_X1    g403(.A(G288), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n724), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT33), .B(G1976), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n824), .A2(new_n827), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT92), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n824), .A2(new_n835), .A3(new_n827), .A4(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT34), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n821), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(KEYINPUT34), .A3(new_n836), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n806), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n805), .A2(KEYINPUT36), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n804), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n839), .A2(new_n805), .A3(KEYINPUT36), .A4(new_n840), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT100), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n842), .ZN(new_n846));
  INV_X1    g421(.A(new_n804), .ZN(new_n847));
  AND4_X1   g422(.A1(KEYINPUT100), .A2(new_n846), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n848), .ZN(G311));
  NAND2_X1  g424(.A1(new_n843), .A2(new_n844), .ZN(G150));
  NAND2_X1  g425(.A1(new_n527), .A2(G55), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n528), .A2(G93), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n544), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n851), .B(new_n852), .C1(new_n519), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n608), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n555), .B(new_n854), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT102), .Z(new_n863));
  INV_X1    g438(.A(G860), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n856), .B1(new_n863), .B2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(new_n635), .B(new_n811), .ZN(new_n867));
  AOI22_X1  g442(.A1(G130), .A2(new_n489), .B1(new_n492), .B2(G142), .ZN(new_n868));
  OAI221_X1 g443(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n461), .C2(G118), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n867), .B(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n788), .B(new_n752), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n509), .B(KEYINPUT103), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n742), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n873), .B(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(G160), .B(G162), .Z(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(new_n649), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(G37), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n879), .B2(new_n876), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g457(.A1(new_n854), .A2(G868), .ZN(new_n883));
  XNOR2_X1  g458(.A(G303), .B(G305), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G288), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n887));
  INV_X1    g462(.A(new_n858), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n627), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n607), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(G299), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n607), .A2(new_n619), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n890), .A2(KEYINPUT104), .A3(G299), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT41), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n894), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n889), .A2(new_n900), .A3(KEYINPUT105), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n627), .B(new_n858), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT105), .B1(new_n889), .B2(new_n900), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n887), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n904), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n909), .A2(KEYINPUT42), .A3(new_n906), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n886), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n905), .A2(new_n887), .A3(new_n907), .ZN(new_n912));
  INV_X1    g487(.A(new_n886), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n909), .B2(new_n906), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n883), .B1(new_n916), .B2(G868), .ZN(G295));
  AOI21_X1  g492(.A(new_n883), .B1(new_n916), .B2(G868), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  INV_X1    g494(.A(new_n903), .ZN(new_n920));
  NAND2_X1  g495(.A1(G286), .A2(G171), .ZN(new_n921));
  NAND2_X1  g496(.A1(G168), .A2(G301), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n888), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n924), .A2(KEYINPUT106), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n858), .A3(new_n922), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(KEYINPUT106), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n920), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n926), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n900), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G37), .B1(new_n931), .B2(new_n886), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n886), .B(KEYINPUT107), .Z(new_n933));
  NAND2_X1  g508(.A1(new_n897), .A2(KEYINPUT41), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n927), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n920), .B1(new_n935), .B2(new_n929), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n898), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n919), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n900), .A2(new_n929), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n925), .A2(new_n927), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n886), .B(new_n940), .C1(new_n941), .C2(new_n920), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n933), .B1(new_n928), .B2(new_n930), .ZN(new_n944));
  AND4_X1   g519(.A1(new_n919), .A2(new_n942), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT44), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT43), .B1(new_n932), .B2(new_n938), .ZN(new_n948));
  AND4_X1   g523(.A1(KEYINPUT43), .A2(new_n942), .A3(new_n943), .A4(new_n944), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n946), .A2(new_n950), .ZN(G397));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n509), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n473), .ZN(new_n956));
  INV_X1    g531(.A(new_n486), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n957), .A3(G40), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(G1996), .A3(new_n752), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT108), .Z(new_n961));
  NOR3_X1   g536(.A1(new_n955), .A2(G1996), .A3(new_n958), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n753), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n788), .A2(G2067), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n786), .A2(new_n790), .A3(new_n787), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n959), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT109), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n811), .B(new_n813), .Z(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n959), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(G290), .B(G1986), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n959), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT63), .ZN(new_n975));
  INV_X1    g550(.A(G40), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n473), .A2(new_n486), .A3(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n464), .A2(new_n470), .A3(G138), .A4(new_n461), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n978), .A2(new_n495), .B1(G2104), .B2(new_n507), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n979), .B2(new_n502), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(G8), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n983));
  OAI211_X1 g558(.A(G48), .B(G543), .C1(new_n572), .C2(new_n525), .ZN(new_n984));
  INV_X1    g559(.A(G86), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n614), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n528), .A2(G86), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(KEYINPUT114), .A3(new_n984), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n988), .A2(new_n990), .B1(new_n520), .B2(new_n589), .ZN(new_n991));
  INV_X1    g566(.A(G1981), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n983), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n591), .A2(new_n992), .A3(new_n592), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n591), .A2(KEYINPUT113), .A3(new_n592), .A4(new_n992), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n589), .A2(new_n520), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n989), .A2(new_n984), .A3(KEYINPUT114), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT114), .B1(new_n989), .B2(new_n984), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1002), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n993), .A2(new_n998), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n982), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n993), .A2(new_n998), .A3(KEYINPUT49), .A4(new_n1003), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G303), .A2(G8), .ZN(new_n1012));
  XOR2_X1   g587(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n1013));
  XNOR2_X1  g588(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT110), .B(G1971), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n958), .B1(new_n953), .B2(new_n954), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n952), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT117), .B(new_n977), .C1(new_n980), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n980), .A2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT117), .B1(new_n1024), .B2(new_n977), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1019), .B1(new_n1026), .B2(new_n796), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1015), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1020), .B1(new_n509), .B2(new_n952), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n958), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1022), .ZN(new_n1032));
  OAI22_X1  g607(.A1(new_n1019), .A2(KEYINPUT111), .B1(new_n1032), .B2(G2090), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1016), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(KEYINPUT111), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(G8), .B(new_n1014), .C1(new_n1033), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n982), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1039), .B(new_n1041), .C1(new_n1040), .C2(G288), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G288), .A2(new_n1040), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n982), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1011), .A2(new_n1029), .A3(new_n1038), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1018), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n980), .A2(KEYINPUT118), .A3(KEYINPUT45), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1017), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n723), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1053), .A2(new_n958), .A3(new_n1030), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n767), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1028), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(G286), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n975), .B1(new_n1047), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1007), .B(new_n1008), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1045), .B1(new_n1060), .B2(new_n1006), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1057), .A2(new_n975), .A3(G286), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1015), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1061), .A2(new_n1062), .A3(new_n1038), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1011), .A2(new_n1040), .A3(new_n829), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n998), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1038), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1068), .A2(new_n1039), .B1(new_n1069), .B2(new_n1061), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n782), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1071));
  NOR2_X1   g646(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n617), .A2(new_n618), .ZN(new_n1077));
  AOI211_X1 g652(.A(KEYINPUT120), .B(new_n1076), .C1(new_n1077), .C2(new_n566), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1076), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(G299), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1073), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT120), .B1(new_n619), .B2(new_n1076), .ZN(new_n1083));
  NAND3_X1  g658(.A1(G299), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1072), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT56), .B(G2072), .Z(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1017), .A2(new_n1018), .A3(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1071), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1086), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1053), .B1(new_n1031), .B2(KEYINPUT117), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1030), .B2(new_n958), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1956), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1089), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1091), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1348), .B1(new_n1031), .B2(new_n1022), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n977), .A2(new_n980), .A3(new_n790), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n890), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1090), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n1103));
  INV_X1    g678(.A(G1996), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n955), .A2(new_n1104), .A3(new_n977), .A4(new_n1018), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n981), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(KEYINPUT121), .A3(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1103), .B1(new_n1112), .B2(new_n556), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1105), .A2(KEYINPUT121), .A3(new_n1107), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT121), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1103), .B(new_n556), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT59), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n556), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT122), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1121), .A3(new_n1116), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1086), .B1(new_n1071), .B2(new_n1089), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1090), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1071), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1097), .A2(KEYINPUT61), .A3(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n607), .B(new_n1099), .C1(new_n1054), .C2(G1348), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1101), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n607), .A2(KEYINPUT60), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1130), .A2(KEYINPUT60), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1126), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1102), .B1(new_n1123), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(G171), .B1(new_n1032), .B2(new_n728), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1017), .A2(new_n762), .A3(new_n1018), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1017), .A2(KEYINPUT53), .A3(new_n762), .A4(new_n1018), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT124), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1032), .A2(new_n728), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1138), .A2(G2078), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1017), .A2(new_n1049), .A3(new_n1050), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1139), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(G171), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1136), .A2(new_n1139), .A3(new_n1148), .A4(new_n1140), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1142), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1139), .A2(new_n1143), .A3(new_n1140), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1151), .B1(new_n1154), .B2(new_n1136), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1150), .A2(new_n1151), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  AND4_X1   g731(.A1(new_n1029), .A2(new_n1011), .A3(new_n1038), .A4(new_n1046), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n540), .A2(G8), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1057), .A2(KEYINPUT51), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT51), .ZN(new_n1160));
  NOR2_X1   g735(.A1(G168), .A2(new_n1028), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1056), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1056), .A2(KEYINPUT123), .A3(new_n540), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT123), .B1(new_n1056), .B2(new_n540), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1159), .B(new_n1162), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1156), .A2(new_n1157), .A3(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1066), .B(new_n1070), .C1(new_n1135), .C2(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1167), .A2(KEYINPUT125), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1047), .A2(new_n1147), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1165), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1165), .A2(new_n1170), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(new_n1167), .B2(KEYINPUT125), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n974), .B1(new_n1168), .B2(new_n1174), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n972), .A2(KEYINPUT127), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n972), .A2(KEYINPUT127), .ZN(new_n1177));
  NOR2_X1   g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n959), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT48), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1176), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n969), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n809), .A2(new_n810), .A3(new_n813), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n965), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n959), .ZN(new_n1185));
  NAND2_X1  g760(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1186));
  INV_X1    g761(.A(new_n962), .ZN(new_n1187));
  NOR2_X1   g762(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n959), .B1(new_n752), .B2(new_n966), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1189), .B(new_n1190), .C1(new_n1187), .C2(new_n1186), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT47), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1181), .A2(new_n1185), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1175), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g769(.A1(G229), .A2(new_n459), .A3(G227), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n881), .A2(new_n671), .A3(new_n1196), .ZN(new_n1197));
  NOR3_X1   g771(.A1(new_n1197), .A2(new_n948), .A3(new_n949), .ZN(G308));
  OR3_X1    g772(.A1(new_n1197), .A2(new_n948), .A3(new_n949), .ZN(G225));
endmodule


