//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT67), .A2(G237), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT67), .A2(G237), .ZN(new_n189));
  AOI21_X1  g003(.A(G953), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  AOI21_X1  g004(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT67), .A2(G237), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT67), .A2(G237), .ZN(new_n194));
  OAI211_X1 g008(.A(G214), .B(new_n192), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n191), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT93), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT18), .A3(G131), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n195), .A2(new_n196), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n204), .A2(new_n199), .A3(KEYINPUT18), .A4(G131), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT78), .ZN(new_n210));
  OR3_X1    g024(.A1(new_n208), .A2(KEYINPUT78), .A3(G140), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT94), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT94), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G146), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n207), .A2(new_n209), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT80), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n201), .B(new_n205), .C1(new_n217), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT95), .B1(new_n198), .B2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT95), .A4(new_n223), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT96), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n204), .B2(G131), .ZN(new_n228));
  AOI211_X1 g042(.A(KEYINPUT96), .B(new_n223), .C1(new_n202), .C2(new_n203), .ZN(new_n229));
  OAI22_X1  g043(.A1(new_n224), .A2(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT17), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT96), .B1(new_n198), .B2(new_n223), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n204), .A2(new_n227), .A3(G131), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(KEYINPUT17), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT16), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT16), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n207), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(G146), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n219), .B1(new_n235), .B2(new_n237), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n234), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n222), .B1(new_n231), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G113), .B(G122), .ZN(new_n244));
  INV_X1    g058(.A(G104), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n246), .B(new_n222), .C1(new_n231), .C2(new_n242), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G902), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n187), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n210), .A2(KEYINPUT94), .A3(new_n211), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT94), .B1(new_n210), .B2(new_n211), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT19), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(KEYINPUT19), .B2(new_n218), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n240), .B1(new_n256), .B2(new_n219), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n220), .B(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n259), .A2(new_n216), .B1(new_n198), .B2(new_n200), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n257), .A2(new_n230), .B1(new_n205), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n246), .B1(new_n261), .B2(KEYINPUT97), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT95), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n263), .B1(new_n204), .B2(G131), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n232), .A2(new_n233), .B1(new_n264), .B2(new_n225), .ZN(new_n265));
  INV_X1    g079(.A(new_n240), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n218), .A2(KEYINPUT19), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n214), .A2(new_n215), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(KEYINPUT19), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n266), .B1(new_n269), .B2(G146), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n222), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT97), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n222), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n234), .A2(new_n241), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT17), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n265), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n262), .A2(new_n273), .B1(new_n278), .B2(new_n246), .ZN(new_n279));
  NOR2_X1   g093(.A1(G475), .A2(G902), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT98), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT20), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(KEYINPUT97), .B(new_n222), .C1(new_n265), .C2(new_n270), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n247), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n257), .A2(new_n230), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT97), .B1(new_n285), .B2(new_n222), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n249), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT20), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n281), .B(KEYINPUT99), .Z(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n252), .B1(new_n282), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT9), .B(G234), .ZN(new_n292));
  INV_X1    g106(.A(G217), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n292), .A2(new_n293), .A3(G953), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n196), .A2(G128), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT101), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT13), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G128), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G143), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n298), .B(new_n300), .C1(new_n297), .C2(new_n295), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n302));
  OAI21_X1  g116(.A(G134), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n295), .A2(new_n300), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G122), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G116), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT100), .ZN(new_n309));
  INV_X1    g123(.A(G107), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G122), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n310), .B1(new_n309), .B2(new_n312), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n303), .B(new_n306), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n304), .B(new_n305), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT14), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n312), .B(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n309), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n317), .B(new_n313), .C1(new_n320), .C2(new_n310), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n294), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n316), .A2(new_n321), .A3(new_n294), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n251), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT15), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G478), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(G478), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n251), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G952), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G953), .ZN(new_n334));
  NAND2_X1  g148(.A1(G234), .A2(G237), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT21), .B(G898), .Z(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(G902), .A3(G953), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n291), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G214), .B1(G237), .B2(G902), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n245), .A2(KEYINPUT85), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT85), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n343), .B1(new_n347), .B2(new_n310), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n346), .A3(G107), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n343), .A2(new_n310), .A3(G104), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G101), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT85), .B(G104), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT3), .B1(new_n353), .B2(G107), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n245), .A2(KEYINPUT3), .A3(G107), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n353), .B2(G107), .ZN(new_n356));
  INV_X1    g170(.A(G101), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n352), .A2(KEYINPUT4), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n360));
  INV_X1    g174(.A(G119), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G116), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n311), .A2(G119), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT2), .B(G113), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G116), .B(G119), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT2), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G113), .ZN(new_n369));
  INV_X1    g183(.A(G113), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(KEYINPUT2), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n367), .B(KEYINPUT66), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n364), .A2(new_n365), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n376), .B(G101), .C1(new_n348), .C2(new_n351), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n362), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT5), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n370), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n367), .A2(KEYINPUT5), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT90), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT90), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n373), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n353), .A2(G107), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n310), .A2(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(G101), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n358), .A2(new_n390), .ZN(new_n391));
  OAI22_X1  g205(.A1(new_n359), .A2(new_n378), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G110), .B(G122), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  OAI221_X1 g209(.A(new_n393), .B1(new_n387), .B2(new_n391), .C1(new_n359), .C2(new_n378), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(KEYINPUT6), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT6), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n398), .A3(new_n394), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT64), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n196), .B2(G146), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n196), .A2(G146), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n219), .A2(KEYINPUT64), .A3(G143), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(KEYINPUT0), .A2(G128), .ZN(new_n405));
  NOR2_X1   g219(.A1(KEYINPUT0), .A2(G128), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G143), .B(G146), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n405), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n208), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G128), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n299), .A2(KEYINPUT1), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n404), .A2(new_n414), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G125), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n192), .A2(G224), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n418), .B(new_n419), .Z(new_n420));
  NAND3_X1  g234(.A1(new_n397), .A2(new_n399), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT7), .B(new_n419), .C1(new_n412), .C2(new_n417), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n404), .A2(new_n407), .B1(new_n409), .B2(new_n405), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G125), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(KEYINPUT7), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n424), .B(new_n425), .C1(G125), .C2(new_n416), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n358), .A2(new_n390), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT91), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n381), .B1(new_n382), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT91), .B1(new_n367), .B2(KEYINPUT5), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n373), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n393), .B(KEYINPUT8), .Z(new_n434));
  INV_X1    g248(.A(new_n387), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n391), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n427), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n437), .B2(new_n396), .ZN(new_n438));
  OAI21_X1  g252(.A(G210), .B1(G237), .B2(G902), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n421), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n421), .B2(new_n438), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(KEYINPUT92), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT92), .ZN(new_n443));
  AOI211_X1 g257(.A(new_n443), .B(new_n439), .C1(new_n421), .C2(new_n438), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n342), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n341), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G472), .ZN(new_n447));
  INV_X1    g261(.A(G137), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT65), .B1(new_n448), .B2(G134), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT65), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n305), .A3(G137), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n448), .A2(KEYINPUT11), .A3(G134), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT11), .B1(new_n448), .B2(G134), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n223), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT11), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n305), .B2(G137), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n448), .A2(KEYINPUT11), .A3(G134), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n449), .A2(new_n458), .A3(new_n451), .A4(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G131), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n423), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n404), .A2(new_n414), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n409), .A2(new_n415), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n452), .A2(new_n455), .A3(new_n223), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n305), .A2(G137), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n448), .A2(G134), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n223), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n462), .A2(new_n463), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n463), .B1(new_n462), .B2(new_n472), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n375), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n462), .A2(new_n472), .A3(new_n374), .A4(new_n373), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n190), .A2(G210), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT27), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT27), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n190), .A2(new_n479), .A3(G210), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT26), .B(G101), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n478), .B2(new_n480), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n475), .A2(KEYINPUT68), .A3(new_n476), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT31), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT69), .B1(new_n483), .B2(new_n484), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n478), .A2(new_n480), .ZN(new_n490));
  INV_X1    g304(.A(new_n481), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n482), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT28), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n460), .A2(G131), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n411), .B1(new_n467), .B2(new_n497), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n461), .A2(new_n416), .A3(new_n470), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n375), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n496), .B1(new_n500), .B2(new_n476), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n476), .A2(new_n496), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n495), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n486), .B2(KEYINPUT31), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n447), .B(new_n251), .C1(new_n488), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT70), .ZN(new_n506));
  INV_X1    g320(.A(new_n476), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT30), .B1(new_n498), .B2(new_n499), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n462), .A2(new_n472), .A3(new_n463), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n510), .B2(new_n375), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT31), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n511), .A2(KEYINPUT68), .A3(new_n512), .A4(new_n485), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n487), .A3(new_n503), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT70), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n447), .A4(new_n251), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n506), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n501), .A2(new_n502), .ZN(new_n519));
  INV_X1    g333(.A(new_n485), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT29), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(G902), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n495), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT72), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n526));
  NOR4_X1   g340(.A1(new_n495), .A2(new_n501), .A3(new_n502), .A4(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT73), .B1(new_n511), .B2(new_n485), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n475), .A2(new_n476), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT73), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n520), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n521), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n523), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G472), .ZN(new_n535));
  INV_X1    g349(.A(new_n505), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT32), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n518), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT22), .B(G137), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n259), .A2(new_n266), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G110), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT74), .B1(new_n299), .B2(G119), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT74), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n361), .A3(G128), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n299), .A2(G119), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT75), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n545), .A2(new_n547), .B1(G119), .B2(new_n299), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n544), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n555), .A2(KEYINPUT79), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n549), .A2(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n549), .A2(KEYINPUT77), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT23), .B1(new_n299), .B2(G119), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n299), .A2(KEYINPUT23), .A3(G119), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT76), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G110), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n555), .A2(KEYINPUT79), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n542), .B1(new_n556), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n560), .A2(new_n562), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G110), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n552), .A2(new_n554), .A3(new_n544), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n569), .C1(new_n239), .C2(new_n240), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n541), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n221), .A2(new_n240), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n563), .A2(new_n564), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n550), .A2(new_n551), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT79), .B(new_n543), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n555), .A2(KEYINPUT79), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n573), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n541), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n570), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n572), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n583), .A2(KEYINPUT81), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(KEYINPUT81), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n293), .B1(G234), .B2(new_n251), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(G902), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT82), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT25), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n583), .B2(new_n251), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n566), .A2(new_n571), .A3(new_n541), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n581), .B1(new_n580), .B2(new_n570), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n590), .B(new_n251), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n595), .A2(new_n587), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n586), .A2(new_n589), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G221), .B1(new_n292), .B2(G902), .ZN(new_n598));
  XOR2_X1   g412(.A(new_n598), .B(KEYINPUT83), .Z(new_n599));
  INV_X1    g413(.A(G469), .ZN(new_n600));
  XNOR2_X1  g414(.A(G110), .B(G140), .ZN(new_n601));
  INV_X1    g415(.A(G227), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G953), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n601), .B(new_n603), .Z(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n456), .A2(new_n461), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n466), .A2(KEYINPUT10), .ZN(new_n607));
  INV_X1    g421(.A(new_n414), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n465), .B1(new_n608), .B2(new_n409), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n358), .A2(new_n390), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT87), .B(KEYINPUT10), .Z(new_n611));
  AOI22_X1  g425(.A1(new_n428), .A2(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n377), .A2(new_n423), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n359), .A2(KEYINPUT86), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT86), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n357), .B1(new_n354), .B2(new_n356), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n411), .B1(new_n616), .B2(new_n376), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n352), .A2(new_n358), .A3(KEYINPUT4), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n606), .B(new_n612), .C1(new_n614), .C2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT86), .B1(new_n359), .B2(new_n613), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n617), .A2(new_n615), .A3(new_n618), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n606), .B1(new_n624), .B2(new_n612), .ZN(new_n625));
  OAI211_X1 g439(.A(KEYINPUT89), .B(new_n605), .C1(new_n621), .C2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n606), .ZN(new_n627));
  INV_X1    g441(.A(new_n610), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n466), .B1(new_n358), .B2(new_n390), .ZN(new_n629));
  OAI211_X1 g443(.A(KEYINPUT12), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT88), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n610), .B1(new_n428), .B2(new_n466), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT88), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT12), .A4(new_n627), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n632), .A2(new_n627), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n631), .B(new_n634), .C1(new_n635), .C2(KEYINPUT12), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n620), .A3(new_n604), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n626), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n612), .B1(new_n614), .B2(new_n619), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n627), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n620), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT89), .B1(new_n641), .B2(new_n605), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n600), .B(new_n251), .C1(new_n638), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n636), .A2(new_n620), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n604), .B(KEYINPUT84), .Z(new_n645));
  AND2_X1   g459(.A1(new_n620), .A2(new_n604), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n644), .A2(new_n645), .B1(new_n646), .B2(new_n640), .ZN(new_n647));
  OAI21_X1  g461(.A(G469), .B1(new_n647), .B2(G902), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n599), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n446), .A2(new_n538), .A3(new_n597), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G101), .ZN(G3));
  INV_X1    g465(.A(new_n649), .ZN(new_n652));
  INV_X1    g466(.A(new_n597), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n514), .A2(new_n251), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(G472), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n506), .A2(new_n656), .A3(new_n516), .ZN(new_n657));
  INV_X1    g471(.A(new_n249), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n275), .A2(new_n277), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n246), .B1(new_n659), .B2(new_n222), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n251), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G475), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n663));
  INV_X1    g477(.A(new_n281), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n288), .B1(new_n287), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n662), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n324), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n322), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(KEYINPUT33), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(KEYINPUT33), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n325), .A2(new_n669), .A3(KEYINPUT33), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(G478), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(G902), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n674), .A2(new_n676), .B1(new_n675), .B2(new_n326), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n666), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n440), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n339), .B(new_n342), .C1(new_n680), .C2(new_n441), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n654), .A2(new_n657), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT34), .B(G104), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G6));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n665), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n273), .A2(new_n247), .A3(new_n283), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n281), .B1(new_n688), .B2(new_n249), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT103), .B1(new_n689), .B2(new_n288), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n287), .A2(new_n288), .A3(new_n664), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n681), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n252), .A2(new_n332), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n654), .A2(new_n695), .A3(new_n657), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT35), .B(G107), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  NAND2_X1  g512(.A1(new_n580), .A2(new_n570), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n589), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n595), .A2(new_n587), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(new_n591), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n446), .A2(new_n649), .A3(new_n657), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  OR2_X1    g521(.A1(new_n338), .A2(G900), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n336), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n691), .B1(new_n665), .B2(new_n686), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n689), .A2(KEYINPUT103), .A3(new_n288), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n694), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n342), .ZN(new_n714));
  INV_X1    g528(.A(new_n441), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n714), .B1(new_n715), .B2(new_n440), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n716), .A2(new_n704), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n713), .A2(new_n538), .A3(new_n649), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  XNOR2_X1  g533(.A(new_n709), .B(KEYINPUT39), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n649), .A2(KEYINPUT105), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT105), .B1(new_n649), .B2(new_n720), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT40), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n723), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT40), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n721), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n524), .B1(new_n476), .B2(new_n500), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n530), .A2(new_n520), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n251), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G472), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n518), .A2(new_n537), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n331), .A2(new_n342), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n291), .A2(new_n704), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n442), .A2(new_n444), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n442), .B2(new_n444), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n732), .A2(new_n734), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n724), .A2(new_n727), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT106), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n724), .A2(new_n727), .A3(new_n743), .A4(new_n740), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n196), .ZN(G45));
  INV_X1    g560(.A(new_n709), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n291), .A2(new_n677), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n538), .A3(new_n649), .A4(new_n717), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G146), .ZN(G48));
  OAI21_X1  g564(.A(new_n251), .B1(new_n638), .B2(new_n642), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  INV_X1    g566(.A(new_n599), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n752), .A2(new_n753), .A3(new_n643), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n682), .A2(new_n754), .A3(new_n597), .A4(new_n538), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n755), .A2(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(KEYINPUT107), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT41), .B(G113), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G15));
  NAND4_X1  g574(.A1(new_n695), .A2(new_n597), .A3(new_n538), .A4(new_n754), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G116), .ZN(G18));
  INV_X1    g576(.A(new_n341), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n754), .A2(new_n763), .A3(new_n538), .A4(new_n717), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G119), .ZN(G21));
  AND3_X1   g579(.A1(new_n597), .A2(new_n505), .A3(new_n656), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n680), .A2(new_n441), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n291), .A2(new_n767), .A3(new_n733), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n766), .A2(new_n754), .A3(new_n768), .A4(new_n339), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT108), .B(G122), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G24));
  NAND3_X1  g585(.A1(new_n666), .A2(new_n678), .A3(new_n709), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n656), .A2(new_n704), .A3(new_n505), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n753), .A2(new_n752), .A3(new_n643), .A4(new_n716), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G125), .ZN(G27));
  AND2_X1   g591(.A1(new_n537), .A2(new_n535), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n536), .A2(KEYINPUT32), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n653), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n442), .A2(new_n714), .A3(new_n444), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n649), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(KEYINPUT42), .A3(new_n748), .A4(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n597), .A3(new_n538), .A4(new_n748), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT42), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n784), .B2(KEYINPUT109), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n783), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT110), .B(G131), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G33));
  NAND4_X1  g604(.A1(new_n782), .A2(new_n713), .A3(new_n597), .A4(new_n538), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  NAND2_X1  g606(.A1(new_n291), .A2(new_n678), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT43), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT43), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n291), .A2(new_n795), .A3(new_n678), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n704), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n657), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(KEYINPUT44), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n794), .A3(new_n796), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n781), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n647), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n647), .A2(new_n805), .ZN(new_n807));
  OAI21_X1  g621(.A(G469), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(G469), .A2(G902), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(KEYINPUT46), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n647), .B(new_n805), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n811), .B(G469), .C1(new_n812), .C2(G902), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n813), .A3(new_n643), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n753), .A4(new_n720), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n753), .A3(new_n720), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT111), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n804), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(KEYINPUT112), .B(G137), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n819), .B(new_n820), .ZN(G39));
  NAND2_X1  g635(.A1(new_n653), .A2(new_n781), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n538), .A3(new_n772), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n814), .A2(KEYINPUT47), .A3(new_n753), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT47), .B1(new_n814), .B2(new_n753), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NAND2_X1  g642(.A1(new_n333), .A2(new_n192), .ZN(new_n829));
  INV_X1    g643(.A(new_n336), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n797), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n754), .A2(new_n781), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT120), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n780), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT48), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OR4_X1    g654(.A1(new_n653), .A2(new_n832), .A3(new_n336), .A4(new_n732), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n334), .B1(new_n841), .B2(new_n679), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n797), .A2(new_n830), .A3(new_n766), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n775), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT48), .B1(new_n837), .B2(new_n838), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n833), .B(new_n834), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT121), .B1(new_n846), .B2(new_n780), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n840), .B(new_n844), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n754), .A2(new_n714), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n738), .A2(new_n739), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT50), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(KEYINPUT119), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n843), .A2(new_n852), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n857), .B(new_n858), .Z(new_n859));
  INV_X1    g673(.A(new_n826), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n824), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n752), .A2(new_n643), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n599), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n781), .B(new_n843), .C1(new_n861), .C2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n656), .A2(new_n505), .A3(new_n704), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n846), .A2(new_n865), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n841), .A2(new_n666), .A3(new_n678), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n859), .A2(new_n864), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n848), .B1(new_n849), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n849), .B2(new_n868), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n538), .A2(new_n717), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n652), .A2(new_n712), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n871), .A2(new_n872), .B1(new_n775), .B2(new_n774), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n798), .A2(new_n709), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n768), .A2(new_n732), .A3(new_n649), .A4(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n873), .A2(KEYINPUT52), .A3(new_n749), .A4(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n718), .A2(new_n776), .A3(new_n749), .A4(new_n876), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n331), .A2(KEYINPUT114), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n328), .A2(new_n883), .A3(new_n330), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n747), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n885), .A2(new_n662), .A3(new_n704), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n782), .A2(new_n538), .A3(new_n692), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT115), .B1(new_n782), .B2(new_n774), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n290), .B1(new_n689), .B2(new_n288), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n677), .B1(new_n889), .B2(new_n662), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n865), .A2(new_n890), .A3(new_n709), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n643), .A2(new_n648), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n781), .A2(new_n892), .A3(new_n753), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n791), .B(new_n887), .C1(new_n888), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n654), .A2(new_n657), .ZN(new_n897));
  INV_X1    g711(.A(new_n445), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n889), .A2(new_n662), .A3(new_n882), .A4(new_n884), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n339), .B(new_n898), .C1(new_n900), .C2(new_n890), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n650), .B(new_n705), .C1(new_n897), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n761), .A2(new_n769), .A3(new_n764), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n756), .B2(new_n757), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n881), .A2(new_n788), .A3(new_n903), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT53), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n788), .A2(new_n903), .A3(new_n905), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n878), .A2(new_n879), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n878), .A2(new_n879), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n877), .A2(new_n880), .A3(KEYINPUT117), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n788), .A2(new_n903), .A3(new_n905), .A4(new_n910), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(KEYINPUT54), .B(new_n907), .C1(new_n911), .C2(new_n919), .ZN(new_n920));
  AND4_X1   g734(.A1(KEYINPUT53), .A2(new_n788), .A3(new_n903), .A4(new_n905), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n917), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n906), .A2(new_n908), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n829), .B1(new_n870), .B2(new_n926), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n653), .A2(new_n599), .A3(new_n714), .ZN(new_n928));
  INV_X1    g742(.A(new_n793), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT49), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n928), .B(new_n929), .C1(new_n930), .C2(new_n862), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT113), .ZN(new_n932));
  INV_X1    g746(.A(new_n732), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n854), .B1(new_n930), .B2(new_n862), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n927), .A2(new_n935), .ZN(G75));
  NOR2_X1   g750(.A1(new_n192), .A2(G952), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n921), .A2(new_n917), .B1(new_n908), .B2(new_n906), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n938), .A2(new_n251), .A3(new_n439), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(KEYINPUT56), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n397), .A2(new_n399), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n420), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT55), .Z(new_n943));
  AOI21_X1  g757(.A(new_n937), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(KEYINPUT56), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT122), .B1(new_n938), .B2(new_n251), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n788), .A2(new_n903), .A3(new_n905), .A4(KEYINPUT53), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n915), .B2(new_n916), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n906), .A2(new_n908), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n947), .B(G902), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n945), .B1(new_n952), .B2(new_n439), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n944), .A2(new_n953), .ZN(G51));
  INV_X1    g768(.A(new_n808), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n946), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n638), .A2(new_n642), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT54), .B1(new_n949), .B2(new_n950), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n925), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n809), .B(KEYINPUT57), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n957), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT123), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n956), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n958), .B2(new_n925), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT123), .B1(new_n965), .B2(new_n957), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n937), .B1(new_n964), .B2(new_n966), .ZN(G54));
  NAND4_X1  g781(.A1(new_n946), .A2(new_n951), .A3(KEYINPUT58), .A4(G475), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n968), .A2(new_n279), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n279), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n937), .ZN(G60));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT59), .Z(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n920), .B2(new_n925), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n674), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(KEYINPUT124), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n974), .B2(new_n674), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n976), .A2(new_n973), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n937), .B1(new_n959), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n977), .A2(new_n979), .A3(new_n981), .ZN(G63));
  NAND2_X1  g796(.A1(G217), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT60), .Z(new_n984));
  OAI211_X1 g798(.A(new_n701), .B(new_n984), .C1(new_n949), .C2(new_n950), .ZN(new_n985));
  INV_X1    g799(.A(new_n937), .ZN(new_n986));
  INV_X1    g800(.A(new_n984), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n938), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n985), .B(new_n986), .C1(new_n988), .C2(new_n586), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n989), .A2(KEYINPUT125), .A3(KEYINPUT61), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT61), .B1(new_n989), .B2(KEYINPUT125), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(G66));
  NAND3_X1  g806(.A1(new_n337), .A2(G224), .A3(G953), .ZN(new_n993));
  INV_X1    g807(.A(new_n902), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n905), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n993), .B1(new_n995), .B2(G953), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n941), .B1(G898), .B2(new_n192), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n996), .B(new_n997), .Z(G69));
  XNOR2_X1  g812(.A(new_n510), .B(new_n269), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n873), .A2(new_n749), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n742), .A2(new_n744), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n742), .A2(KEYINPUT62), .A3(new_n1001), .A4(new_n744), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n818), .A2(new_n816), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1007), .A2(new_n781), .A3(new_n803), .A4(new_n800), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n781), .B1(new_n900), .B2(new_n890), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n649), .A2(new_n720), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n597), .A3(new_n538), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1006), .A2(new_n1008), .A3(new_n827), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1000), .B1(new_n1013), .B2(new_n192), .ZN(new_n1014));
  INV_X1    g828(.A(new_n791), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n861), .B2(new_n823), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1008), .A2(new_n1016), .A3(new_n788), .A4(new_n1001), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n780), .A2(new_n768), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1018), .B1(new_n1007), .B2(new_n1020), .ZN(new_n1021));
  AOI211_X1 g835(.A(KEYINPUT127), .B(new_n1019), .C1(new_n818), .C2(new_n816), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n192), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n192), .A2(G900), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n999), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(KEYINPUT126), .B1(new_n1014), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1008), .A2(new_n827), .A3(new_n1012), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1029), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n999), .B1(new_n1030), .B2(G953), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT126), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n827), .A2(new_n1001), .A3(new_n791), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1033), .A2(new_n819), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n1034), .B(new_n788), .C1(new_n1022), .C2(new_n1021), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1025), .B1(new_n1035), .B2(new_n192), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1031), .B(new_n1032), .C1(new_n1036), .C2(new_n999), .ZN(new_n1037));
  INV_X1    g851(.A(G900), .ZN(new_n1038));
  OAI21_X1  g852(.A(G953), .B1(new_n602), .B2(new_n1038), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1028), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1039), .B1(new_n1028), .B2(new_n1037), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1040), .A2(new_n1041), .ZN(G72));
  NOR2_X1   g856(.A1(new_n911), .A2(new_n919), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1043), .B1(KEYINPUT53), .B2(new_n906), .ZN(new_n1044));
  NAND2_X1  g858(.A1(G472), .A2(G902), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n1045), .B(KEYINPUT63), .Z(new_n1046));
  NAND2_X1  g860(.A1(new_n529), .A2(new_n532), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n1044), .B(new_n1046), .C1(new_n1047), .C2(new_n729), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1046), .B1(new_n1013), .B2(new_n995), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1049), .A2(new_n485), .A3(new_n530), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1046), .B1(new_n1035), .B2(new_n995), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n530), .A2(new_n485), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n937), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AND3_X1   g867(.A1(new_n1048), .A2(new_n1050), .A3(new_n1053), .ZN(G57));
endmodule


