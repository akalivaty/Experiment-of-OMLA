//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT82), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(KEYINPUT82), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G107), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n190), .A2(new_n193), .A3(KEYINPUT82), .A4(G104), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT83), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n193), .B2(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n194), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n198), .A2(new_n201), .ZN(new_n204));
  OAI21_X1  g018(.A(G101), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n200), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n211), .A2(KEYINPUT65), .A3(G143), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT65), .B1(new_n211), .B2(G143), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n208), .B(new_n210), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n211), .A2(G143), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n207), .B2(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n211), .A2(KEYINPUT65), .A3(G143), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(G143), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n209), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n214), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n206), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT10), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n195), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n199), .A2(new_n198), .ZN(new_n227));
  OAI21_X1  g041(.A(G101), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT4), .A3(new_n200), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n207), .A2(KEYINPUT64), .A3(G146), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT64), .B1(new_n207), .B2(G146), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n220), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n232), .A2(new_n235), .B1(new_n219), .B2(new_n233), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n237), .B(G101), .C1(new_n226), .C2(new_n227), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n229), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G137), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT11), .A3(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n242), .A2(new_n244), .A3(new_n248), .A4(new_n245), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n207), .A2(G146), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n208), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n207), .A2(KEYINPUT64), .A3(G146), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n251), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n214), .B1(new_n255), .B2(new_n221), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n206), .A2(KEYINPUT10), .A3(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n225), .A2(new_n239), .A3(new_n250), .A4(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G110), .B(G140), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G227), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n200), .A2(new_n205), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  OAI21_X1  g081(.A(G128), .B1(new_n251), .B2(new_n267), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n232), .A2(new_n268), .B1(new_n219), .B2(new_n210), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT84), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT84), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(new_n273), .A3(new_n223), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n247), .A2(new_n249), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n274), .A2(KEYINPUT12), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT12), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n265), .B1(new_n278), .B2(KEYINPUT85), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n276), .B2(new_n277), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n189), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT12), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n266), .A2(new_n272), .A3(new_n269), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n222), .A2(new_n200), .A3(new_n205), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n272), .B1(new_n266), .B2(new_n269), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n283), .B1(new_n287), .B2(new_n250), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n274), .A2(KEYINPUT12), .A3(new_n275), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(KEYINPUT85), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n265), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n281), .A2(new_n290), .A3(new_n189), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n264), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n225), .A2(new_n239), .A3(new_n257), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(new_n275), .ZN(new_n295));
  INV_X1    g109(.A(new_n258), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n187), .B(new_n188), .C1(new_n282), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(G469), .A2(G902), .ZN(new_n300));
  OR3_X1    g114(.A1(new_n295), .A2(new_n296), .A3(new_n293), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n278), .A2(new_n296), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(new_n264), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n303), .A2(new_n187), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT9), .B(G234), .ZN(new_n306));
  OAI21_X1  g120(.A(G221), .B1(new_n306), .B2(G902), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n309));
  INV_X1    g123(.A(G119), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G128), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(G128), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n309), .B(new_n311), .C1(new_n312), .C2(KEYINPUT23), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G110), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT24), .B(G110), .Z(new_n315));
  XNOR2_X1  g129(.A(G119), .B(G128), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G125), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G140), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT77), .A4(KEYINPUT16), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT16), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT16), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(new_n320), .A3(G125), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n211), .B(new_n324), .C1(new_n325), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n321), .A2(new_n323), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n328), .B(new_n327), .C1(new_n332), .C2(new_n326), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n211), .B1(new_n333), .B2(new_n324), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n319), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n324), .B1(new_n325), .B2(new_n329), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G146), .ZN(new_n337));
  OAI22_X1  g151(.A1(new_n313), .A2(G110), .B1(new_n315), .B2(new_n316), .ZN(new_n338));
  XNOR2_X1  g152(.A(G125), .B(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n211), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT78), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT22), .B(G137), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n344), .B(new_n345), .Z(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n344), .B(new_n345), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n335), .A2(new_n341), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT74), .B(G217), .ZN(new_n351));
  INV_X1    g165(.A(G234), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(G902), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT75), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n188), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n358));
  INV_X1    g172(.A(new_n349), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n348), .B1(new_n335), .B2(new_n341), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n188), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n354), .B(KEYINPUT76), .Z(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n358), .B1(new_n350), .B2(new_n188), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n357), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G116), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT67), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT67), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G116), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n369), .A3(G119), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n310), .A2(G116), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT68), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT69), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT2), .B(G113), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n370), .A2(KEYINPUT68), .A3(new_n371), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n370), .A2(KEYINPUT68), .A3(new_n371), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT68), .B1(new_n370), .B2(new_n371), .ZN(new_n380));
  INV_X1    g194(.A(new_n376), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n370), .A3(new_n371), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT69), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n378), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT66), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n243), .A3(G134), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT66), .B1(new_n241), .B2(G137), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n243), .A2(G134), .ZN(new_n390));
  OAI211_X1 g204(.A(G131), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n249), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n256), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n236), .A2(new_n275), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n396), .B1(new_n394), .B2(new_n395), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n386), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n256), .A2(new_n393), .B1(new_n236), .B2(new_n275), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n385), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g215(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n402));
  NOR2_X1   g216(.A1(G237), .A2(G953), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G210), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n402), .B(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT26), .B(G101), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n401), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT31), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n233), .B(new_n208), .C1(new_n212), .C2(new_n213), .ZN(new_n411));
  INV_X1    g225(.A(new_n235), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n255), .B2(new_n412), .ZN(new_n413));
  OAI22_X1  g227(.A1(new_n250), .A2(new_n413), .B1(new_n269), .B2(new_n392), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT69), .A3(new_n383), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n416), .B2(new_n378), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(KEYINPUT30), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n420), .B2(new_n386), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT31), .A3(new_n407), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n414), .A2(new_n416), .A3(new_n378), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n401), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT28), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT28), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n401), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n407), .B(KEYINPUT71), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n410), .A2(new_n422), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(G472), .A2(G902), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT32), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n427), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n426), .B1(new_n401), .B2(new_n423), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n429), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT31), .B1(new_n421), .B2(new_n407), .ZN(new_n437));
  AND4_X1   g251(.A1(KEYINPUT31), .A2(new_n399), .A3(new_n401), .A4(new_n407), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT32), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n431), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n433), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n399), .A2(new_n401), .ZN(new_n443));
  INV_X1    g257(.A(new_n407), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT29), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n445), .B(new_n446), .C1(new_n428), .C2(new_n429), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT72), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n425), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT73), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n427), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n401), .A2(KEYINPUT73), .A3(new_n426), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n435), .A2(KEYINPUT72), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n444), .A2(new_n446), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n449), .A2(new_n453), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n447), .A2(new_n456), .A3(new_n188), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G472), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n365), .B1(new_n442), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n367), .A2(new_n369), .A3(G122), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT93), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT93), .A4(G122), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n366), .A2(G122), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n193), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g281(.A(G107), .B(new_n465), .C1(new_n462), .C2(new_n463), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT94), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT67), .B(G116), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT93), .B1(new_n470), .B2(G122), .ZN(new_n471));
  AND4_X1   g285(.A1(KEYINPUT93), .A2(new_n367), .A3(new_n369), .A4(G122), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G107), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n464), .A2(new_n193), .A3(new_n466), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT95), .B1(new_n207), .B2(G128), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT95), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n209), .A3(G143), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT13), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(new_n241), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n478), .A2(new_n480), .B1(G128), .B2(new_n207), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n469), .A2(new_n477), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n464), .A2(KEYINPUT14), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT14), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n462), .A2(new_n487), .A3(new_n463), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n488), .A3(new_n466), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G107), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n483), .B(G134), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(new_n468), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n351), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n494), .A2(G953), .A3(new_n306), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n485), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n485), .B2(new_n493), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n188), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT15), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(G478), .ZN(new_n500));
  INV_X1    g314(.A(G478), .ZN(new_n501));
  OAI221_X1 g315(.A(new_n188), .B1(KEYINPUT15), .B2(new_n501), .C1(new_n496), .C2(new_n497), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G952), .ZN(new_n505));
  AOI211_X1 g319(.A(G953), .B(new_n505), .C1(G234), .C2(G237), .ZN(new_n506));
  AOI211_X1 g320(.A(new_n188), .B(new_n260), .C1(G234), .C2(G237), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT21), .B(G898), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT20), .ZN(new_n511));
  XNOR2_X1  g325(.A(G113), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n197), .ZN(new_n513));
  INV_X1    g327(.A(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n260), .A3(G214), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(KEYINPUT89), .B2(new_n207), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT89), .B(G143), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT18), .A3(G131), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n332), .A2(G146), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n340), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(KEYINPUT18), .A2(G131), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n516), .B(new_n524), .C1(new_n515), .C2(new_n517), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n340), .A3(KEYINPUT90), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n519), .A2(new_n523), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n517), .A2(new_n515), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT89), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n403), .A2(G214), .B1(new_n530), .B2(G143), .ZN(new_n531));
  OAI21_X1  g345(.A(G131), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n337), .B(new_n330), .C1(new_n528), .C2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n516), .B(new_n248), .C1(new_n515), .C2(new_n517), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n513), .B(new_n527), .C1(new_n533), .C2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT19), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n332), .A2(KEYINPUT91), .A3(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(KEYINPUT91), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n538), .A2(KEYINPUT91), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n339), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n211), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n535), .A2(new_n337), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n527), .A3(KEYINPUT92), .ZN(new_n545));
  INV_X1    g359(.A(new_n513), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT92), .B1(new_n544), .B2(new_n527), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n537), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(G475), .A2(G902), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n511), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n511), .A3(new_n550), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n527), .B1(new_n533), .B2(new_n536), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n546), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n537), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n188), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n552), .A2(new_n553), .B1(G475), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n504), .A2(new_n510), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT87), .ZN(new_n560));
  OAI21_X1  g374(.A(G113), .B1(new_n371), .B2(KEYINPUT5), .ZN(new_n561));
  INV_X1    g375(.A(new_n371), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n470), .B2(G119), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n561), .B1(new_n563), .B2(KEYINPUT5), .ZN(new_n564));
  INV_X1    g378(.A(new_n383), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT5), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n372), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(KEYINPUT87), .B(new_n383), .C1(new_n568), .C2(new_n561), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n569), .A3(new_n206), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n374), .B2(new_n377), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n383), .B(new_n266), .C1(new_n571), .C2(new_n561), .ZN(new_n572));
  XNOR2_X1  g386(.A(G110), .B(G122), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT88), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT88), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n570), .A2(new_n572), .A3(new_n577), .A4(new_n574), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n383), .B(new_n206), .C1(new_n571), .C2(new_n561), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n229), .A2(new_n238), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n580), .B(new_n573), .C1(new_n385), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n269), .A2(new_n322), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n413), .A2(G125), .ZN(new_n584));
  INV_X1    g398(.A(G224), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(G953), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT7), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n583), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n583), .B2(new_n584), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n579), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n580), .B1(new_n385), .B2(new_n581), .ZN(new_n594));
  INV_X1    g408(.A(new_n573), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(KEYINPUT6), .A3(new_n582), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n583), .A2(new_n584), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n586), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT6), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n594), .A2(new_n600), .A3(new_n595), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n597), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G210), .B1(G237), .B2(G902), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n593), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n593), .B2(new_n602), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G214), .B1(G237), .B2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n559), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n308), .A2(new_n459), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  OAI21_X1  g426(.A(G472), .B1(new_n430), .B2(G902), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n430), .B2(new_n432), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n365), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n593), .A2(new_n602), .ZN(new_n616));
  INV_X1    g430(.A(new_n603), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(KEYINPUT96), .A3(new_n604), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n616), .A2(new_n620), .A3(new_n617), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n608), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT97), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n623), .A2(KEYINPUT97), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n624), .B(new_n625), .C1(new_n496), .C2(new_n497), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n485), .A2(new_n493), .ZN(new_n627));
  INV_X1    g441(.A(new_n495), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n485), .A2(new_n493), .A3(new_n495), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(KEYINPUT97), .A3(new_n623), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n501), .A2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n498), .A2(new_n501), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n557), .A2(G475), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n549), .A2(new_n511), .A3(new_n550), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(new_n551), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n622), .A2(new_n509), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n308), .A2(new_n615), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT98), .Z(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  AND3_X1   g459(.A1(new_n619), .A2(new_n608), .A3(new_n621), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n558), .A2(new_n510), .A3(new_n503), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT99), .B1(new_n622), .B2(new_n648), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n308), .A3(new_n615), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n348), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n342), .B(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OAI22_X1  g472(.A1(new_n363), .A2(new_n364), .B1(new_n658), .B2(new_n355), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n614), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n308), .A2(new_n610), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  AOI22_X1  g478(.A1(new_n433), .A2(new_n441), .B1(new_n457), .B2(G472), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n506), .B1(new_n507), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n558), .A2(new_n503), .A3(new_n668), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n622), .A2(new_n665), .A3(new_n660), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n308), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XOR2_X1   g486(.A(new_n667), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n308), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n607), .B(KEYINPUT38), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n407), .A2(new_n421), .B1(new_n429), .B2(new_n424), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n442), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n503), .A2(new_n639), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n659), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n608), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n675), .A2(new_n676), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT100), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  NOR3_X1   g501(.A1(new_n622), .A2(new_n665), .A3(new_n660), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n636), .A2(KEYINPUT101), .A3(new_n639), .A4(new_n668), .ZN(new_n689));
  INV_X1    g503(.A(new_n633), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n626), .B2(new_n631), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n498), .A2(new_n501), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n639), .B(new_n668), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n308), .A2(new_n688), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  OAI21_X1  g512(.A(new_n188), .B1(new_n282), .B2(new_n298), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G469), .ZN(new_n700));
  AND4_X1   g514(.A1(new_n459), .A2(new_n307), .A3(new_n299), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n641), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND2_X1  g518(.A1(new_n652), .A2(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT102), .B(G116), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G18));
  NOR4_X1   g521(.A1(new_n622), .A2(new_n665), .A3(new_n559), .A4(new_n660), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n700), .A2(new_n307), .A3(new_n299), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n365), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g528(.A(KEYINPUT103), .B(new_n357), .C1(new_n363), .C2(new_n364), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n429), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n451), .A2(new_n452), .B1(new_n435), .B2(KEYINPUT72), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n717), .B1(new_n718), .B2(new_n449), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n437), .A2(new_n438), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n431), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AND4_X1   g535(.A1(new_n510), .A2(new_n716), .A3(new_n721), .A4(new_n613), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n307), .A3(new_n299), .A4(new_n700), .ZN(new_n723));
  INV_X1    g537(.A(new_n681), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n646), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n712), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n622), .A2(new_n681), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n709), .A2(KEYINPUT104), .A3(new_n727), .A4(new_n722), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  AND3_X1   g544(.A1(new_n721), .A2(new_n613), .A3(new_n659), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n731), .A2(new_n689), .A3(new_n695), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n709), .A2(new_n732), .A3(new_n646), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  OAI21_X1  g548(.A(KEYINPUT105), .B1(new_n302), .B2(new_n264), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n736), .B(new_n293), .C1(new_n278), .C2(new_n296), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n735), .A2(G469), .A3(new_n301), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n299), .A2(new_n300), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n299), .A2(KEYINPUT106), .A3(new_n300), .A4(new_n738), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n665), .ZN(new_n744));
  AND4_X1   g558(.A1(new_n744), .A2(new_n689), .A3(new_n695), .A4(new_n716), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n605), .A2(new_n609), .A3(new_n606), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n743), .A2(new_n745), .A3(new_n307), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n696), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n746), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n751), .A2(new_n665), .A3(new_n365), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n750), .A2(new_n307), .A3(new_n743), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT107), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n748), .A2(new_n756), .A3(new_n753), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  INV_X1    g573(.A(new_n669), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n743), .A2(new_n307), .A3(new_n752), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND2_X1  g576(.A1(new_n636), .A2(new_n558), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT43), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n636), .A2(new_n765), .A3(new_n558), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n764), .A2(new_n614), .A3(new_n659), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n751), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n768), .B2(new_n767), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n187), .B1(new_n303), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n735), .A2(KEYINPUT45), .A3(new_n301), .A4(new_n737), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n300), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n299), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n307), .B(new_n673), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n770), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(KEYINPUT108), .B(G137), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n781), .B(new_n782), .ZN(G39));
  NAND4_X1  g597(.A1(new_n696), .A2(new_n665), .A3(new_n365), .A4(new_n746), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n307), .B1(new_n778), .B2(new_n779), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(KEYINPUT47), .B(new_n307), .C1(new_n778), .C2(new_n779), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n320), .ZN(G42));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n697), .A2(new_n671), .A3(new_n733), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n680), .A2(new_n668), .A3(new_n682), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n622), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n743), .A2(new_n794), .A3(new_n307), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n791), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n743), .A2(new_n794), .A3(new_n307), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n308), .B(new_n688), .C1(new_n760), .C2(new_n696), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT52), .A4(new_n733), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(KEYINPUT111), .A3(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(KEYINPUT111), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n701), .A2(new_n641), .B1(new_n708), .B2(new_n709), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n729), .A2(new_n804), .A3(new_n611), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n743), .A2(new_n307), .A3(new_n732), .A4(new_n746), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n503), .A2(new_n639), .A3(new_n667), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n746), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT110), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n665), .A2(new_n660), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(KEYINPUT110), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n308), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n761), .A2(new_n806), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n558), .B1(new_n635), .B2(new_n634), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT109), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT109), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n640), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n558), .A2(new_n503), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n608), .B(new_n510), .C1(new_n605), .C2(new_n606), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n308), .A2(new_n615), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n705), .A2(new_n662), .A3(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n805), .A2(new_n813), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n802), .A2(new_n803), .A3(new_n758), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n796), .A2(new_n799), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n824), .A2(new_n755), .A3(new_n826), .A4(new_n757), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n803), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n754), .A2(new_n803), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n824), .A2(new_n800), .A3(new_n832), .A4(new_n801), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n764), .A2(new_n506), .A3(new_n766), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n716), .A2(new_n613), .A3(new_n721), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n835), .A2(new_n836), .A3(new_n751), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT112), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n787), .A2(new_n788), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n700), .A2(new_n299), .ZN(new_n840));
  INV_X1    g654(.A(new_n307), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n838), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT50), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n709), .A2(new_n677), .A3(new_n609), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n835), .A2(new_n836), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n845), .B2(new_n846), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n844), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n845), .A2(new_n846), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT50), .A3(new_n849), .A4(new_n847), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n709), .A2(new_n746), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n357), .B(new_n506), .C1(new_n363), .C2(new_n364), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n855), .A2(new_n680), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n636), .A2(new_n639), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n855), .A2(new_n835), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n731), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n843), .A2(new_n854), .A3(KEYINPUT51), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n744), .A2(new_n716), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT48), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT114), .B1(new_n860), .B2(new_n866), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT48), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n709), .A2(new_n646), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n505), .B(G953), .C1(new_n874), .C2(new_n849), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n857), .A2(new_n814), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n864), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n862), .B1(new_n851), .B2(new_n853), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT51), .B1(new_n880), .B2(new_n843), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n829), .A2(new_n834), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n505), .A2(new_n260), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT49), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n840), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n840), .A2(new_n886), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n716), .A2(new_n307), .A3(new_n608), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n680), .A2(new_n889), .A3(new_n763), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n887), .A2(new_n677), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT115), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n885), .A2(new_n894), .A3(new_n891), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(G75));
  NOR2_X1   g710(.A1(new_n260), .A2(G952), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT118), .Z(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n597), .A2(new_n601), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT116), .Z(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT117), .Z(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(G210), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n904), .B(new_n188), .C1(new_n830), .C2(new_n833), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n599), .B(KEYINPUT55), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n905), .A2(KEYINPUT56), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n830), .A2(new_n833), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(G210), .A3(G902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n903), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n907), .B1(new_n905), .B2(KEYINPUT56), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n911), .A3(new_n906), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n915), .A3(new_n902), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n899), .B1(new_n913), .B2(new_n916), .ZN(G51));
  XOR2_X1   g731(.A(new_n300), .B(KEYINPUT57), .Z(new_n918));
  AND3_X1   g732(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n831), .B1(new_n830), .B2(new_n833), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n282), .A2(new_n298), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT119), .B(new_n918), .C1(new_n919), .C2(new_n920), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n909), .A2(G902), .A3(new_n773), .A4(new_n772), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n897), .B1(new_n926), .B2(new_n927), .ZN(G54));
  INV_X1    g742(.A(new_n897), .ZN(new_n929));
  AND4_X1   g743(.A1(KEYINPUT58), .A2(new_n909), .A3(G475), .A4(G902), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n549), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n549), .B2(new_n930), .ZN(G60));
  XOR2_X1   g746(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n933));
  NOR2_X1   g747(.A1(new_n501), .A2(new_n188), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n632), .B(new_n935), .C1(new_n919), .C2(new_n920), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n898), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n829), .A2(new_n834), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n632), .B1(new_n938), .B2(new_n935), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(G63));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n830), .A2(new_n833), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n943));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n898), .B1(new_n946), .B2(new_n350), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n942), .A2(new_n658), .A3(new_n945), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT122), .B1(new_n946), .B2(new_n350), .ZN(new_n950));
  INV_X1    g764(.A(new_n948), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  INV_X1    g766(.A(new_n350), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n952), .B(new_n953), .C1(new_n942), .C2(new_n945), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n899), .A2(new_n941), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n950), .A2(new_n951), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n949), .A2(new_n956), .ZN(G66));
  OAI21_X1  g771(.A(G953), .B1(new_n508), .B2(new_n585), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n805), .A2(new_n823), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT123), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n958), .B1(new_n961), .B2(G953), .ZN(new_n962));
  INV_X1    g776(.A(new_n901), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(G898), .B2(new_n260), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  NOR2_X1   g779(.A1(new_n539), .A2(new_n542), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT124), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n420), .B(new_n967), .Z(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n789), .A2(new_n781), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n819), .A2(new_n752), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n674), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n792), .B(KEYINPUT125), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n686), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n686), .A2(new_n973), .A3(KEYINPUT62), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n969), .B1(new_n978), .B2(G953), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n780), .A2(new_n725), .A3(new_n865), .ZN(new_n980));
  INV_X1    g794(.A(new_n761), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n758), .A2(new_n970), .A3(new_n973), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n260), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(G900), .B2(new_n260), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n968), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n979), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(G227), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n988), .B2(new_n666), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT126), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n990), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n979), .A2(new_n986), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n960), .B2(new_n983), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(new_n444), .A3(new_n421), .ZN(new_n998));
  INV_X1    g812(.A(new_n996), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n445), .B2(new_n408), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n825), .A2(new_n828), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n998), .A2(new_n929), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n421), .A2(new_n444), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n978), .A2(new_n961), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1003), .B(new_n1004), .C1(new_n1005), .C2(new_n999), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n999), .B1(new_n978), .B2(new_n961), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1004), .ZN(new_n1008));
  OAI21_X1  g822(.A(KEYINPUT127), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1002), .B1(new_n1006), .B2(new_n1009), .ZN(G57));
endmodule


