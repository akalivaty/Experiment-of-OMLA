//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n614, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT68), .Z(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT69), .Z(G261));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n452), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT70), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n463), .A3(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(new_n466), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT71), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(G101), .A3(G2104), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT72), .Z(new_n478));
  AND3_X1   g053(.A1(new_n470), .A2(new_n476), .A3(new_n478), .ZN(G160));
  NAND4_X1  g054(.A1(new_n475), .A2(new_n472), .A3(G2105), .A4(new_n466), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n484), .B1(new_n486), .B2(G136), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AND4_X1   g065(.A1(G2105), .A2(new_n475), .A3(new_n472), .A4(new_n466), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G126), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n475), .A2(new_n472), .A3(new_n466), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(G138), .A3(new_n474), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n464), .A2(new_n466), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n492), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(KEYINPUT4), .A2(new_n495), .B1(new_n500), .B2(new_n501), .ZN(new_n506));
  INV_X1    g081(.A(new_n488), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n507), .B1(G114), .B2(new_n474), .ZN(new_n508));
  INV_X1    g083(.A(G126), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n480), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT74), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  NAND2_X1  g088(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n521), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n523), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n522), .A2(G543), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n535), .A2(G51), .B1(new_n518), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g112(.A(KEYINPUT76), .B(new_n530), .C1(new_n523), .C2(new_n531), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT77), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n534), .A2(new_n537), .A3(new_n541), .A4(new_n538), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(G168));
  AOI22_X1  g118(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n520), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n523), .A2(new_n546), .B1(new_n525), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n520), .ZN(new_n551));
  INV_X1    g126(.A(new_n523), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G81), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT78), .B(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n535), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  AOI22_X1  g137(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n520), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n563), .A2(KEYINPUT79), .A3(new_n520), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n525), .A2(KEYINPUT9), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n525), .B2(new_n569), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n570), .A2(new_n571), .B1(new_n552), .B2(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  NAND2_X1  g151(.A1(new_n552), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n535), .A2(G49), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n520), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n523), .A2(new_n583), .B1(new_n525), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  AND2_X1   g162(.A1(new_n518), .A2(G60), .ZN(new_n588));
  AND2_X1   g163(.A1(G72), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(KEYINPUT80), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n552), .A2(G85), .B1(new_n535), .B2(G47), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n596), .A2(new_n520), .B1(new_n525), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n552), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n523), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n595), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n595), .B1(new_n609), .B2(G868), .ZN(G321));
  MUX2_X1   g186(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g187(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n609), .B1(new_n614), .B2(G860), .ZN(G148));
  OAI21_X1  g190(.A(G868), .B1(new_n608), .B2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g193(.A1(new_n465), .A2(G2105), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n501), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n480), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n486), .B2(G135), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(G2096), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n624), .A2(new_n631), .A3(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT83), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n635), .B2(new_n636), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n653), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n656), .B2(new_n652), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT86), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n670), .A2(new_n672), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n668), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n673), .A3(new_n668), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n674), .B1(new_n673), .B2(new_n668), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1981), .B(G1986), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G34), .ZN(new_n688));
  AOI21_X1  g263(.A(G29), .B1(new_n688), .B2(KEYINPUT24), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(KEYINPUT24), .B2(new_n688), .ZN(new_n690));
  INV_X1    g265(.A(G160), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(G2084), .Z(new_n694));
  AOI22_X1  g269(.A1(new_n501), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(new_n474), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT95), .Z(new_n697));
  NAND3_X1  g272(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT25), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n486), .B2(G139), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(new_n692), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n692), .B2(G33), .ZN(new_n703));
  INV_X1    g278(.A(G2072), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n694), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(G28), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n692), .B1(new_n706), .B2(G28), .ZN(new_n708));
  AND2_X1   g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  NOR2_X1   g284(.A1(KEYINPUT31), .A2(G11), .ZN(new_n710));
  OAI22_X1  g285(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n629), .B2(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(G16), .A2(G19), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n557), .B2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n712), .B1(new_n714), .B2(G1341), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(G1341), .ZN(new_n716));
  INV_X1    g291(.A(G1961), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NOR2_X1   g293(.A1(G171), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G5), .B2(new_n718), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n717), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT101), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n692), .A2(G26), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  AND2_X1   g300(.A1(new_n486), .A2(G140), .ZN(new_n726));
  INV_X1    g301(.A(G104), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n727), .A2(new_n474), .A3(KEYINPUT94), .ZN(new_n728));
  AOI21_X1  g303(.A(KEYINPUT94), .B1(new_n727), .B2(new_n474), .ZN(new_n729));
  OAI221_X1 g304(.A(G2104), .B1(G116), .B2(new_n474), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G128), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n480), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n725), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2067), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n705), .A2(new_n721), .A3(new_n723), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n703), .A2(new_n704), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT96), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n491), .A2(G129), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G105), .B2(new_n619), .ZN(new_n745));
  INV_X1    g320(.A(G141), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n740), .B(new_n745), .C1(new_n485), .C2(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT97), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(KEYINPUT97), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(new_n692), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n692), .B2(G32), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n737), .B(new_n739), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n755));
  NAND2_X1  g330(.A1(G168), .A2(G16), .ZN(new_n756));
  MUX2_X1   g331(.A(KEYINPUT98), .B(new_n755), .S(new_n756), .Z(new_n757));
  XOR2_X1   g332(.A(KEYINPUT99), .B(G1966), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT100), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n692), .A2(G35), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n692), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n752), .A2(new_n753), .B1(G2090), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G27), .A2(G29), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G164), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2078), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n757), .A2(new_n758), .ZN(new_n769));
  NOR2_X1   g344(.A1(G4), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n609), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT93), .B(G1348), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n771), .A2(new_n772), .B1(new_n763), .B2(G2090), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n718), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT23), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  AND4_X1   g353(.A1(new_n769), .A2(new_n773), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n754), .A2(new_n760), .A3(new_n768), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G6), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n586), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT89), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT32), .B(G1981), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n718), .A2(G23), .ZN(new_n786));
  INV_X1    g361(.A(G288), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n718), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n718), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n718), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1971), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n790), .B2(new_n791), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n785), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n785), .A2(new_n792), .A3(KEYINPUT91), .A4(new_n796), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n799), .A2(KEYINPUT34), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT92), .ZN(new_n802));
  AOI21_X1  g377(.A(KEYINPUT34), .B1(new_n799), .B2(new_n800), .ZN(new_n803));
  NAND2_X1  g378(.A1(G290), .A2(G16), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n718), .A2(G24), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G1986), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n692), .A2(G25), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n486), .A2(G131), .ZN(new_n810));
  INV_X1    g385(.A(G119), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n474), .A2(G107), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n480), .A2(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n809), .B1(new_n815), .B2(new_n692), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT35), .B(G1991), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n806), .A2(new_n807), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n803), .A2(new_n808), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n802), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n802), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n780), .B1(new_n822), .B2(new_n824), .ZN(G311));
  INV_X1    g400(.A(new_n780), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(G150));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n535), .A2(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n523), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n518), .A2(G67), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n520), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n829), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n835), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n552), .A2(G93), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT102), .A4(new_n830), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(new_n556), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT103), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n553), .A2(new_n555), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(new_n551), .C1(new_n835), .C2(new_n832), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n841), .B1(new_n840), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n614), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  AOI21_X1  g425(.A(G860), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n836), .A2(new_n839), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(G145));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n492), .A2(new_n503), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT104), .B1(new_n506), .B2(new_n510), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n748), .A2(new_n749), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n733), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n733), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n750), .A2(new_n734), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n861), .A3(new_n864), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT105), .B1(new_n701), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(KEYINPUT105), .B2(new_n701), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n874), .A2(new_n867), .A3(new_n869), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n491), .A2(G130), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n474), .A2(G118), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(G142), .B2(new_n486), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n621), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n815), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n873), .A2(new_n875), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G162), .B(new_n629), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n691), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n887), .A2(KEYINPUT107), .A3(new_n889), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT107), .B1(new_n887), .B2(new_n889), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n857), .B(new_n890), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g469(.A(G290), .B(new_n787), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n586), .B(G166), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n897), .B2(new_n898), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT42), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n609), .A2(new_n614), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n846), .B(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G299), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT108), .B1(new_n906), .B2(new_n608), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n609), .A2(G299), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n609), .A2(G299), .A3(KEYINPUT108), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(KEYINPUT41), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n906), .A2(new_n608), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n908), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n905), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n903), .A2(new_n913), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n903), .B1(new_n913), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(G868), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n853), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(G868), .B2(new_n923), .ZN(G295));
  OAI21_X1  g499(.A(new_n922), .B1(G868), .B2(new_n923), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  INV_X1    g502(.A(new_n902), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n540), .A2(new_n929), .A3(new_n542), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n844), .B2(new_n845), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n840), .A2(new_n843), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT103), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n930), .ZN(new_n936));
  AOI21_X1  g511(.A(G301), .B1(G168), .B2(KEYINPUT110), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n937), .B1(new_n932), .B2(new_n936), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n911), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(new_n936), .ZN(new_n942));
  INV_X1    g517(.A(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n944), .A2(new_n938), .B1(new_n914), .B2(new_n917), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n928), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n946), .A2(new_n857), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n941), .A2(new_n945), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n902), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n927), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n908), .A2(new_n915), .ZN(new_n951));
  OAI211_X1 g526(.A(KEYINPUT41), .B(new_n951), .C1(new_n939), .C2(new_n940), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n916), .B1(new_n944), .B2(new_n938), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n952), .B(new_n902), .C1(new_n953), .C2(new_n911), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n954), .A2(new_n946), .A3(new_n857), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n926), .B1(new_n950), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(KEYINPUT111), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n954), .A2(new_n946), .A3(new_n960), .A4(new_n857), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT43), .A4(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n949), .A2(new_n946), .A3(new_n927), .A4(new_n857), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n927), .B1(new_n955), .B2(KEYINPUT111), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n959), .B1(new_n966), .B2(new_n961), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n957), .B1(new_n965), .B2(new_n967), .ZN(G397));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT45), .B1(new_n861), .B2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n470), .A2(new_n476), .A3(new_n478), .A4(G40), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n733), .B(G2067), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n750), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n976), .B2(new_n750), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n815), .B(new_n817), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT113), .B1(G290), .B2(G1986), .ZN(new_n981));
  NAND2_X1  g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n981), .B(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n980), .B1(new_n973), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT114), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n969), .B1(new_n506), .B2(new_n510), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n971), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(G1384), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n505), .B2(new_n511), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI211_X1 g569(.A(KEYINPUT116), .B(new_n991), .C1(new_n505), .C2(new_n511), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n758), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT117), .B(new_n758), .C1(new_n994), .C2(new_n995), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n492), .B2(new_n503), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n971), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT118), .B(G2084), .Z(new_n1003));
  AOI21_X1  g578(.A(G1384), .B1(new_n505), .B2(new_n511), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1002), .B(new_n1003), .C1(new_n1004), .C2(new_n1001), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n998), .A2(new_n999), .A3(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n986), .B(G8), .C1(new_n1006), .C2(G286), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT122), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G168), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1005), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n996), .B2(new_n997), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n1008), .B(new_n1011), .C1(new_n1013), .C2(new_n999), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT122), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1007), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1009), .B1(new_n1013), .B2(new_n999), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1017), .A2(new_n986), .A3(new_n1010), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT123), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT62), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1008), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1006), .A2(KEYINPUT122), .A3(new_n1010), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1017), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(KEYINPUT51), .A3(new_n1011), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT123), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .A4(new_n1007), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1019), .A2(new_n1020), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1020), .B1(new_n1019), .B2(new_n1028), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n859), .A2(new_n860), .A3(new_n990), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1031), .B(new_n972), .C1(new_n1004), .C2(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g607(.A(G1971), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n512), .A2(new_n969), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n1002), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1009), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G166), .A2(new_n1009), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT55), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1004), .A2(new_n1001), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n971), .B1(new_n987), .B2(KEYINPUT50), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1037), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1034), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1041), .B1(new_n1047), .B2(G8), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  OAI221_X1 g624(.A(G8), .B1(G288), .B2(new_n1049), .C1(new_n971), .C2(new_n987), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT52), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G305), .A2(G1981), .ZN(new_n1052));
  INV_X1    g627(.A(G1981), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n586), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n987), .A2(new_n971), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(new_n1009), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1052), .A2(KEYINPUT49), .A3(new_n1054), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(new_n787), .B2(G1976), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1050), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(KEYINPUT115), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1050), .A2(new_n1066), .A3(new_n1063), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1051), .B(new_n1061), .C1(new_n1065), .C2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1043), .A2(new_n1048), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1032), .B2(G2078), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT124), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n1070), .C1(new_n1032), .C2(G2078), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1036), .A2(new_n1002), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1072), .A2(new_n1074), .B1(new_n717), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n994), .A2(new_n995), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1070), .A2(G2078), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1069), .A2(G171), .A3(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1029), .A2(new_n1030), .A3(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(G171), .B(KEYINPUT54), .Z(new_n1083));
  AND3_X1   g658(.A1(new_n1076), .A2(new_n1079), .A3(new_n1083), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1070), .B(G2078), .C1(new_n971), .C2(KEYINPUT125), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1031), .C1(KEYINPUT125), .C2(new_n971), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1086), .A2(new_n970), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1083), .B1(new_n1076), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1069), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n568), .B2(new_n572), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n572), .B(new_n1090), .C1(new_n566), .C2(new_n567), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT56), .B(G2072), .Z(new_n1096));
  NOR2_X1   g671(.A1(new_n1032), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1956), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1098), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1100), .B(new_n1094), .C1(new_n1032), .C2(new_n1096), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1099), .A2(new_n1101), .A3(KEYINPUT61), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT61), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1348), .ZN(new_n1105));
  INV_X1    g680(.A(G2067), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1075), .A2(new_n1105), .B1(new_n1106), .B2(new_n1058), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n609), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1107), .A2(new_n609), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1108), .B1(new_n1107), .B2(new_n609), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1032), .A2(G1996), .B1(new_n1058), .B2(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1115), .A2(KEYINPUT121), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(KEYINPUT121), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1113), .B1(new_n1118), .B2(new_n557), .ZN(new_n1119));
  AOI211_X1 g694(.A(KEYINPUT59), .B(new_n556), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1104), .B(new_n1112), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1099), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1107), .A2(new_n608), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1101), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1089), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1019), .A2(new_n1028), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1061), .A2(new_n1049), .A3(new_n787), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1054), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1059), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1042), .B2(new_n1068), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1069), .A2(G168), .A3(new_n1017), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT63), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1043), .A2(new_n1135), .A3(new_n1068), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(G168), .A3(new_n1017), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1131), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1127), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n985), .B1(new_n1082), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n973), .A2(new_n976), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT46), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n975), .A2(new_n750), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1142), .B1(new_n974), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT47), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1148), .A2(KEYINPUT126), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(KEYINPUT126), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n810), .A2(new_n817), .A3(new_n814), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n978), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n733), .A2(new_n1106), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n974), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n974), .A2(G1986), .A3(G290), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT48), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(KEYINPUT127), .B2(new_n980), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1154), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1149), .A2(new_n1150), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1140), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g736(.A(G319), .ZN(new_n1163));
  NOR3_X1   g737(.A1(G229), .A2(new_n1163), .A3(G227), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n893), .A2(new_n650), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g739(.A1(new_n950), .A2(new_n956), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n1165), .A2(new_n1166), .ZN(G308));
  OR2_X1    g741(.A1(new_n1165), .A2(new_n1166), .ZN(G225));
endmodule


