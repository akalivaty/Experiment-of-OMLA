

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U325 ( .A(n578), .B(n577), .ZN(n579) );
  NOR2_X1 U326 ( .A1(n457), .A2(n542), .ZN(n569) );
  NOR2_X1 U327 ( .A1(n572), .A2(n571), .ZN(n580) );
  XNOR2_X1 U328 ( .A(n379), .B(n378), .ZN(n539) );
  NOR2_X1 U329 ( .A1(n377), .A2(n376), .ZN(n379) );
  XNOR2_X1 U330 ( .A(n369), .B(n368), .ZN(n377) );
  NOR2_X1 U331 ( .A1(n294), .A2(n293), .ZN(n369) );
  XNOR2_X1 U332 ( .A(n349), .B(n295), .ZN(n294) );
  INV_X1 U333 ( .A(n348), .ZN(n295) );
  XNOR2_X1 U334 ( .A(n370), .B(KEYINPUT41), .ZN(n460) );
  XNOR2_X1 U335 ( .A(n329), .B(n436), .ZN(n370) );
  XNOR2_X1 U336 ( .A(n320), .B(n296), .ZN(n298) );
  XNOR2_X1 U337 ( .A(n319), .B(n297), .ZN(n296) );
  INV_X1 U338 ( .A(KEYINPUT74), .ZN(n297) );
  XNOR2_X1 U339 ( .A(G176GAT), .B(G92GAT), .ZN(n318) );
  INV_X1 U340 ( .A(n366), .ZN(n293) );
  XNOR2_X1 U341 ( .A(G134GAT), .B(G92GAT), .ZN(n310) );
  INV_X1 U342 ( .A(KEYINPUT45), .ZN(n371) );
  NOR2_X1 U343 ( .A1(n581), .A2(n566), .ZN(n366) );
  INV_X1 U344 ( .A(KEYINPUT76), .ZN(n303) );
  XOR2_X1 U345 ( .A(n324), .B(KEYINPUT32), .Z(n299) );
  XNOR2_X1 U346 ( .A(n371), .B(KEYINPUT114), .ZN(n372) );
  XNOR2_X1 U347 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n318), .B(G64GAT), .ZN(n385) );
  XNOR2_X1 U350 ( .A(n322), .B(n305), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U352 ( .A(n313), .B(n312), .ZN(n317) );
  XNOR2_X1 U353 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n458) );
  XNOR2_X1 U354 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U355 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XOR2_X1 U356 ( .A(KEYINPUT10), .B(n428), .Z(n301) );
  XOR2_X1 U357 ( .A(G36GAT), .B(G190GAT), .Z(n390) );
  XNOR2_X1 U358 ( .A(n390), .B(G218GAT), .ZN(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n307) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G85GAT), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n302), .B(KEYINPUT73), .ZN(n322) );
  NAND2_X1 U362 ( .A1(G232GAT), .A2(G233GAT), .ZN(n304) );
  XOR2_X1 U363 ( .A(n307), .B(n306), .Z(n313) );
  XOR2_X1 U364 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n309) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U367 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n315) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(G29GAT), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U370 ( .A(KEYINPUT7), .B(n316), .ZN(n345) );
  XNOR2_X1 U371 ( .A(n317), .B(n345), .ZN(n566) );
  XOR2_X1 U372 ( .A(G57GAT), .B(KEYINPUT13), .Z(n352) );
  XOR2_X1 U373 ( .A(n385), .B(n352), .Z(n320) );
  NAND2_X1 U374 ( .A1(G230GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n322), .B(KEYINPUT31), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n298), .B(n323), .ZN(n324) );
  XOR2_X1 U377 ( .A(G120GAT), .B(G71GAT), .Z(n448) );
  XNOR2_X1 U378 ( .A(n448), .B(KEYINPUT33), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n299), .B(n325), .ZN(n329) );
  XOR2_X1 U380 ( .A(G78GAT), .B(KEYINPUT72), .Z(n327) );
  XNOR2_X1 U381 ( .A(G148GAT), .B(G106GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U383 ( .A(G204GAT), .B(n328), .ZN(n436) );
  XOR2_X1 U384 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n331) );
  XNOR2_X1 U385 ( .A(KEYINPUT68), .B(KEYINPUT71), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n344) );
  XOR2_X1 U387 ( .A(G197GAT), .B(G36GAT), .Z(n333) );
  XNOR2_X1 U388 ( .A(G169GAT), .B(G50GAT), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U390 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n335) );
  XNOR2_X1 U391 ( .A(G8GAT), .B(KEYINPUT67), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U393 ( .A(n337), .B(n336), .Z(n342) );
  XOR2_X1 U394 ( .A(G113GAT), .B(G1GAT), .Z(n412) );
  XOR2_X1 U395 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U396 ( .A(n431), .B(G15GAT), .Z(n339) );
  NAND2_X1 U397 ( .A1(G229GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n412), .B(n340), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n346) );
  XOR2_X1 U402 ( .A(n346), .B(n345), .Z(n509) );
  INV_X1 U403 ( .A(n509), .ZN(n573) );
  NAND2_X1 U404 ( .A1(n460), .A2(n573), .ZN(n349) );
  XOR2_X1 U405 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n347) );
  XNOR2_X1 U406 ( .A(KEYINPUT111), .B(n347), .ZN(n348) );
  XOR2_X1 U407 ( .A(KEYINPUT14), .B(G78GAT), .Z(n351) );
  XNOR2_X1 U408 ( .A(G22GAT), .B(G71GAT), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U410 ( .A(n353), .B(n352), .Z(n356) );
  XOR2_X1 U411 ( .A(G15GAT), .B(G127GAT), .Z(n439) );
  XNOR2_X1 U412 ( .A(G8GAT), .B(G183GAT), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n354), .B(KEYINPUT77), .ZN(n384) );
  XNOR2_X1 U414 ( .A(n439), .B(n384), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n358) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U419 ( .A(n360), .B(n359), .Z(n365) );
  XOR2_X1 U420 ( .A(G211GAT), .B(G64GAT), .Z(n362) );
  XNOR2_X1 U421 ( .A(G1GAT), .B(G155GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n363), .B(KEYINPUT12), .ZN(n364) );
  XOR2_X1 U424 ( .A(n365), .B(n364), .Z(n581) );
  INV_X1 U425 ( .A(n581), .ZN(n492) );
  XNOR2_X1 U426 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n368) );
  NAND2_X1 U427 ( .A1(n509), .A2(n370), .ZN(n375) );
  XOR2_X1 U428 ( .A(n566), .B(KEYINPUT36), .Z(n586) );
  NOR2_X1 U429 ( .A1(n492), .A2(n586), .ZN(n373) );
  NOR2_X1 U430 ( .A1(n375), .A2(n374), .ZN(n376) );
  XNOR2_X1 U431 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n378) );
  XNOR2_X1 U432 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n380) );
  XNOR2_X1 U433 ( .A(n380), .B(KEYINPUT17), .ZN(n381) );
  XOR2_X1 U434 ( .A(n381), .B(KEYINPUT19), .Z(n383) );
  XNOR2_X1 U435 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n383), .B(n382), .ZN(n456) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n394) );
  XOR2_X1 U438 ( .A(G211GAT), .B(KEYINPUT21), .Z(n387) );
  XNOR2_X1 U439 ( .A(G197GAT), .B(G218GAT), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n430) );
  XNOR2_X1 U441 ( .A(n430), .B(KEYINPUT92), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n388), .B(G204GAT), .ZN(n389) );
  XOR2_X1 U443 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U444 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U447 ( .A(n456), .B(n395), .Z(n515) );
  INV_X1 U448 ( .A(n515), .ZN(n529) );
  NAND2_X1 U449 ( .A1(n539), .A2(n529), .ZN(n397) );
  XOR2_X1 U450 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n421) );
  XOR2_X1 U452 ( .A(KEYINPUT80), .B(KEYINPUT0), .Z(n399) );
  XNOR2_X1 U453 ( .A(G134GAT), .B(KEYINPUT79), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n447) );
  XNOR2_X1 U455 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n400), .B(KEYINPUT3), .ZN(n425) );
  XNOR2_X1 U457 ( .A(n447), .B(n425), .ZN(n420) );
  XOR2_X1 U458 ( .A(G148GAT), .B(KEYINPUT89), .Z(n402) );
  XNOR2_X1 U459 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U461 ( .A(G57GAT), .B(G127GAT), .Z(n404) );
  XNOR2_X1 U462 ( .A(G141GAT), .B(G120GAT), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U464 ( .A(n406), .B(n405), .Z(n418) );
  XOR2_X1 U465 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n408) );
  XNOR2_X1 U466 ( .A(KEYINPUT88), .B(KEYINPUT6), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n416) );
  XOR2_X1 U468 ( .A(KEYINPUT4), .B(G162GAT), .Z(n410) );
  XNOR2_X1 U469 ( .A(G29GAT), .B(G85GAT), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U471 ( .A(n412), .B(n411), .Z(n414) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U476 ( .A(n420), .B(n419), .Z(n527) );
  INV_X1 U477 ( .A(n527), .ZN(n558) );
  NAND2_X1 U478 ( .A1(n421), .A2(n558), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n422), .B(KEYINPUT64), .ZN(n572) );
  XOR2_X1 U480 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n424) );
  XNOR2_X1 U481 ( .A(KEYINPUT87), .B(KEYINPUT23), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n435) );
  XOR2_X1 U483 ( .A(n425), .B(KEYINPUT24), .Z(n427) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U486 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n472) );
  NOR2_X1 U491 ( .A1(n572), .A2(n472), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n438), .B(KEYINPUT55), .ZN(n457) );
  XNOR2_X1 U493 ( .A(n439), .B(G99GAT), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n440), .B(G190GAT), .ZN(n444) );
  XOR2_X1 U495 ( .A(G183GAT), .B(G176GAT), .Z(n442) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G113GAT), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U498 ( .A(n444), .B(n443), .Z(n454) );
  XOR2_X1 U499 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n446) );
  XNOR2_X1 U500 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n452) );
  XOR2_X1 U502 ( .A(n448), .B(n447), .Z(n450) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U507 ( .A(n456), .B(n455), .Z(n531) );
  INV_X1 U508 ( .A(n531), .ZN(n542) );
  NAND2_X1 U509 ( .A1(n566), .A2(n569), .ZN(n459) );
  NAND2_X1 U510 ( .A1(n569), .A2(n460), .ZN(n464) );
  XOR2_X1 U511 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n462) );
  XOR2_X1 U512 ( .A(G176GAT), .B(KEYINPUT56), .Z(n461) );
  XNOR2_X1 U513 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U514 ( .A(n464), .B(n463), .ZN(G1349GAT) );
  XOR2_X1 U515 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n482) );
  NAND2_X1 U516 ( .A1(n370), .A2(n573), .ZN(n495) );
  NOR2_X1 U517 ( .A1(n492), .A2(n566), .ZN(n465) );
  XNOR2_X1 U518 ( .A(n465), .B(KEYINPUT16), .ZN(n479) );
  NAND2_X1 U519 ( .A1(n472), .A2(n542), .ZN(n466) );
  XNOR2_X1 U520 ( .A(n466), .B(KEYINPUT26), .ZN(n571) );
  XNOR2_X1 U521 ( .A(KEYINPUT27), .B(n515), .ZN(n474) );
  NOR2_X1 U522 ( .A1(n571), .A2(n474), .ZN(n556) );
  NOR2_X1 U523 ( .A1(n515), .A2(n542), .ZN(n467) );
  NOR2_X1 U524 ( .A1(n472), .A2(n467), .ZN(n468) );
  XOR2_X1 U525 ( .A(KEYINPUT25), .B(n468), .Z(n469) );
  NOR2_X1 U526 ( .A1(n556), .A2(n469), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n470), .A2(n527), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT94), .B(n471), .Z(n478) );
  XNOR2_X1 U529 ( .A(KEYINPUT65), .B(KEYINPUT28), .ZN(n473) );
  XOR2_X1 U530 ( .A(n473), .B(n472), .Z(n534) );
  OR2_X1 U531 ( .A1(n474), .A2(n534), .ZN(n475) );
  NOR2_X1 U532 ( .A1(n558), .A2(n475), .ZN(n540) );
  NAND2_X1 U533 ( .A1(n540), .A2(n542), .ZN(n476) );
  XOR2_X1 U534 ( .A(KEYINPUT93), .B(n476), .Z(n477) );
  NAND2_X1 U535 ( .A1(n478), .A2(n477), .ZN(n491) );
  NAND2_X1 U536 ( .A1(n479), .A2(n491), .ZN(n510) );
  NOR2_X1 U537 ( .A1(n495), .A2(n510), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT95), .B(n480), .Z(n489) );
  NAND2_X1 U539 ( .A1(n489), .A2(n527), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U541 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  XOR2_X1 U542 ( .A(G8GAT), .B(KEYINPUT97), .Z(n485) );
  NAND2_X1 U543 ( .A1(n489), .A2(n529), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U546 ( .A1(n489), .A2(n531), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  NAND2_X1 U549 ( .A1(n489), .A2(n534), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U551 ( .A1(n492), .A2(n491), .ZN(n493) );
  NOR2_X1 U552 ( .A1(n586), .A2(n493), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n494), .ZN(n526) );
  NOR2_X1 U554 ( .A1(n526), .A2(n495), .ZN(n497) );
  XNOR2_X1 U555 ( .A(KEYINPUT38), .B(KEYINPUT99), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(n507) );
  NOR2_X1 U557 ( .A1(n507), .A2(n558), .ZN(n501) );
  XOR2_X1 U558 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n499) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT100), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n503) );
  NOR2_X1 U563 ( .A1(n515), .A2(n507), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(n504), .ZN(G1329GAT) );
  NOR2_X1 U566 ( .A1(n507), .A2(n542), .ZN(n505) );
  XOR2_X1 U567 ( .A(KEYINPUT40), .B(n505), .Z(n506) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  INV_X1 U569 ( .A(n534), .ZN(n521) );
  NOR2_X1 U570 ( .A1(n507), .A2(n521), .ZN(n508) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  NAND2_X1 U572 ( .A1(n509), .A2(n460), .ZN(n525) );
  NOR2_X1 U573 ( .A1(n525), .A2(n510), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(KEYINPUT105), .ZN(n520) );
  NOR2_X1 U575 ( .A1(n558), .A2(n520), .ZN(n513) );
  XNOR2_X1 U576 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n514), .Z(G1332GAT) );
  NOR2_X1 U579 ( .A1(n515), .A2(n520), .ZN(n516) );
  XOR2_X1 U580 ( .A(KEYINPUT106), .B(n516), .Z(n517) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(n517), .ZN(G1333GAT) );
  NOR2_X1 U582 ( .A1(n542), .A2(n520), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1334GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U586 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(n524), .ZN(G1335GAT) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n535), .A2(n527), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n535), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U594 ( .A(G99GAT), .B(KEYINPUT109), .Z(n533) );
  NAND2_X1 U595 ( .A1(n535), .A2(n531), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1338GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n537) );
  NAND2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U600 ( .A(G106GAT), .B(n538), .Z(G1339GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n544) );
  NAND2_X1 U602 ( .A1(n539), .A2(n540), .ZN(n541) );
  NOR2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n553) );
  NAND2_X1 U604 ( .A1(n553), .A2(n573), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U606 ( .A(G113GAT), .B(n545), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n547) );
  NAND2_X1 U608 ( .A1(n553), .A2(n460), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(n548), .ZN(G1341GAT) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(KEYINPUT120), .ZN(n552) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U613 ( .A1(n553), .A2(n581), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(n552), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U617 ( .A1(n553), .A2(n566), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U619 ( .A1(n539), .A2(n556), .ZN(n557) );
  NOR2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n573), .A2(n565), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n561) );
  NAND2_X1 U624 ( .A1(n565), .A2(n460), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT53), .Z(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n581), .A2(n565), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U631 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U632 ( .A1(n569), .A2(n573), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(n568), .ZN(G1348GAT) );
  NAND2_X1 U634 ( .A1(n581), .A2(n569), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  NAND2_X1 U637 ( .A1(n580), .A2(n573), .ZN(n574) );
  XNOR2_X1 U638 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n578) );
  INV_X1 U641 ( .A(n580), .ZN(n585) );
  OR2_X1 U642 ( .A1(n585), .A2(n370), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U645 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n584) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n588) );
  NOR2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U650 ( .A(n588), .B(n587), .Z(G1355GAT) );
endmodule

