//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1174, new_n1175;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR3_X1    g032(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n456), .B1(new_n453), .B2(new_n457), .ZN(new_n459));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  OAI211_X1 g035(.A(new_n458), .B(new_n459), .C1(new_n452), .C2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n470), .A2(new_n472), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(new_n464), .B2(new_n465), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n483), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n492), .B2(G114), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n478), .C2(new_n479), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n478), .B2(new_n479), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n500), .B(new_n503), .C1(new_n479), .C2(new_n478), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n498), .B1(new_n502), .B2(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n510), .A2(G651), .B1(new_n514), .B2(G50), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n507), .A2(new_n517), .A3(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n515), .B1(new_n516), .B2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n512), .A2(KEYINPUT71), .A3(new_n513), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n526), .A2(G543), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n520), .A2(G89), .A3(new_n521), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n507), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  XNOR2_X1  g112(.A(KEYINPUT72), .B(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n528), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n520), .A2(G90), .A3(new_n521), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(new_n528), .A2(G43), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n542), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n545), .B(new_n547), .C1(new_n548), .C2(new_n522), .ZN(new_n549));
  INV_X1    g124(.A(G860), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n549), .A2(new_n550), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT73), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND3_X1  g131(.A1(new_n526), .A2(G543), .A3(new_n527), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT74), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n511), .B1(new_n517), .B2(new_n525), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n560), .A2(new_n561), .A3(G53), .A4(new_n527), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(KEYINPUT9), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n520), .A2(G91), .A3(new_n521), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n508), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  OAI211_X1 g145(.A(KEYINPUT74), .B(new_n570), .C1(new_n557), .C2(new_n558), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(G299));
  NAND3_X1  g147(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(G301));
  OAI21_X1  g148(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n574));
  INV_X1    g149(.A(G49), .ZN(new_n575));
  INV_X1    g150(.A(G87), .ZN(new_n576));
  OAI221_X1 g151(.A(new_n574), .B1(new_n575), .B2(new_n557), .C1(new_n522), .C2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n507), .A2(G61), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n578), .A2(new_n579), .B1(G73), .B2(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n507), .A2(KEYINPUT75), .A3(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n542), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT76), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT77), .ZN(new_n585));
  INV_X1    g160(.A(new_n522), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n585), .B1(G86), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n586), .A2(G85), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n528), .A2(G47), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n542), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n528), .A2(G54), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n507), .A2(G66), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT79), .Z(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n522), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n520), .A2(G92), .A3(new_n521), .A4(new_n601), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n600), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n594), .B1(new_n606), .B2(G868), .ZN(G321));
  XNOR2_X1  g182(.A(G321), .B(KEYINPUT80), .ZN(G284));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n549), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n604), .A2(new_n605), .ZN(new_n617));
  INV_X1    g192(.A(new_n600), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n616), .B1(new_n620), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g197(.A1(new_n481), .A2(G135), .B1(G123), .B2(new_n484), .ZN(new_n623));
  OR3_X1    g198(.A1(new_n483), .A2(KEYINPUT82), .A3(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT82), .B1(new_n483), .B2(G111), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n624), .A2(G2104), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n623), .A2(KEYINPUT83), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n470), .A2(new_n474), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT13), .B(G2100), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n633), .A2(new_n634), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n675), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n679), .C1(new_n672), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G27), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT95), .Z(new_n690));
  INV_X1    g265(.A(new_n504), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n503), .B1(new_n470), .B2(new_n500), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n497), .B(new_n496), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n690), .B1(new_n693), .B2(G29), .ZN(new_n694));
  INV_X1    g269(.A(G2078), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G28), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT30), .ZN(new_n698));
  AOI21_X1  g273(.A(G29), .B1(new_n697), .B2(KEYINPUT30), .ZN(new_n699));
  OR2_X1    g274(.A1(KEYINPUT31), .A2(G11), .ZN(new_n700));
  NAND2_X1  g275(.A1(KEYINPUT31), .A2(G11), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n698), .A2(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT26), .Z(new_n705));
  INV_X1    g280(.A(G129), .ZN(new_n706));
  INV_X1    g281(.A(new_n484), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n703), .B(new_n705), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(new_n688), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n688), .B2(G32), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n702), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n696), .B(new_n713), .C1(new_n711), .C2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(G115), .A2(G2104), .ZN(new_n715));
  INV_X1    g290(.A(G127), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n480), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n483), .B1(new_n717), .B2(KEYINPUT93), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(KEYINPUT93), .B2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n720));
  NAND2_X1  g295(.A1(G103), .A2(G2104), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G2105), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n483), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n481), .A2(G139), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G33), .B(new_n725), .S(G29), .Z(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(G2072), .Z(new_n727));
  AND2_X1   g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n688), .B1(KEYINPUT24), .B2(G34), .ZN(new_n729));
  OAI22_X1  g304(.A1(G160), .A2(new_n688), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI22_X1  g305(.A1(new_n730), .A2(G2084), .B1(new_n694), .B2(new_n695), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n632), .A2(new_n688), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n731), .B(new_n732), .C1(G2084), .C2(new_n730), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n714), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(G19), .B(new_n549), .S(G16), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1341), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n484), .A2(G128), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n483), .A2(G116), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n739));
  INV_X1    g314(.A(G140), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n470), .A2(new_n483), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n737), .B1(new_n738), .B2(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT91), .Z(new_n744));
  XOR2_X1   g319(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n688), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2067), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n734), .A2(new_n736), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G20), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT97), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT23), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n610), .B2(new_n751), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1956), .Z(new_n756));
  INV_X1    g331(.A(G2090), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n688), .A2(G35), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT96), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n488), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT29), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n756), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT98), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G4), .A2(G16), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n606), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT90), .B(G1348), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G168), .A2(new_n751), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n751), .B2(G21), .ZN(new_n770));
  INV_X1    g345(.A(G1966), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT94), .Z(new_n773));
  AOI22_X1  g348(.A1(new_n770), .A2(new_n771), .B1(new_n757), .B2(new_n761), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n751), .A2(G5), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G171), .B2(new_n751), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AND4_X1   g353(.A1(new_n768), .A2(new_n773), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n762), .A2(new_n763), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n750), .A2(new_n764), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G6), .B(G305), .S(G16), .Z(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT32), .B(G1981), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT89), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n782), .A2(new_n784), .ZN(new_n786));
  MUX2_X1   g361(.A(G23), .B(G288), .S(G16), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT33), .B(G1976), .Z(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n751), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n751), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G1971), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n787), .A2(new_n788), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(G1971), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR4_X1   g370(.A1(new_n785), .A2(new_n786), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n751), .A2(G24), .ZN(new_n799));
  INV_X1    g374(.A(G290), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n751), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G1986), .Z(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT87), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n484), .A2(G119), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n483), .A2(G107), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(G131), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n804), .B1(new_n805), .B2(new_n806), .C1(new_n807), .C2(new_n741), .ZN(new_n808));
  MUX2_X1   g383(.A(G25), .B(new_n808), .S(G29), .Z(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT86), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n809), .B(new_n811), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n802), .A2(KEYINPUT87), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n798), .A2(new_n803), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n796), .A2(new_n797), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n814), .A2(KEYINPUT36), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT36), .B1(new_n814), .B2(new_n815), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n781), .B1(new_n817), .B2(new_n818), .ZN(G311));
  INV_X1    g394(.A(new_n781), .ZN(new_n820));
  INV_X1    g395(.A(new_n818), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n816), .ZN(G150));
  NOR2_X1   g397(.A1(new_n619), .A2(new_n613), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT38), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n528), .A2(G55), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(new_n542), .ZN(new_n827));
  INV_X1    g402(.A(G93), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n825), .B(new_n827), .C1(new_n828), .C2(new_n522), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n549), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n824), .B(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(new_n550), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n829), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n708), .B(new_n742), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n693), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n839), .A2(KEYINPUT100), .A3(new_n719), .A4(new_n724), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n725), .B(KEYINPUT100), .Z(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n484), .A2(G130), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n483), .A2(G118), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  INV_X1    g420(.A(G142), .ZN(new_n846));
  OAI221_X1 g421(.A(new_n843), .B1(new_n844), .B2(new_n845), .C1(new_n846), .C2(new_n741), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n808), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n637), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT101), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n842), .A2(new_n850), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n842), .A2(KEYINPUT102), .A3(new_n850), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT99), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G160), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n849), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n853), .C1(new_n842), .C2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n861), .A2(KEYINPUT40), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT40), .B1(new_n861), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(G395));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n610), .A2(new_n619), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n606), .A2(G299), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(KEYINPUT103), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n606), .A2(G299), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n870), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n871), .A2(new_n872), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n870), .ZN(new_n879));
  AOI211_X1 g454(.A(KEYINPUT104), .B(KEYINPUT41), .C1(new_n871), .C2(new_n872), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n549), .A2(new_n829), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n549), .A2(new_n829), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n620), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(KEYINPUT105), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n873), .A2(new_n875), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n886), .A2(KEYINPUT105), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(G166), .B(G288), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n583), .A2(new_n587), .A3(G290), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(G290), .B1(new_n583), .B2(new_n587), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  XNOR2_X1  g471(.A(G288), .B(G303), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n892), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT42), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n887), .A2(new_n890), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(new_n887), .B2(new_n890), .ZN(new_n902));
  OAI21_X1  g477(.A(G868), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n829), .A2(new_n615), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(G295));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n904), .ZN(G331));
  NAND2_X1  g481(.A1(G301), .A2(G286), .ZN(new_n907));
  NAND2_X1  g482(.A1(G168), .A2(G171), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n884), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n907), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n882), .B2(new_n883), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n830), .A2(KEYINPUT106), .A3(new_n910), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n889), .A2(new_n909), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n909), .A2(new_n911), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n915), .B(new_n899), .C1(new_n881), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n914), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n909), .A2(new_n875), .A3(new_n873), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n888), .A2(KEYINPUT41), .ZN(new_n922));
  INV_X1    g497(.A(new_n880), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n878), .A2(new_n870), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT104), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n921), .B1(new_n926), .B2(new_n916), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n893), .A2(new_n891), .A3(new_n894), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n897), .B1(new_n896), .B2(new_n892), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n895), .A2(new_n898), .A3(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n918), .B(new_n864), .C1(new_n927), .C2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n913), .A2(new_n909), .A3(new_n914), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n888), .A2(new_n870), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n878), .A2(KEYINPUT41), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n920), .B1(new_n830), .B2(new_n910), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n932), .B(new_n931), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  AND4_X1   g517(.A1(KEYINPUT43), .A2(new_n942), .A3(new_n864), .A4(new_n918), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT44), .B1(new_n936), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT108), .B1(new_n934), .B2(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n918), .A2(new_n864), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n926), .A2(new_n916), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n933), .B1(new_n947), .B2(new_n915), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT43), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n942), .A2(new_n935), .A3(new_n864), .A4(new_n918), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n945), .B1(new_n951), .B2(KEYINPUT108), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n944), .B1(new_n952), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n691), .A2(new_n692), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(new_n498), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n469), .A2(KEYINPUT110), .A3(G40), .A4(new_n475), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n960));
  OAI21_X1  g535(.A(G125), .B1(new_n478), .B2(new_n479), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n483), .B1(new_n961), .B2(new_n467), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n472), .B1(new_n478), .B2(new_n479), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n474), .A2(G101), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(G40), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n960), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n959), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n958), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n708), .B(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n742), .B(G2067), .Z(new_n971));
  AND2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n808), .B(new_n810), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(G290), .B(G1986), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT124), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n959), .A2(new_n966), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n496), .A2(new_n497), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n502), .A2(new_n504), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n979), .B(KEYINPUT116), .C1(KEYINPUT45), .C2(new_n982), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n956), .A2(new_n957), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n956), .A2(new_n986), .B1(new_n959), .B2(new_n966), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(KEYINPUT116), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n771), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n990));
  INV_X1    g565(.A(G2084), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n693), .A2(new_n992), .A3(new_n954), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n990), .A2(new_n991), .A3(new_n993), .A4(new_n979), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT117), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n956), .A2(KEYINPUT50), .B1(new_n959), .B2(new_n966), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n991), .A4(new_n993), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n978), .B1(new_n989), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G286), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n989), .A2(G168), .A3(new_n999), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n978), .A2(KEYINPUT120), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1002), .A2(KEYINPUT51), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1001), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n693), .B2(new_n954), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n967), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(new_n695), .A3(new_n984), .A4(new_n983), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT121), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n956), .A2(new_n957), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n987), .B2(KEYINPUT116), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n695), .A4(new_n1010), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(new_n1016), .A3(KEYINPUT53), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n996), .A2(new_n993), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n982), .A2(KEYINPUT45), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n958), .A2(new_n1019), .A3(new_n695), .A4(new_n979), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n777), .A2(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G301), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n958), .A2(new_n1019), .ZN(new_n1024));
  AND4_X1   g599(.A1(KEYINPUT53), .A2(G160), .A3(G40), .A4(new_n695), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT122), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1028), .A3(new_n1025), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1022), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(G171), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1007), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n958), .A2(new_n979), .A3(new_n1019), .ZN(new_n1033));
  INV_X1    g608(.A(G1971), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n996), .A2(new_n757), .A3(new_n993), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n978), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G303), .A2(G8), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT55), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1035), .A2(KEYINPUT111), .A3(new_n1036), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT112), .B(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n978), .B1(new_n979), .B2(new_n982), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1046), .B(new_n1047), .C1(new_n1048), .C2(G288), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G288), .A2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n979), .A2(new_n982), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G8), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT52), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n585), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT113), .B(G86), .Z(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n522), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(G1981), .B1(new_n1057), .B2(new_n582), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n582), .A2(KEYINPUT76), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT76), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1061), .B(new_n542), .C1(new_n580), .C2(new_n581), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n587), .B(new_n1059), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1052), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1058), .A2(new_n1063), .A3(KEYINPUT49), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1054), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1037), .A2(G8), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1041), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1044), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1006), .A2(new_n1032), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1017), .A2(G301), .A3(new_n1022), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT123), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1017), .A2(new_n1075), .A3(G301), .A4(new_n1022), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1007), .B1(new_n1030), .B2(G171), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n977), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1044), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1002), .A2(KEYINPUT51), .A3(new_n1003), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1080), .B1(new_n1085), .B2(new_n1001), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1086), .A2(KEYINPUT124), .A3(new_n1087), .A4(new_n1032), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1018), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT56), .B(G2072), .Z(new_n1090));
  OAI22_X1  g665(.A1(new_n1089), .A2(G1956), .B1(new_n1033), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(G299), .B(KEYINPUT57), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1051), .A2(G2067), .ZN(new_n1098));
  INV_X1    g673(.A(G1348), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1018), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(new_n606), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1024), .A2(new_n969), .A3(new_n979), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n1051), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n549), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1102), .B1(new_n1106), .B2(KEYINPUT59), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(KEYINPUT59), .B2(new_n1106), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1100), .A2(new_n619), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1100), .A2(new_n619), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT60), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1093), .A2(KEYINPUT61), .A3(new_n1094), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1097), .A2(new_n1108), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1093), .A2(new_n1110), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1094), .A3(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1079), .A2(new_n1088), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1085), .A2(new_n1118), .A3(new_n1001), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1117), .A2(new_n1119), .A3(new_n1023), .A4(new_n1071), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1121));
  NOR2_X1   g696(.A1(G288), .A2(G1976), .ZN(new_n1122));
  XOR2_X1   g697(.A(new_n1122), .B(KEYINPUT114), .Z(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1063), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1052), .B1(new_n1125), .B2(KEYINPUT115), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1127), .A3(new_n1063), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1044), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1126), .A2(new_n1128), .B1(new_n1129), .B2(new_n1068), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1000), .A2(G168), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(KEYINPUT63), .A3(new_n1044), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(G8), .A4(new_n1043), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1041), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1068), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT119), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(new_n1068), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1132), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT63), .B1(new_n1071), .B2(new_n1131), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1120), .B(new_n1130), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n976), .B1(new_n1116), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n968), .A2(KEYINPUT46), .A3(new_n969), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT126), .Z(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT46), .B1(new_n968), .B2(new_n969), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT125), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n971), .A2(new_n709), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1150), .A2(new_n968), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1147), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1152), .A2(KEYINPUT47), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(KEYINPUT47), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G290), .A2(G1986), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n968), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n974), .A2(new_n968), .B1(KEYINPUT48), .B2(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1157), .A2(KEYINPUT48), .ZN(new_n1159));
  INV_X1    g734(.A(new_n810), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n808), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n972), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(G2067), .B2(new_n742), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1158), .A2(new_n1159), .B1(new_n1163), .B2(new_n968), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1153), .A2(new_n1154), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT127), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1145), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g742(.A1(G227), .A2(new_n461), .ZN(new_n1169));
  NOR3_X1   g743(.A1(G229), .A2(G401), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g744(.A(new_n859), .B1(new_n854), .B2(new_n855), .ZN(new_n1171));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n1171), .B2(new_n865), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n952), .A2(new_n1172), .ZN(G308));
  INV_X1    g747(.A(KEYINPUT108), .ZN(new_n1174));
  AOI21_X1  g748(.A(new_n1174), .B1(new_n949), .B2(new_n950), .ZN(new_n1175));
  OAI221_X1 g749(.A(new_n1170), .B1(new_n1171), .B2(new_n865), .C1(new_n1175), .C2(new_n945), .ZN(G225));
endmodule


