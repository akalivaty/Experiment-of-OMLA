//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G219), .A2(G218), .A3(G220), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n455), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(KEYINPUT69), .A2(G113), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT69), .B1(G113), .B2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n463), .C1(new_n467), .C2(new_n468), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  MUX2_X1   g054(.A(G100), .B(G112), .S(G2105), .Z(new_n480));
  AOI22_X1  g055(.A1(G136), .A2(new_n479), .B1(new_n480), .B2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n477), .A2(new_n478), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n484), .A2(KEYINPUT70), .A3(G124), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT70), .B1(new_n484), .B2(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n481), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n477), .B2(new_n478), .ZN(new_n490));
  AND2_X1   g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n477), .B2(new_n478), .ZN(new_n494));
  AND2_X1   g069(.A1(G102), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n463), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n463), .C1(new_n467), .C2(new_n468), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n492), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G651), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(G543), .A3(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n508), .A2(new_n511), .A3(new_n509), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n502), .A2(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  OR3_X1    g091(.A1(new_n515), .A2(new_n516), .A3(new_n506), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n515), .B2(new_n506), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(G166));
  INV_X1    g094(.A(new_n512), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  INV_X1    g096(.A(new_n510), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(new_n526), .B1(new_n511), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n521), .A2(new_n523), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n505), .A2(new_n507), .B1(new_n504), .B2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(G52), .A3(G543), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n531), .A2(G90), .A3(new_n511), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n532), .B(new_n533), .C1(new_n506), .C2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n534), .A2(new_n506), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n538), .A2(KEYINPUT73), .A3(new_n532), .A4(new_n533), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  AND2_X1   g116(.A1(KEYINPUT5), .A2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(KEYINPUT5), .A2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g123(.A(KEYINPUT74), .B(new_n541), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G651), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n552), .A2(new_n510), .B1(new_n512), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND4_X1  g136(.A1(new_n508), .A2(G53), .A3(G543), .A4(new_n509), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(G91), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n512), .A2(new_n564), .B1(new_n565), .B2(new_n506), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G166), .ZN(G303));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n506), .B1(new_n544), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n522), .B2(G49), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n508), .A2(G87), .A3(new_n511), .A4(new_n509), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT75), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n531), .A2(new_n576), .A3(G87), .A4(new_n511), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n531), .A2(G86), .A3(new_n511), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n531), .A2(G48), .A3(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n583), .B(G61), .C1(new_n542), .C2(new_n543), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(KEYINPUT77), .A2(G73), .A3(G543), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n584), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n583), .B1(new_n511), .B2(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n582), .B1(KEYINPUT78), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n593), .B(G651), .C1(new_n589), .C2(new_n590), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n522), .A2(G47), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT79), .B(G85), .Z(new_n597));
  NAND2_X1  g172(.A1(new_n520), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n596), .B(new_n598), .C1(new_n506), .C2(new_n599), .ZN(G290));
  NAND3_X1  g175(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n512), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n544), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n601), .A2(new_n604), .B1(G651), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n510), .B(KEYINPUT80), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G54), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G171), .ZN(G284));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G171), .ZN(G321));
  NOR2_X1   g190(.A1(G286), .A2(new_n612), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n566), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n612), .B2(new_n619), .ZN(G297));
  AOI21_X1  g195(.A(new_n616), .B1(new_n612), .B2(new_n619), .ZN(G280));
  INV_X1    g196(.A(new_n611), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR3_X1   g199(.A1(new_n551), .A2(G868), .A3(new_n554), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n611), .A2(G559), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g203(.A(new_n479), .ZN(new_n629));
  OAI21_X1  g204(.A(KEYINPUT12), .B1(new_n629), .B2(new_n476), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT12), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n479), .A2(new_n631), .A3(G2104), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  MUX2_X1   g212(.A(G99), .B(G111), .S(G2105), .Z(new_n638));
  AOI22_X1  g213(.A1(new_n484), .A2(G123), .B1(G2104), .B2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G135), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n629), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n636), .A2(new_n637), .A3(new_n643), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2427), .ZN(new_n648));
  INV_X1    g223(.A(G2430), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT81), .ZN(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT82), .Z(new_n663));
  NOR2_X1   g238(.A1(G2072), .A2(G2078), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n442), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n665), .B(KEYINPUT17), .Z(new_n670));
  OAI211_X1 g245(.A(new_n667), .B(new_n669), .C1(new_n663), .C2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n663), .A3(new_n668), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n665), .A2(new_n668), .A3(new_n662), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n642), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2100), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n679), .A2(KEYINPUT83), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  INV_X1    g261(.A(new_n682), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n679), .B2(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n685), .A2(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n684), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT84), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n693), .B(new_n697), .ZN(G229));
  NOR2_X1   g273(.A1(G6), .A2(G16), .ZN(new_n699));
  INV_X1    g274(.A(G305), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G23), .B(G288), .S(G16), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT85), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G22), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G166), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G1971), .Z(new_n710));
  NAND3_X1  g285(.A1(new_n703), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n713));
  MUX2_X1   g288(.A(G24), .B(G290), .S(G16), .Z(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G1986), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(G1986), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n479), .A2(G131), .ZN(new_n717));
  AND2_X1   g292(.A1(G107), .A2(G2105), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G95), .B2(new_n463), .ZN(new_n719));
  INV_X1    g294(.A(G119), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n717), .B1(new_n476), .B2(new_n719), .C1(new_n720), .C2(new_n483), .ZN(new_n721));
  MUX2_X1   g296(.A(G25), .B(new_n721), .S(G29), .Z(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  NOR4_X1   g300(.A1(new_n715), .A2(new_n716), .A3(new_n725), .A4(KEYINPUT86), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n712), .A2(new_n713), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT87), .B(KEYINPUT36), .Z(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G5), .A2(G16), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT101), .Z(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(G301), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT102), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1961), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G33), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT89), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n479), .A2(G139), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT90), .Z(new_n739));
  NAND3_X1  g314(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT25), .Z(new_n741));
  AOI22_X1  g316(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n739), .B(new_n741), .C1(new_n463), .C2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G29), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n737), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT91), .Z(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(G2072), .ZN(new_n747));
  NOR2_X1   g322(.A1(G16), .A2(G19), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n555), .B2(G16), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n746), .B2(G2072), .ZN(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G35), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G162), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT29), .Z(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n747), .A2(new_n751), .A3(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n744), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT93), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G29), .B2(G160), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G2084), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n763), .A2(G2084), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n732), .A2(G21), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G286), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G27), .A2(G29), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G164), .B2(G29), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT99), .ZN(new_n777));
  INV_X1    g352(.A(G28), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n778), .B2(KEYINPUT30), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(KEYINPUT100), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n780), .A2(KEYINPUT100), .B1(KEYINPUT30), .B2(new_n778), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n777), .B1(new_n781), .B2(new_n782), .C1(new_n641), .C2(new_n744), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n766), .A2(new_n770), .A3(new_n775), .A4(new_n783), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n765), .B(new_n784), .C1(new_n769), .C2(new_n768), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n744), .A2(G26), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT28), .Z(new_n787));
  MUX2_X1   g362(.A(G104), .B(G116), .S(G2105), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G2104), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT88), .Z(new_n790));
  AOI22_X1  g365(.A1(new_n484), .A2(G128), .B1(G140), .B2(new_n479), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n787), .B1(new_n792), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2067), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n774), .B2(new_n773), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n744), .A2(G32), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT97), .B(KEYINPUT26), .Z(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n484), .A2(G129), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT96), .Z(new_n803));
  NAND3_X1  g378(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n479), .A2(G141), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT95), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n797), .B1(new_n808), .B2(new_n744), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT27), .B(G1996), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT98), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n796), .B(new_n812), .C1(new_n755), .C2(new_n754), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n785), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G4), .A2(G16), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n622), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1348), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n732), .A2(G20), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT23), .Z(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G299), .B2(G16), .ZN(new_n820));
  INV_X1    g395(.A(G1956), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  AND4_X1   g398(.A1(new_n735), .A2(new_n757), .A3(new_n814), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n727), .A2(new_n728), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n729), .A2(new_n824), .A3(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n544), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G651), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n531), .A2(G55), .A3(G543), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n531), .A2(G93), .A3(new_n511), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  OAI21_X1  g411(.A(new_n834), .B1(new_n551), .B2(new_n554), .ZN(new_n837));
  INV_X1    g412(.A(new_n834), .ZN(new_n838));
  INV_X1    g413(.A(new_n554), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(new_n839), .A3(new_n550), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n611), .A2(new_n623), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n836), .B1(new_n846), .B2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n641), .B(G160), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G162), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n743), .A2(KEYINPUT103), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n807), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n633), .B(new_n721), .ZN(new_n855));
  MUX2_X1   g430(.A(G106), .B(G118), .S(G2105), .Z(new_n856));
  AOI22_X1  g431(.A1(new_n484), .A2(G130), .B1(G2104), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n479), .A2(KEYINPUT104), .A3(G142), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT104), .B1(new_n479), .B2(G142), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n855), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n792), .B(G164), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n862), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n854), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n853), .A3(new_n863), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n851), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(G37), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n868), .A3(new_n851), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(G395));
  NAND2_X1  g451(.A1(new_n834), .A2(new_n612), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n700), .A2(G166), .ZN(new_n878));
  NAND2_X1  g453(.A1(G305), .A2(G303), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G290), .B(G288), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n879), .A3(new_n878), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT42), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n837), .A2(new_n840), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n626), .B(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n608), .A2(new_n619), .A3(new_n610), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n619), .B1(new_n608), .B2(new_n610), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n888), .A2(KEYINPUT107), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT41), .B1(new_n890), .B2(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n611), .A2(G299), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n889), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT107), .B1(new_n888), .B2(new_n893), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n894), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n886), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n886), .B2(new_n902), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n886), .A2(new_n902), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n877), .B1(new_n907), .B2(new_n612), .ZN(G295));
  OAI21_X1  g483(.A(new_n877), .B1(new_n907), .B2(new_n612), .ZN(G331));
  AOI21_X1  g484(.A(G286), .B1(new_n537), .B2(new_n539), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n537), .A2(G286), .A3(new_n539), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n841), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n887), .B1(new_n914), .B2(new_n910), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n899), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n892), .A3(new_n915), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n885), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G37), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n885), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n895), .A2(new_n898), .B1(new_n913), .B2(new_n915), .ZN(new_n923));
  INV_X1    g498(.A(new_n918), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(KEYINPUT43), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n919), .A2(new_n920), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n895), .A2(new_n929), .A3(new_n898), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n892), .A2(KEYINPUT109), .A3(new_n897), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n916), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n885), .B1(new_n932), .B2(new_n918), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n927), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT44), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n936));
  INV_X1    g511(.A(new_n933), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n921), .B2(new_n937), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n928), .A2(new_n933), .A3(KEYINPUT110), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n921), .A2(new_n927), .A3(new_n925), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n935), .B1(new_n942), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n945));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n500), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n500), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G125), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n477), .B2(new_n478), .ZN(new_n951));
  NAND2_X1  g526(.A1(G113), .A2(G2104), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT69), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(KEYINPUT69), .A2(G113), .A3(G2104), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(G2105), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n472), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n479), .B2(G137), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n959), .A3(G40), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT112), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n957), .A2(new_n959), .A3(new_n962), .A4(G40), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n949), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n808), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n792), .A2(G2067), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n790), .A2(new_n794), .A3(new_n791), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n965), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(new_n966), .A3(new_n808), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n972), .A2(KEYINPUT113), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(KEYINPUT113), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT114), .B(new_n971), .C1(new_n973), .C2(new_n974), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n721), .A2(new_n724), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n721), .A2(new_n724), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n965), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  NOR2_X1   g558(.A1(G290), .A2(G1986), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n965), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(G286), .A2(G8), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT125), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT50), .B1(new_n500), .B2(new_n946), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n500), .A2(KEYINPUT50), .A3(new_n946), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n964), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT118), .B(G2084), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n500), .A2(new_n946), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n944), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n961), .A3(new_n963), .A4(new_n997), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n992), .A2(new_n994), .B1(new_n998), .B2(new_n769), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT51), .B(new_n988), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n962), .B1(G160), .B2(G40), .ZN(new_n1003));
  INV_X1    g578(.A(new_n963), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n500), .A2(KEYINPUT50), .A3(new_n946), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1005), .B(new_n994), .C1(new_n989), .C2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n997), .A2(new_n961), .A3(new_n963), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n500), .B2(new_n946), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n769), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1000), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT125), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n987), .B(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1002), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n1013), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1001), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1005), .A2(new_n774), .A3(new_n996), .A4(new_n997), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1008), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1021), .A2(KEYINPUT53), .A3(new_n774), .A4(new_n996), .ZN(new_n1022));
  INV_X1    g597(.A(G1961), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1006), .A2(new_n989), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n964), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1020), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G171), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n960), .A2(new_n1019), .A3(G2078), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1028), .A2(new_n997), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1018), .A2(new_n1019), .B1(new_n949), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT126), .B1(new_n992), .B2(G1961), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT126), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1032), .B(new_n1023), .C1(new_n1024), .C2(new_n964), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1030), .A2(G301), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT54), .B1(new_n1027), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n580), .A2(new_n581), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1036), .A2(new_n1037), .A3(new_n594), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n591), .ZN(new_n1040));
  OAI21_X1  g615(.A(G1981), .B1(new_n1040), .B2(new_n582), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1039), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT49), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n961), .A2(new_n946), .A3(new_n500), .A4(new_n963), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n573), .A2(new_n578), .A3(G1976), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(G8), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT117), .B(G1976), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(G288), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1051), .A2(G8), .A3(new_n1044), .A4(new_n1047), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n1055));
  OR3_X1    g630(.A1(G166), .A2(new_n1000), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(G166), .B2(new_n1000), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT115), .B(G1971), .Z(new_n1059));
  AOI22_X1  g634(.A1(new_n992), .A2(new_n755), .B1(new_n998), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1060), .B2(new_n1000), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n998), .A2(new_n1059), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1005), .B(new_n755), .C1(new_n989), .C2(new_n1006), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(G8), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1054), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1035), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n949), .A2(new_n1029), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1031), .A2(new_n1020), .A3(new_n1069), .A4(new_n1033), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1005), .B1(new_n989), .B2(new_n1006), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1019), .A2(new_n1018), .B1(new_n1072), .B2(new_n1023), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(G301), .A3(new_n1022), .ZN(new_n1074));
  AND4_X1   g649(.A1(KEYINPUT127), .A2(new_n1071), .A3(KEYINPUT54), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1070), .B2(G171), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT127), .B1(new_n1077), .B2(new_n1074), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1017), .B(new_n1068), .C1(new_n1075), .C2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G299), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n619), .A2(KEYINPUT57), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1005), .A2(new_n996), .A3(new_n997), .A4(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1084), .B(new_n1086), .C1(new_n992), .C2(G1956), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT122), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1072), .A2(new_n821), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1086), .A4(new_n1084), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1086), .B1(new_n992), .B2(G1956), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1084), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1080), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1087), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1008), .A2(G1996), .A3(new_n1009), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  AND2_X1   g676(.A1(new_n1044), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n555), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT59), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1105), .B(new_n555), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1099), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT124), .B1(new_n1096), .B2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1087), .A2(new_n1098), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1084), .B1(new_n1089), .B2(new_n1086), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1110), .B(new_n1111), .C1(new_n1113), .C2(new_n1080), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1044), .A2(G2067), .ZN(new_n1115));
  INV_X1    g690(.A(G1348), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1072), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n611), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n611), .B(KEYINPUT60), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1118), .A2(KEYINPUT60), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1109), .A2(new_n1114), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1092), .B1(new_n1118), .B2(new_n1112), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1079), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n1000), .B(G286), .C1(new_n1007), .C2(new_n1010), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1054), .A2(new_n1061), .A3(new_n1066), .A4(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT120), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1054), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1129), .A2(KEYINPUT121), .A3(KEYINPUT63), .A4(new_n1124), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1125), .A2(new_n1134), .A3(new_n1126), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1128), .A2(new_n1130), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1046), .ZN(new_n1137));
  NOR2_X1   g712(.A1(G288), .A2(G1976), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1137), .A2(new_n1138), .B1(new_n1037), .B2(new_n700), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1054), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1139), .A2(new_n1045), .B1(new_n1140), .B2(new_n1066), .ZN(new_n1141));
  AOI21_X1  g716(.A(G301), .B1(new_n1073), .B2(new_n1022), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1142), .A2(new_n1054), .A3(new_n1061), .A4(new_n1066), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1001), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1141), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1136), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n986), .B1(new_n1123), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT46), .ZN(new_n1151));
  INV_X1    g726(.A(new_n965), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(G1996), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n965), .A2(KEYINPUT46), .A3(new_n966), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n965), .B1(new_n807), .B2(new_n970), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT47), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n965), .A2(new_n984), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT48), .Z(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n982), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1152), .B1(new_n1161), .B2(new_n969), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1150), .A2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g739(.A1(G401), .A2(G229), .A3(new_n461), .A4(G227), .ZN(new_n1166));
  NAND4_X1  g740(.A1(new_n874), .A2(new_n1166), .A3(new_n934), .A4(new_n926), .ZN(G225));
  INV_X1    g741(.A(G225), .ZN(G308));
endmodule


