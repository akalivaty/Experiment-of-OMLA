

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n746), .ZN(n765) );
  BUF_X1 U553 ( .A(n746), .Z(n784) );
  INV_X1 U554 ( .A(G2104), .ZN(n575) );
  NOR2_X1 U555 ( .A1(n763), .A2(n762), .ZN(n531) );
  NAND2_X1 U556 ( .A1(n742), .A2(n741), .ZN(n746) );
  NOR2_X2 U557 ( .A1(n575), .A2(G2105), .ZN(n910) );
  OR2_X1 U558 ( .A1(n772), .A2(G168), .ZN(n528) );
  NOR2_X1 U559 ( .A1(n535), .A2(n532), .ZN(n771) );
  INV_X1 U560 ( .A(n740), .ZN(n742) );
  INV_X1 U561 ( .A(KEYINPUT102), .ZN(n547) );
  NAND2_X1 U562 ( .A1(n575), .A2(n554), .ZN(n553) );
  INV_X1 U563 ( .A(G2105), .ZN(n554) );
  INV_X1 U564 ( .A(G1966), .ZN(n543) );
  INV_X1 U565 ( .A(KEYINPUT92), .ZN(n538) );
  AND2_X1 U566 ( .A1(n541), .A2(KEYINPUT92), .ZN(n540) );
  NAND2_X1 U567 ( .A1(n534), .A2(n533), .ZN(n532) );
  NAND2_X1 U568 ( .A1(n784), .A2(n542), .ZN(n534) );
  NAND2_X1 U569 ( .A1(n784), .A2(n538), .ZN(n533) );
  AND2_X1 U570 ( .A1(n543), .A2(G8), .ZN(n542) );
  NAND2_X1 U571 ( .A1(n539), .A2(n536), .ZN(n535) );
  AND2_X1 U572 ( .A1(G8), .A2(n537), .ZN(n536) );
  NAND2_X1 U573 ( .A1(n765), .A2(n540), .ZN(n539) );
  NAND2_X1 U574 ( .A1(n538), .A2(G2084), .ZN(n537) );
  XNOR2_X1 U575 ( .A(n527), .B(KEYINPUT31), .ZN(n526) );
  NAND2_X1 U576 ( .A1(n528), .A2(n520), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n784), .A2(G8), .ZN(n812) );
  NAND2_X1 U578 ( .A1(n546), .A2(n522), .ZN(n545) );
  NAND2_X1 U579 ( .A1(n519), .A2(n518), .ZN(n544) );
  AND2_X1 U580 ( .A1(n574), .A2(n521), .ZN(n525) );
  AND2_X1 U581 ( .A1(n802), .A2(n522), .ZN(n518) );
  AND2_X1 U582 ( .A1(n552), .A2(n524), .ZN(n519) );
  OR2_X1 U583 ( .A1(G171), .A2(n773), .ZN(n520) );
  AND2_X1 U584 ( .A1(n577), .A2(n576), .ZN(n521) );
  AND2_X1 U585 ( .A1(n573), .A2(n525), .ZN(G160) );
  NAND2_X1 U586 ( .A1(G160), .A2(G40), .ZN(n740) );
  AND2_X1 U587 ( .A1(n832), .A2(n825), .ZN(n522) );
  NOR2_X1 U588 ( .A1(n810), .A2(n812), .ZN(n523) );
  AND2_X1 U589 ( .A1(n801), .A2(n547), .ZN(n524) );
  INV_X1 U590 ( .A(G2084), .ZN(n541) );
  NAND2_X1 U591 ( .A1(n529), .A2(n526), .ZN(n790) );
  NAND2_X1 U592 ( .A1(n530), .A2(n769), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n531), .B(KEYINPUT29), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n545), .A2(n544), .ZN(n820) );
  NAND2_X1 U595 ( .A1(n548), .A2(n550), .ZN(n546) );
  NAND2_X1 U596 ( .A1(n549), .A2(KEYINPUT102), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n552), .A2(n801), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n551), .A2(KEYINPUT102), .ZN(n550) );
  INV_X1 U599 ( .A(n802), .ZN(n551) );
  NAND2_X1 U600 ( .A1(n818), .A2(n817), .ZN(n552) );
  XNOR2_X2 U601 ( .A(n553), .B(KEYINPUT17), .ZN(n909) );
  XNOR2_X1 U602 ( .A(KEYINPUT30), .B(KEYINPUT95), .ZN(n770) );
  XNOR2_X1 U603 ( .A(n771), .B(n770), .ZN(n772) );
  INV_X1 U604 ( .A(KEYINPUT103), .ZN(n819) );
  XOR2_X1 U605 ( .A(KEYINPUT15), .B(n599), .Z(n990) );
  XOR2_X1 U606 ( .A(G543), .B(KEYINPUT0), .Z(n656) );
  NOR2_X2 U607 ( .A1(G651), .A2(n656), .ZN(n668) );
  NAND2_X1 U608 ( .A1(G53), .A2(n668), .ZN(n557) );
  INV_X1 U609 ( .A(G651), .ZN(n558) );
  NOR2_X1 U610 ( .A1(G543), .A2(n558), .ZN(n555) );
  XOR2_X1 U611 ( .A(KEYINPUT1), .B(n555), .Z(n667) );
  NAND2_X1 U612 ( .A1(G65), .A2(n667), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n563) );
  NOR2_X2 U614 ( .A1(n656), .A2(n558), .ZN(n672) );
  NAND2_X1 U615 ( .A1(n672), .A2(G78), .ZN(n561) );
  NOR2_X1 U616 ( .A1(G651), .A2(G543), .ZN(n559) );
  XNOR2_X1 U617 ( .A(n559), .B(KEYINPUT64), .ZN(n669) );
  NAND2_X1 U618 ( .A1(G91), .A2(n669), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U620 ( .A1(n563), .A2(n562), .ZN(G299) );
  NAND2_X1 U621 ( .A1(G52), .A2(n668), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G64), .A2(n667), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U624 ( .A1(n672), .A2(G77), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G90), .A2(n669), .ZN(n566) );
  NAND2_X1 U626 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U627 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U628 ( .A1(n570), .A2(n569), .ZN(G171) );
  AND2_X1 U629 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U630 ( .A(G57), .ZN(G237) );
  INV_X1 U631 ( .A(G132), .ZN(G219) );
  NAND2_X1 U632 ( .A1(G101), .A2(n910), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT23), .B(n571), .Z(n574) );
  NAND2_X1 U634 ( .A1(G137), .A2(n909), .ZN(n572) );
  XOR2_X1 U635 ( .A(n572), .B(KEYINPUT65), .Z(n573) );
  AND2_X1 U636 ( .A1(n575), .A2(G2105), .ZN(n905) );
  NAND2_X1 U637 ( .A1(G125), .A2(n905), .ZN(n577) );
  AND2_X1 U638 ( .A1(G2104), .A2(G2105), .ZN(n906) );
  NAND2_X1 U639 ( .A1(G113), .A2(n906), .ZN(n576) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U642 ( .A(G223), .ZN(n842) );
  NAND2_X1 U643 ( .A1(n842), .A2(G567), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  NAND2_X1 U645 ( .A1(G43), .A2(n668), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n580), .B(KEYINPUT70), .ZN(n587) );
  NAND2_X1 U647 ( .A1(G81), .A2(n669), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G68), .A2(n672), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT69), .B(KEYINPUT13), .Z(n584) );
  XNOR2_X1 U652 ( .A(n585), .B(n584), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n667), .A2(G56), .ZN(n588) );
  XOR2_X1 U655 ( .A(KEYINPUT14), .B(n588), .Z(n589) );
  NOR2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U657 ( .A(KEYINPUT71), .B(n591), .ZN(n997) );
  INV_X1 U658 ( .A(G860), .ZN(n637) );
  OR2_X1 U659 ( .A1(n997), .A2(n637), .ZN(G153) );
  INV_X1 U660 ( .A(G171), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U662 ( .A1(G79), .A2(n672), .ZN(n593) );
  NAND2_X1 U663 ( .A1(G54), .A2(n668), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U665 ( .A(n594), .B(KEYINPUT72), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n667), .A2(G66), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G92), .A2(n669), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  OR2_X1 U670 ( .A1(n990), .A2(G868), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n601), .A2(n600), .ZN(G284) );
  NAND2_X1 U672 ( .A1(n669), .A2(G89), .ZN(n602) );
  XOR2_X1 U673 ( .A(KEYINPUT73), .B(n602), .Z(n603) );
  XNOR2_X1 U674 ( .A(n603), .B(KEYINPUT4), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G76), .A2(n672), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT5), .ZN(n611) );
  NAND2_X1 U678 ( .A1(G51), .A2(n668), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G63), .A2(n667), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U681 ( .A(KEYINPUT6), .B(n609), .Z(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n612), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U684 ( .A(G168), .B(KEYINPUT8), .Z(n613) );
  XNOR2_X1 U685 ( .A(KEYINPUT74), .B(n613), .ZN(G286) );
  XNOR2_X1 U686 ( .A(KEYINPUT75), .B(G868), .ZN(n614) );
  NOR2_X1 U687 ( .A1(G286), .A2(n614), .ZN(n616) );
  NOR2_X1 U688 ( .A1(G868), .A2(G299), .ZN(n615) );
  NOR2_X1 U689 ( .A1(n616), .A2(n615), .ZN(G297) );
  NAND2_X1 U690 ( .A1(G559), .A2(n637), .ZN(n617) );
  XNOR2_X1 U691 ( .A(KEYINPUT76), .B(n617), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n618), .A2(n990), .ZN(n619) );
  XNOR2_X1 U693 ( .A(KEYINPUT16), .B(n619), .ZN(G148) );
  INV_X1 U694 ( .A(G868), .ZN(n687) );
  NOR2_X1 U695 ( .A1(G559), .A2(n687), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n990), .A2(n620), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT77), .ZN(n623) );
  NOR2_X1 U698 ( .A1(n997), .A2(G868), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U700 ( .A1(n906), .A2(G111), .ZN(n624) );
  XOR2_X1 U701 ( .A(KEYINPUT79), .B(n624), .Z(n626) );
  NAND2_X1 U702 ( .A1(n910), .A2(G99), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U704 ( .A(KEYINPUT80), .B(n627), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n905), .A2(G123), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT18), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G135), .A2(n909), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U709 ( .A(KEYINPUT78), .B(n631), .ZN(n632) );
  NOR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n1011) );
  XNOR2_X1 U711 ( .A(n1011), .B(G2096), .ZN(n635) );
  INV_X1 U712 ( .A(G2100), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(G156) );
  NAND2_X1 U714 ( .A1(G559), .A2(n990), .ZN(n636) );
  XOR2_X1 U715 ( .A(n997), .B(n636), .Z(n684) );
  NAND2_X1 U716 ( .A1(n637), .A2(n684), .ZN(n645) );
  NAND2_X1 U717 ( .A1(n668), .A2(G55), .ZN(n639) );
  NAND2_X1 U718 ( .A1(G93), .A2(n669), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G80), .A2(n672), .ZN(n640) );
  XNOR2_X1 U721 ( .A(KEYINPUT81), .B(n640), .ZN(n641) );
  NOR2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n667), .A2(G67), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n686) );
  XNOR2_X1 U725 ( .A(n645), .B(n686), .ZN(G145) );
  NAND2_X1 U726 ( .A1(n672), .A2(G75), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G88), .A2(n669), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G50), .A2(n668), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G62), .A2(n667), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U732 ( .A1(n651), .A2(n650), .ZN(G166) );
  INV_X1 U733 ( .A(G166), .ZN(G303) );
  NAND2_X1 U734 ( .A1(G49), .A2(n668), .ZN(n653) );
  NAND2_X1 U735 ( .A1(G74), .A2(G651), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U737 ( .A1(n667), .A2(n654), .ZN(n655) );
  XNOR2_X1 U738 ( .A(n655), .B(KEYINPUT82), .ZN(n658) );
  NAND2_X1 U739 ( .A1(G87), .A2(n656), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(G288) );
  NAND2_X1 U741 ( .A1(n668), .A2(G47), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n672), .A2(G72), .ZN(n660) );
  NAND2_X1 U743 ( .A1(G85), .A2(n669), .ZN(n659) );
  NAND2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U745 ( .A1(G60), .A2(n667), .ZN(n661) );
  XOR2_X1 U746 ( .A(KEYINPUT66), .B(n661), .Z(n662) );
  NOR2_X1 U747 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U748 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U749 ( .A(KEYINPUT67), .B(n666), .Z(G290) );
  NAND2_X1 U750 ( .A1(n667), .A2(G61), .ZN(n677) );
  NAND2_X1 U751 ( .A1(n668), .A2(G48), .ZN(n671) );
  NAND2_X1 U752 ( .A1(G86), .A2(n669), .ZN(n670) );
  NAND2_X1 U753 ( .A1(n671), .A2(n670), .ZN(n675) );
  NAND2_X1 U754 ( .A1(n672), .A2(G73), .ZN(n673) );
  XOR2_X1 U755 ( .A(KEYINPUT2), .B(n673), .Z(n674) );
  NOR2_X1 U756 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U757 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U758 ( .A(KEYINPUT83), .B(n678), .Z(G305) );
  XNOR2_X1 U759 ( .A(KEYINPUT19), .B(G303), .ZN(n679) );
  XNOR2_X1 U760 ( .A(n679), .B(G288), .ZN(n680) );
  XNOR2_X1 U761 ( .A(n680), .B(G299), .ZN(n681) );
  XNOR2_X1 U762 ( .A(n681), .B(n686), .ZN(n682) );
  XNOR2_X1 U763 ( .A(n682), .B(G290), .ZN(n683) );
  XNOR2_X1 U764 ( .A(n683), .B(G305), .ZN(n922) );
  XNOR2_X1 U765 ( .A(n684), .B(n922), .ZN(n685) );
  NAND2_X1 U766 ( .A1(n685), .A2(G868), .ZN(n689) );
  NAND2_X1 U767 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U768 ( .A1(n689), .A2(n688), .ZN(G295) );
  NAND2_X1 U769 ( .A1(G2078), .A2(G2084), .ZN(n690) );
  XOR2_X1 U770 ( .A(KEYINPUT20), .B(n690), .Z(n691) );
  NAND2_X1 U771 ( .A1(G2090), .A2(n691), .ZN(n693) );
  XNOR2_X1 U772 ( .A(KEYINPUT21), .B(KEYINPUT84), .ZN(n692) );
  XNOR2_X1 U773 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U774 ( .A1(G2072), .A2(n694), .ZN(G158) );
  XNOR2_X1 U775 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U776 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  NOR2_X1 U777 ( .A1(G220), .A2(G219), .ZN(n695) );
  XOR2_X1 U778 ( .A(KEYINPUT22), .B(n695), .Z(n696) );
  NOR2_X1 U779 ( .A1(G218), .A2(n696), .ZN(n697) );
  NAND2_X1 U780 ( .A1(G96), .A2(n697), .ZN(n846) );
  NAND2_X1 U781 ( .A1(G2106), .A2(n846), .ZN(n701) );
  NAND2_X1 U782 ( .A1(G69), .A2(G120), .ZN(n698) );
  NOR2_X1 U783 ( .A1(G237), .A2(n698), .ZN(n699) );
  NAND2_X1 U784 ( .A1(G108), .A2(n699), .ZN(n847) );
  NAND2_X1 U785 ( .A1(G567), .A2(n847), .ZN(n700) );
  NAND2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n848) );
  NAND2_X1 U787 ( .A1(G661), .A2(G483), .ZN(n702) );
  NOR2_X1 U788 ( .A1(n848), .A2(n702), .ZN(n845) );
  NAND2_X1 U789 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U790 ( .A1(G138), .A2(n909), .ZN(n704) );
  NAND2_X1 U791 ( .A1(G102), .A2(n910), .ZN(n703) );
  NAND2_X1 U792 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U793 ( .A1(G126), .A2(n905), .ZN(n706) );
  NAND2_X1 U794 ( .A1(G114), .A2(n906), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U796 ( .A1(n708), .A2(n707), .ZN(G164) );
  NOR2_X1 U797 ( .A1(G164), .A2(G1384), .ZN(n741) );
  NOR2_X1 U798 ( .A1(n741), .A2(n740), .ZN(n837) );
  NAND2_X1 U799 ( .A1(G140), .A2(n909), .ZN(n711) );
  NAND2_X1 U800 ( .A1(G104), .A2(n910), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U802 ( .A(KEYINPUT34), .B(n712), .ZN(n718) );
  NAND2_X1 U803 ( .A1(G128), .A2(n905), .ZN(n714) );
  NAND2_X1 U804 ( .A1(G116), .A2(n906), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U806 ( .A(KEYINPUT35), .B(n715), .ZN(n716) );
  XNOR2_X1 U807 ( .A(KEYINPUT85), .B(n716), .ZN(n717) );
  NOR2_X1 U808 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U809 ( .A(KEYINPUT36), .B(n719), .ZN(n892) );
  XNOR2_X1 U810 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NOR2_X1 U811 ( .A1(n892), .A2(n824), .ZN(n1008) );
  NAND2_X1 U812 ( .A1(n837), .A2(n1008), .ZN(n832) );
  NAND2_X1 U813 ( .A1(G119), .A2(n905), .ZN(n720) );
  XNOR2_X1 U814 ( .A(n720), .B(KEYINPUT86), .ZN(n727) );
  NAND2_X1 U815 ( .A1(G131), .A2(n909), .ZN(n722) );
  NAND2_X1 U816 ( .A1(G107), .A2(n906), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U818 ( .A1(G95), .A2(n910), .ZN(n723) );
  XNOR2_X1 U819 ( .A(KEYINPUT87), .B(n723), .ZN(n724) );
  NOR2_X1 U820 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U821 ( .A1(n727), .A2(n726), .ZN(n891) );
  NAND2_X1 U822 ( .A1(G1991), .A2(n891), .ZN(n728) );
  XNOR2_X1 U823 ( .A(n728), .B(KEYINPUT88), .ZN(n738) );
  NAND2_X1 U824 ( .A1(G105), .A2(n910), .ZN(n729) );
  XNOR2_X1 U825 ( .A(n729), .B(KEYINPUT38), .ZN(n736) );
  NAND2_X1 U826 ( .A1(G141), .A2(n909), .ZN(n731) );
  NAND2_X1 U827 ( .A1(G129), .A2(n905), .ZN(n730) );
  NAND2_X1 U828 ( .A1(n731), .A2(n730), .ZN(n734) );
  NAND2_X1 U829 ( .A1(G117), .A2(n906), .ZN(n732) );
  XNOR2_X1 U830 ( .A(KEYINPUT89), .B(n732), .ZN(n733) );
  NOR2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U832 ( .A1(n736), .A2(n735), .ZN(n916) );
  NAND2_X1 U833 ( .A1(G1996), .A2(n916), .ZN(n737) );
  NAND2_X1 U834 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U835 ( .A(KEYINPUT90), .B(n739), .ZN(n1031) );
  NAND2_X1 U836 ( .A1(n837), .A2(n1031), .ZN(n825) );
  INV_X1 U837 ( .A(G1348), .ZN(n934) );
  NOR2_X1 U838 ( .A1(n765), .A2(n934), .ZN(n744) );
  AND2_X1 U839 ( .A1(n765), .A2(G2067), .ZN(n743) );
  NOR2_X1 U840 ( .A1(n744), .A2(n743), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n990), .A2(n750), .ZN(n754) );
  INV_X1 U842 ( .A(G1996), .ZN(n962) );
  NOR2_X1 U843 ( .A1(n746), .A2(n962), .ZN(n745) );
  XOR2_X1 U844 ( .A(n745), .B(KEYINPUT26), .Z(n748) );
  NAND2_X1 U845 ( .A1(n784), .A2(G1341), .ZN(n747) );
  NAND2_X1 U846 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U847 ( .A1(n997), .A2(n749), .ZN(n752) );
  AND2_X1 U848 ( .A1(n990), .A2(n750), .ZN(n751) );
  NOR2_X1 U849 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U850 ( .A1(n754), .A2(n753), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n765), .A2(G2072), .ZN(n755) );
  XOR2_X1 U852 ( .A(KEYINPUT27), .B(n755), .Z(n757) );
  NAND2_X1 U853 ( .A1(G1956), .A2(n784), .ZN(n756) );
  NAND2_X1 U854 ( .A1(n757), .A2(n756), .ZN(n760) );
  NOR2_X1 U855 ( .A1(G299), .A2(n760), .ZN(n758) );
  NOR2_X1 U856 ( .A1(n759), .A2(n758), .ZN(n763) );
  NAND2_X1 U857 ( .A1(G299), .A2(n760), .ZN(n761) );
  XOR2_X1 U858 ( .A(KEYINPUT28), .B(n761), .Z(n762) );
  OR2_X1 U859 ( .A1(n765), .A2(G1961), .ZN(n767) );
  XOR2_X1 U860 ( .A(G2078), .B(KEYINPUT25), .Z(n764) );
  XNOR2_X1 U861 ( .A(KEYINPUT93), .B(n764), .ZN(n959) );
  NAND2_X1 U862 ( .A1(n765), .A2(n959), .ZN(n766) );
  NAND2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n773) );
  AND2_X1 U864 ( .A1(n773), .A2(G171), .ZN(n768) );
  XOR2_X1 U865 ( .A(KEYINPUT94), .B(n768), .Z(n769) );
  NAND2_X1 U866 ( .A1(n790), .A2(G286), .ZN(n774) );
  XNOR2_X1 U867 ( .A(n774), .B(KEYINPUT96), .ZN(n780) );
  NOR2_X1 U868 ( .A1(G1971), .A2(n812), .ZN(n776) );
  NOR2_X1 U869 ( .A1(G2090), .A2(n784), .ZN(n775) );
  NOR2_X1 U870 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U871 ( .A1(n777), .A2(G303), .ZN(n778) );
  XOR2_X1 U872 ( .A(KEYINPUT97), .B(n778), .Z(n779) );
  NAND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n781), .A2(G8), .ZN(n782) );
  XNOR2_X1 U875 ( .A(n782), .B(KEYINPUT32), .ZN(n792) );
  NAND2_X1 U876 ( .A1(KEYINPUT92), .A2(G1966), .ZN(n783) );
  NAND2_X1 U877 ( .A1(n783), .A2(n784), .ZN(n787) );
  XNOR2_X1 U878 ( .A(KEYINPUT92), .B(n541), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n785), .A2(n765), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n788), .A2(G8), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n809) );
  NOR2_X1 U884 ( .A1(G2090), .A2(G303), .ZN(n793) );
  XNOR2_X1 U885 ( .A(KEYINPUT100), .B(n793), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n794), .A2(G8), .ZN(n795) );
  XOR2_X1 U887 ( .A(KEYINPUT101), .B(n795), .Z(n796) );
  NAND2_X1 U888 ( .A1(n809), .A2(n796), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n797), .A2(n812), .ZN(n802) );
  NOR2_X1 U890 ( .A1(G1981), .A2(G305), .ZN(n798) );
  XNOR2_X1 U891 ( .A(n798), .B(KEYINPUT91), .ZN(n799) );
  XNOR2_X1 U892 ( .A(KEYINPUT24), .B(n799), .ZN(n800) );
  OR2_X1 U893 ( .A1(n812), .A2(n800), .ZN(n801) );
  NOR2_X1 U894 ( .A1(G288), .A2(G1976), .ZN(n803) );
  XNOR2_X1 U895 ( .A(n803), .B(KEYINPUT98), .ZN(n984) );
  NOR2_X1 U896 ( .A1(G1971), .A2(G303), .ZN(n804) );
  XOR2_X1 U897 ( .A(n804), .B(KEYINPUT99), .Z(n805) );
  NOR2_X1 U898 ( .A1(n984), .A2(n805), .ZN(n807) );
  INV_X1 U899 ( .A(KEYINPUT33), .ZN(n806) );
  AND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n818) );
  NAND2_X1 U902 ( .A1(G1976), .A2(G288), .ZN(n991) );
  INV_X1 U903 ( .A(n991), .ZN(n810) );
  OR2_X1 U904 ( .A1(KEYINPUT33), .A2(n523), .ZN(n816) );
  INV_X1 U905 ( .A(n984), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U907 ( .A1(KEYINPUT33), .A2(n813), .ZN(n814) );
  XNOR2_X1 U908 ( .A(G1981), .B(G305), .ZN(n982) );
  NOR2_X1 U909 ( .A1(n814), .A2(n982), .ZN(n815) );
  AND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U911 ( .A(n820), .B(n819), .ZN(n822) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n985) );
  NAND2_X1 U913 ( .A1(n837), .A2(n985), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U915 ( .A(n823), .B(KEYINPUT104), .ZN(n840) );
  AND2_X1 U916 ( .A1(n892), .A2(n824), .ZN(n1009) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n916), .ZN(n1023) );
  INV_X1 U918 ( .A(n825), .ZN(n829) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n891), .ZN(n1019) );
  NOR2_X1 U920 ( .A1(G1986), .A2(G290), .ZN(n826) );
  XOR2_X1 U921 ( .A(n826), .B(KEYINPUT105), .Z(n827) );
  NOR2_X1 U922 ( .A1(n1019), .A2(n827), .ZN(n828) );
  NOR2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U924 ( .A1(n1023), .A2(n830), .ZN(n831) );
  XNOR2_X1 U925 ( .A(KEYINPUT39), .B(n831), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U927 ( .A(KEYINPUT106), .B(n834), .Z(n835) );
  NOR2_X1 U928 ( .A1(n1009), .A2(n835), .ZN(n836) );
  XNOR2_X1 U929 ( .A(KEYINPUT107), .B(n836), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U932 ( .A(n841), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U935 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U937 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  NOR2_X1 U942 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U944 ( .A(KEYINPUT109), .B(n848), .ZN(G319) );
  XNOR2_X1 U945 ( .A(G1348), .B(G2454), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n849), .B(G2430), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n850), .B(G1341), .ZN(n856) );
  XOR2_X1 U948 ( .A(G2443), .B(G2427), .Z(n852) );
  XNOR2_X1 U949 ( .A(G2438), .B(G2446), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n854) );
  XOR2_X1 U951 ( .A(G2451), .B(G2435), .Z(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n857) );
  NAND2_X1 U954 ( .A1(n857), .A2(G14), .ZN(n858) );
  XOR2_X1 U955 ( .A(KEYINPUT108), .B(n858), .Z(G401) );
  XOR2_X1 U956 ( .A(G2100), .B(G2096), .Z(n860) );
  XNOR2_X1 U957 ( .A(KEYINPUT42), .B(G2678), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U959 ( .A(KEYINPUT43), .B(G2090), .Z(n862) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2072), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U963 ( .A(G2078), .B(G2084), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(G227) );
  XOR2_X1 U965 ( .A(G2474), .B(KEYINPUT110), .Z(n868) );
  XNOR2_X1 U966 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(n869), .B(KEYINPUT111), .Z(n871) );
  XNOR2_X1 U969 ( .A(G1996), .B(G1991), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n879) );
  XOR2_X1 U971 ( .A(G1976), .B(G1971), .Z(n873) );
  XNOR2_X1 U972 ( .A(G1986), .B(G1961), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n877) );
  XOR2_X1 U974 ( .A(KEYINPUT112), .B(G1981), .Z(n875) );
  XNOR2_X1 U975 ( .A(G1956), .B(G1966), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(n877), .B(n876), .Z(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(G229) );
  NAND2_X1 U979 ( .A1(G100), .A2(n910), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G112), .A2(n906), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G124), .A2(n905), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n882), .B(KEYINPUT44), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G136), .A2(n909), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n883), .B(KEYINPUT114), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n886) );
  NOR2_X1 U987 ( .A1(n887), .A2(n886), .ZN(G162) );
  XOR2_X1 U988 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n889) );
  XNOR2_X1 U989 ( .A(G162), .B(KEYINPUT48), .ZN(n888) );
  XNOR2_X1 U990 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U991 ( .A(G164), .B(n890), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n891), .B(n1011), .ZN(n894) );
  XOR2_X1 U993 ( .A(G160), .B(n892), .Z(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n920) );
  NAND2_X1 U996 ( .A1(G139), .A2(n909), .ZN(n898) );
  NAND2_X1 U997 ( .A1(G103), .A2(n910), .ZN(n897) );
  NAND2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n904) );
  NAND2_X1 U999 ( .A1(G127), .A2(n905), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n906), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1002 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  XNOR2_X1 U1003 ( .A(KEYINPUT116), .B(n902), .ZN(n903) );
  NOR2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n1012) );
  NAND2_X1 U1005 ( .A1(G130), .A2(n905), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(G118), .A2(n906), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n915) );
  NAND2_X1 U1008 ( .A1(G142), .A2(n909), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(G106), .A2(n910), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1011 ( .A(n913), .B(KEYINPUT45), .Z(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1014 ( .A(n1012), .B(n918), .Z(n919) );
  XNOR2_X1 U1015 ( .A(n920), .B(n919), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n921), .ZN(G395) );
  XNOR2_X1 U1017 ( .A(G286), .B(n922), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(n990), .B(G171), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(n924), .B(n923), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(n925), .B(n997), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(G37), .A2(n926), .ZN(G397) );
  INV_X1 U1022 ( .A(G401), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(G319), .A2(n927), .ZN(n930) );
  NOR2_X1 U1024 ( .A1(G227), .A2(G229), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT49), .B(n928), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1031 ( .A(G5), .B(G1961), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(n933), .B(KEYINPUT123), .ZN(n948) );
  XNOR2_X1 U1033 ( .A(G1966), .B(G21), .ZN(n946) );
  XNOR2_X1 U1034 ( .A(KEYINPUT59), .B(G4), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(n935), .B(n934), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(G1341), .B(G19), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(G1981), .B(G6), .ZN(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n938), .B(KEYINPUT125), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1041 ( .A(G1956), .B(KEYINPUT124), .Z(n941) );
  XNOR2_X1 U1042 ( .A(G20), .B(n941), .ZN(n942) );
  NAND2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT60), .B(n944), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(G1971), .B(G22), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(G23), .B(G1976), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n952) );
  XOR2_X1 U1050 ( .A(G1986), .B(G24), .Z(n951) );
  NAND2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n953), .ZN(n954) );
  NOR2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1054 ( .A(n956), .B(KEYINPUT61), .Z(n957) );
  XNOR2_X1 U1055 ( .A(KEYINPUT126), .B(n957), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(G16), .A2(n958), .ZN(n1039) );
  INV_X1 U1057 ( .A(KEYINPUT55), .ZN(n1033) );
  XOR2_X1 U1058 ( .A(G27), .B(n959), .Z(n969) );
  XNOR2_X1 U1059 ( .A(G2067), .B(G26), .ZN(n961) );
  XNOR2_X1 U1060 ( .A(G33), .B(G2072), .ZN(n960) );
  NOR2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(G32), .B(n962), .ZN(n963) );
  NAND2_X1 U1063 ( .A1(n963), .A2(G28), .ZN(n965) );
  XNOR2_X1 U1064 ( .A(G25), .B(G1991), .ZN(n964) );
  NOR2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n970) );
  XNOR2_X1 U1069 ( .A(n971), .B(n970), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(G35), .B(G2090), .ZN(n972) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(G34), .B(KEYINPUT54), .ZN(n974) );
  XNOR2_X1 U1073 ( .A(n974), .B(n541), .ZN(n975) );
  NAND2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1075 ( .A(n1033), .B(n977), .ZN(n979) );
  INV_X1 U1076 ( .A(G29), .ZN(n978) );
  NAND2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1078 ( .A1(G11), .A2(n980), .ZN(n1007) );
  XOR2_X1 U1079 ( .A(G16), .B(KEYINPUT56), .Z(n1004) );
  XOR2_X1 U1080 ( .A(G1966), .B(G168), .Z(n981) );
  NOR2_X1 U1081 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1082 ( .A(KEYINPUT57), .B(n983), .Z(n1001) );
  NOR2_X1 U1083 ( .A1(n985), .A2(n984), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(G171), .B(G1961), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(G299), .B(G1956), .ZN(n987) );
  XNOR2_X1 U1086 ( .A(G303), .B(G1971), .ZN(n986) );
  NOR2_X1 U1087 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1088 ( .A1(n989), .A2(n988), .ZN(n994) );
  XNOR2_X1 U1089 ( .A(n990), .B(G1348), .ZN(n992) );
  NAND2_X1 U1090 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1091 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(G1341), .B(n997), .ZN(n998) );
  NOR2_X1 U1094 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1096 ( .A(n1002), .B(KEYINPUT121), .ZN(n1003) );
  NOR2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1098 ( .A(n1005), .B(KEYINPUT122), .ZN(n1006) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1037) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1029) );
  XNOR2_X1 U1101 ( .A(G160), .B(n541), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1021) );
  XOR2_X1 U1103 ( .A(n1012), .B(KEYINPUT118), .Z(n1013) );
  XOR2_X1 U1104 ( .A(G2072), .B(n1013), .Z(n1015) );
  XNOR2_X1 U1105 ( .A(G2078), .B(G164), .ZN(n1014) );
  NAND2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1107 ( .A(n1016), .B(KEYINPUT119), .Z(n1017) );
  XNOR2_X1 U1108 ( .A(KEYINPUT50), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(G2090), .B(G162), .ZN(n1022) );
  XNOR2_X1 U1112 ( .A(n1022), .B(KEYINPUT117), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1114 ( .A(KEYINPUT51), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1118 ( .A(KEYINPUT52), .B(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1120 ( .A1(n1035), .A2(G29), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1122 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1123 ( .A(KEYINPUT62), .B(n1040), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

