//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT78), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G140), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(new_n195), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G104), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(G107), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n196), .A2(new_n199), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n195), .A2(G107), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n198), .A2(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(G101), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n206), .B1(G128), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(G146), .ZN(new_n213));
  AND4_X1   g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(G128), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n202), .B(new_n205), .C1(new_n209), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT10), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n202), .A2(new_n205), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n210), .B1(G143), .B2(new_n211), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(KEYINPUT68), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n208), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n206), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n219), .B(KEYINPUT10), .C1(new_n225), .C2(new_n214), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n212), .A2(new_n213), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT0), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n220), .A3(KEYINPUT64), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT64), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(KEYINPUT0), .B2(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n212), .A2(new_n213), .B1(KEYINPUT0), .B2(G128), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n229), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n196), .A2(new_n199), .A3(new_n201), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G101), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n240), .A3(G101), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G134), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G137), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(G137), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n244), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G137), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G134), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT11), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(G131), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n249), .A2(G134), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n250), .B2(new_n252), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n251), .A2(KEYINPUT11), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n245), .B1(new_n247), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT66), .B(G131), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n217), .A2(new_n226), .A3(new_n242), .A4(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(G128), .B1(new_n208), .B2(new_n223), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT68), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n227), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n214), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n218), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n215), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n270), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT12), .B1(new_n270), .B2(new_n262), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n264), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n194), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n264), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n217), .A2(new_n226), .A3(new_n242), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n262), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n194), .A2(new_n273), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n190), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n271), .B2(new_n272), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n270), .A2(new_n262), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT12), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n270), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(KEYINPUT77), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n283), .A2(new_n288), .A3(new_n275), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n277), .A2(new_n264), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n194), .ZN(new_n291));
  AOI211_X1 g105(.A(G469), .B(G902), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n281), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G221), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT76), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n294), .B1(new_n297), .B2(new_n280), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT6), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n302));
  INV_X1    g116(.A(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G116), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G113), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(G116), .B(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n302), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT2), .B(G113), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n218), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n314), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n306), .A2(KEYINPUT2), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G113), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n308), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n319), .A2(new_n324), .A3(KEYINPUT69), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT69), .B1(new_n319), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n327), .A2(KEYINPUT79), .A3(new_n239), .A4(new_n241), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n323), .A2(new_n308), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(new_n315), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n319), .A2(new_n324), .A3(KEYINPUT69), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n239), .A3(new_n332), .A4(new_n241), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n318), .B1(new_n328), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G122), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n301), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n333), .A2(new_n334), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n333), .A2(new_n334), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n317), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n337), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n234), .A2(new_n227), .A3(new_n228), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n206), .A2(KEYINPUT0), .A3(G128), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT81), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n212), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n224), .A2(G128), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n214), .B1(new_n351), .B2(new_n227), .ZN(new_n352));
  INV_X1    g166(.A(G125), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n347), .A2(new_n355), .A3(G125), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n349), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n192), .A2(G224), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT82), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n357), .B(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n341), .A2(new_n301), .A3(new_n342), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n344), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT83), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n344), .A2(new_n365), .A3(new_n361), .A4(new_n362), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n315), .B1(new_n307), .B2(new_n309), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n218), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT5), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n307), .B1(new_n372), .B2(new_n313), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n316), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT84), .B1(new_n368), .B2(new_n219), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n337), .B(KEYINPUT8), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n357), .A2(new_n360), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n376), .A2(new_n377), .B1(new_n378), .B2(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n336), .A2(new_n337), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n354), .A2(KEYINPUT85), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n348), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n354), .A2(KEYINPUT85), .ZN(new_n383));
  XOR2_X1   g197(.A(KEYINPUT86), .B(KEYINPUT7), .Z(new_n384));
  OAI22_X1  g198(.A1(new_n382), .A2(new_n383), .B1(new_n360), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n379), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n280), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n300), .B1(new_n367), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n300), .ZN(new_n390));
  AOI211_X1 g204(.A(new_n390), .B(new_n387), .C1(new_n364), .C2(new_n366), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n189), .B(new_n299), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n331), .A2(new_n332), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n244), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n243), .A2(KEYINPUT67), .A3(G137), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n250), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G131), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n261), .B(new_n399), .C1(new_n225), .C2(new_n214), .ZN(new_n400));
  INV_X1    g214(.A(new_n260), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n248), .A2(new_n401), .A3(new_n254), .ZN(new_n402));
  INV_X1    g216(.A(G131), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n257), .B2(new_n259), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n236), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n394), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n405), .A3(new_n394), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT71), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT28), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT71), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n409), .A2(new_n412), .B1(new_n410), .B2(new_n408), .ZN(new_n413));
  NOR2_X1   g227(.A1(G237), .A2(G953), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G210), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT27), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT26), .B(G101), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n408), .A2(new_n418), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT70), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n261), .A2(new_n399), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(new_n352), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n347), .B1(new_n261), .B2(new_n255), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT30), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n400), .A2(new_n405), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n422), .B1(new_n429), .B2(new_n327), .ZN(new_n430));
  AOI211_X1 g244(.A(KEYINPUT70), .B(new_n394), .C1(new_n426), .C2(new_n428), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n421), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT31), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n400), .A2(new_n405), .A3(new_n427), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n427), .B1(new_n400), .B2(new_n405), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n327), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT70), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n429), .A2(new_n422), .A3(new_n327), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT31), .A3(new_n421), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n419), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(G472), .A2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT32), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n413), .A2(new_n418), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT31), .B1(new_n440), .B2(new_n421), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n433), .B(new_n420), .C1(new_n438), .C2(new_n439), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT32), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n443), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT29), .B1(new_n413), .B2(new_n418), .ZN(new_n452));
  INV_X1    g266(.A(new_n408), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n438), .B2(new_n439), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n418), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n407), .A2(KEYINPUT72), .A3(new_n408), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT72), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n406), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n458), .A3(KEYINPUT28), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n408), .A2(new_n410), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n459), .A2(KEYINPUT29), .A3(new_n418), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n280), .A3(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n445), .A2(new_n451), .B1(new_n462), .B2(G472), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT22), .B(G137), .ZN(new_n464));
  INV_X1    g278(.A(G234), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n294), .A2(new_n465), .A3(G953), .ZN(new_n466));
  XOR2_X1   g280(.A(new_n464), .B(new_n466), .Z(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n303), .A2(G128), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT74), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n303), .A2(G128), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT24), .B(G110), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT23), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(new_n303), .B2(G128), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT75), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(KEYINPUT75), .A3(new_n476), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G110), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT16), .ZN(new_n485));
  INV_X1    g299(.A(G140), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(G125), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(G125), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n353), .A2(G140), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(G146), .B(new_n487), .C1(new_n490), .C2(new_n485), .ZN(new_n491));
  XNOR2_X1  g305(.A(G125), .B(G140), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n211), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n484), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI22_X1  g308(.A1(new_n473), .A2(new_n474), .B1(new_n481), .B2(new_n482), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n487), .B1(new_n490), .B2(new_n485), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n211), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n497), .A2(new_n491), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n468), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n499), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n484), .A2(new_n491), .A3(new_n493), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(new_n467), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n503), .A3(new_n280), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT25), .A4(new_n280), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G217), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(G234), .B2(new_n280), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT73), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n500), .A2(new_n503), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n510), .A2(G902), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n508), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n463), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(KEYINPUT87), .A2(G143), .ZN(new_n517));
  NOR2_X1   g331(.A1(KEYINPUT87), .A2(G143), .ZN(new_n518));
  OAI211_X1 g332(.A(G214), .B(new_n414), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G237), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n192), .A3(G214), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT87), .A2(G143), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n401), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n260), .A3(new_n523), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(KEYINPUT17), .A3(new_n401), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n498), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(G113), .B(G122), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(G104), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT90), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT89), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n519), .A2(new_n536), .A3(new_n523), .ZN(new_n537));
  NAND2_X1  g351(.A1(KEYINPUT18), .A2(G131), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n519), .A2(new_n523), .A3(new_n536), .A4(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n490), .A2(G146), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n493), .ZN(new_n543));
  AND4_X1   g357(.A1(new_n535), .A2(new_n540), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n537), .A2(new_n539), .B1(new_n493), .B2(new_n542), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n535), .B1(new_n545), .B2(new_n541), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n530), .B(new_n534), .C1(new_n544), .C2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n532), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n530), .B1(new_n544), .B2(new_n546), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(KEYINPUT92), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT92), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n530), .B(new_n552), .C1(new_n544), .C2(new_n546), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n548), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT93), .B1(new_n554), .B2(G902), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT89), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n545), .A2(new_n535), .A3(new_n541), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n529), .A2(new_n497), .A3(new_n491), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(new_n528), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n532), .B1(new_n560), .B2(new_n552), .ZN(new_n561));
  INV_X1    g375(.A(new_n553), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n547), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n280), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT91), .B(G475), .Z(new_n566));
  NAND3_X1  g380(.A1(new_n555), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n525), .A2(new_n527), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n492), .B(KEYINPUT19), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n211), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n570), .A3(new_n491), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n544), .B2(new_n546), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n532), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n547), .ZN(new_n574));
  NOR2_X1   g388(.A1(G475), .A2(G902), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT20), .ZN(new_n577));
  INV_X1    g391(.A(G952), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(G953), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n465), .B2(new_n520), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n280), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT21), .B(G898), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT95), .ZN(new_n585));
  XNOR2_X1  g399(.A(G116), .B(G122), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n198), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n220), .A2(G143), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n207), .A2(G128), .ZN(new_n591));
  OR3_X1    g405(.A1(new_n590), .A2(new_n591), .A3(G134), .ZN(new_n592));
  OAI21_X1  g406(.A(G134), .B1(new_n590), .B2(new_n591), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT14), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n586), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n311), .A2(G122), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n198), .B1(new_n596), .B2(KEYINPUT14), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n592), .A2(new_n593), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n586), .B(new_n198), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n220), .A2(G143), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n590), .B2(KEYINPUT13), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(KEYINPUT13), .B2(new_n590), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n600), .B(new_n592), .C1(new_n603), .C2(new_n243), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n296), .A2(new_n509), .A3(G953), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n599), .A2(new_n606), .A3(new_n604), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT15), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G478), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n609), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n606), .B1(new_n599), .B2(new_n604), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n280), .B(new_n612), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n585), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n280), .B1(new_n614), .B2(new_n615), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n611), .A3(G478), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT95), .A3(new_n616), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n584), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n567), .A2(new_n577), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT96), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n393), .A2(new_n516), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  NAND2_X1  g440(.A1(new_n449), .A2(new_n443), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n442), .B2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT97), .ZN(new_n629));
  INV_X1    g443(.A(new_n298), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n514), .B(new_n630), .C1(new_n292), .C2(new_n281), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n633), .B(G472), .C1(new_n442), .C2(G902), .ZN(new_n634));
  AND4_X1   g448(.A1(new_n627), .A2(new_n629), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT98), .Z(new_n636));
  OAI211_X1 g450(.A(KEYINPUT33), .B(new_n609), .C1(new_n608), .C2(KEYINPUT100), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n608), .A2(KEYINPUT100), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n608), .B2(new_n609), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(G478), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(G902), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n642), .A2(new_n644), .B1(new_n643), .B2(new_n619), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n567), .B2(new_n577), .ZN(new_n646));
  INV_X1    g460(.A(new_n584), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n647), .B(new_n189), .C1(new_n389), .C2(new_n391), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n636), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NAND3_X1  g466(.A1(new_n576), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n567), .B(new_n653), .C1(new_n577), .C2(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n618), .A2(new_n621), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n636), .A2(new_n649), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT102), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT35), .B(G107), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n623), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n392), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n629), .A2(new_n627), .A3(new_n634), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n508), .A2(new_n511), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n501), .A2(new_n502), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n468), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n513), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NOR2_X1   g489(.A1(new_n463), .A2(new_n671), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n582), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n580), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n654), .A2(new_n655), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n393), .A2(new_n676), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NAND2_X1  g497(.A1(new_n567), .A2(new_n577), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n655), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n189), .A3(new_n671), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n679), .B(KEYINPUT39), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n299), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n687), .B1(KEYINPUT40), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n445), .A2(new_n451), .ZN(new_n691));
  INV_X1    g505(.A(new_n418), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n454), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n456), .A2(new_n458), .ZN(new_n694));
  AOI21_X1  g508(.A(G902), .B1(new_n694), .B2(new_n692), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n690), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n367), .A2(new_n388), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n390), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n367), .A2(new_n300), .A3(new_n388), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT38), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  INV_X1    g523(.A(new_n645), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n684), .A2(new_n710), .A3(new_n679), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n393), .A2(new_n676), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  NAND4_X1  g528(.A1(new_n705), .A2(new_n647), .A3(new_n189), .A4(new_n646), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n462), .A2(G472), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n442), .A2(KEYINPUT32), .A3(new_n444), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n450), .B1(new_n449), .B2(new_n443), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n289), .A2(new_n291), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n190), .B1(new_n720), .B2(new_n280), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n292), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT103), .B1(new_n722), .B2(new_n630), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NOR4_X1   g538(.A1(new_n721), .A2(new_n292), .A3(new_n724), .A4(new_n298), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n719), .A2(new_n514), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n715), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT41), .B(G113), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND4_X1  g544(.A1(new_n705), .A2(new_n647), .A3(new_n189), .A4(new_n656), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n727), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n311), .ZN(G18));
  OAI21_X1  g547(.A(new_n189), .B1(new_n389), .B2(new_n391), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n720), .A2(new_n280), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n720), .A2(new_n190), .A3(new_n280), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n630), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n724), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n722), .A2(KEYINPUT103), .A3(new_n630), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n624), .A3(new_n676), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  OAI211_X1 g558(.A(new_n686), .B(new_n189), .C1(new_n389), .C2(new_n391), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n447), .A2(new_n448), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n418), .B1(new_n459), .B2(new_n460), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n443), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n628), .A2(new_n749), .A3(new_n514), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n741), .A2(new_n750), .A3(new_n584), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n746), .A2(KEYINPUT104), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  INV_X1    g567(.A(new_n750), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n647), .A3(new_n726), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n753), .B1(new_n755), .B2(new_n745), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  NAND2_X1  g572(.A1(new_n711), .A2(KEYINPUT105), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n646), .A2(new_n760), .A3(new_n679), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n628), .A2(new_n749), .A3(new_n670), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n742), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G125), .ZN(G27));
  NAND4_X1  g579(.A1(new_n703), .A2(new_n189), .A3(new_n704), .A4(new_n299), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n768));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n762), .A3(new_n516), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n719), .A2(new_n514), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n759), .A2(new_n761), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n770), .A2(new_n771), .A3(new_n766), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(KEYINPUT106), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n769), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  NAND3_X1  g590(.A1(new_n767), .A2(new_n516), .A3(new_n681), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NAND2_X1  g592(.A1(new_n685), .A2(new_n710), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n664), .A3(new_n670), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT107), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n703), .A2(new_n189), .A3(new_n704), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n278), .A2(KEYINPUT45), .ZN(new_n789));
  OAI21_X1  g603(.A(G469), .B1(new_n278), .B2(KEYINPUT45), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n789), .A2(new_n790), .B1(new_n190), .B2(new_n280), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n292), .B1(new_n791), .B2(new_n792), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n298), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n788), .A2(new_n795), .A3(new_n688), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n783), .B2(new_n782), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n786), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  AND2_X1   g613(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n788), .A2(new_n463), .A3(new_n515), .A4(new_n712), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT108), .B(G140), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G42));
  NOR2_X1   g620(.A1(new_n613), .A2(new_n617), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n685), .A2(KEYINPUT111), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n684), .B2(new_n807), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n809), .B(new_n811), .C1(new_n685), .C2(new_n645), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n635), .A2(new_n649), .A3(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n673), .A2(new_n813), .A3(new_n625), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n727), .B1(new_n715), .B2(new_n731), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n624), .A2(new_n719), .A3(new_n670), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n705), .A2(new_n189), .A3(new_n726), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n814), .A2(new_n819), .A3(new_n757), .A4(new_n775), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n767), .A2(new_n762), .A3(new_n763), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n777), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n654), .A2(new_n808), .A3(new_n680), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n719), .A2(new_n670), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT112), .B1(new_n825), .B2(new_n766), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n767), .A2(new_n676), .A3(new_n827), .A4(new_n824), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n822), .A2(new_n823), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n826), .A2(new_n828), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n821), .A2(new_n777), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT113), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n820), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n670), .A2(new_n680), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n684), .A3(new_n621), .A4(new_n618), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n691), .B2(new_n697), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n393), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n764), .A2(new_n682), .A3(new_n713), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(KEYINPUT114), .A3(new_n840), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n713), .A2(new_n838), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(KEYINPUT52), .A3(new_n682), .A4(new_n764), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n834), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n833), .A2(new_n830), .ZN(new_n849));
  INV_X1    g663(.A(new_n820), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n841), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT54), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n463), .A2(new_n741), .A3(new_n515), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n856), .B(new_n649), .C1(new_n646), .C2(new_n656), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n663), .B1(new_n672), .B2(new_n516), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n743), .A4(new_n813), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n752), .A2(new_n756), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n822), .A2(new_n823), .A3(new_n829), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n823), .B1(new_n822), .B2(new_n829), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n861), .B(new_n775), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n851), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n852), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n834), .A2(KEYINPUT53), .A3(new_n847), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n787), .A2(new_n741), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n515), .A2(new_n580), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n646), .A3(new_n698), .A4(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n872), .A2(new_n579), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n779), .B(KEYINPUT43), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n874), .A2(new_n580), .A3(new_n750), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n742), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n580), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n516), .A3(new_n870), .ZN(new_n878));
  XOR2_X1   g692(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n879));
  OAI211_X1 g693(.A(new_n873), .B(new_n876), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(KEYINPUT48), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n880), .B1(new_n882), .B2(new_n878), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n877), .A2(new_n763), .A3(new_n870), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n684), .A2(new_n710), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n870), .A2(new_n698), .A3(new_n871), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n877), .A2(new_n754), .A3(new_n788), .ZN(new_n887));
  INV_X1    g701(.A(new_n722), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n630), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n800), .A2(new_n801), .A3(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n884), .B(new_n886), .C1(new_n887), .C2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT50), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n741), .A2(new_n189), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n707), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n875), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n893), .B1(new_n707), .B2(new_n894), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n707), .A2(new_n894), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT116), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(KEYINPUT50), .A3(new_n875), .A4(new_n895), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n891), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n883), .B1(new_n902), .B2(KEYINPUT51), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT51), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n904), .B(new_n891), .C1(new_n898), .C2(new_n901), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n855), .A2(new_n869), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n578), .A2(new_n192), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OR4_X1    g723(.A1(new_n515), .A2(new_n779), .A3(new_n188), .A4(new_n298), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n910), .A2(KEYINPUT109), .B1(KEYINPUT49), .B2(new_n888), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(KEYINPUT109), .B2(new_n910), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT110), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n888), .A2(KEYINPUT49), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(new_n707), .A3(new_n698), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT118), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n909), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(G75));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n866), .A2(new_n867), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(G902), .ZN(new_n923));
  INV_X1    g737(.A(G210), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n344), .A2(new_n362), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(new_n361), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n925), .A2(new_n928), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n192), .A2(G952), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(G51));
  NOR2_X1   g746(.A1(new_n789), .A2(new_n790), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n922), .A2(G902), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT119), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n190), .A2(new_n280), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT57), .Z(new_n940));
  OAI21_X1  g754(.A(new_n720), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n931), .B1(new_n935), .B2(new_n941), .ZN(G54));
  INV_X1    g756(.A(new_n931), .ZN(new_n943));
  AND4_X1   g757(.A1(KEYINPUT58), .A2(new_n922), .A3(G475), .A4(G902), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n574), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n574), .B2(new_n944), .ZN(G60));
  XOR2_X1   g760(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n947));
  NOR2_X1   g761(.A1(new_n643), .A2(new_n280), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n642), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(new_n869), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT121), .B1(new_n952), .B2(new_n931), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT121), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n954), .B(new_n943), .C1(new_n938), .C2(new_n950), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n855), .A2(new_n869), .ZN(new_n956));
  INV_X1    g770(.A(new_n949), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n956), .A2(new_n957), .B1(new_n639), .B2(new_n641), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n953), .A2(new_n955), .A3(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT122), .Z(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT60), .Z(new_n962));
  NAND3_X1  g776(.A1(new_n922), .A2(new_n668), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n866), .B2(new_n867), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n963), .B(new_n943), .C1(new_n512), .C2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n967), .A3(new_n943), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n966), .A2(new_n968), .A3(KEYINPUT61), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n965), .A2(new_n512), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n931), .B1(new_n965), .B2(new_n668), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n970), .B(new_n971), .C1(new_n967), .C2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n969), .A2(new_n973), .ZN(G66));
  INV_X1    g788(.A(G224), .ZN(new_n975));
  OAI21_X1  g789(.A(G953), .B1(new_n583), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n861), .B2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n926), .B1(G898), .B2(new_n192), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G69));
  AOI21_X1  g793(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n429), .B(new_n569), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n804), .B1(new_n786), .B2(new_n797), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n764), .A2(new_n682), .A3(new_n713), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n708), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n812), .A2(KEYINPUT124), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n770), .A2(new_n766), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n812), .A2(KEYINPUT124), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n987), .A2(new_n688), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n982), .A2(new_n985), .A3(new_n986), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n981), .B1(new_n991), .B2(new_n192), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n746), .A2(new_n516), .A3(new_n688), .A4(new_n795), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n982), .A2(new_n983), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n775), .A2(new_n777), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT126), .Z(new_n997));
  NOR3_X1   g811(.A1(new_n995), .A2(G953), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n981), .B1(new_n677), .B2(new_n192), .ZN(new_n999));
  OAI22_X1  g813(.A1(new_n992), .A2(new_n993), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n992), .A2(new_n993), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n980), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n992), .A2(new_n993), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n998), .A2(new_n999), .ZN(new_n1005));
  INV_X1    g819(.A(new_n980), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1001), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1003), .A2(new_n1007), .ZN(G72));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  OR2_X1    g824(.A1(new_n995), .A2(new_n997), .ZN(new_n1011));
  INV_X1    g825(.A(new_n861), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n454), .A2(new_n692), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1010), .B1(new_n991), .B2(new_n1012), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1018), .B(new_n1010), .C1(new_n991), .C2(new_n1012), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1017), .A2(new_n693), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n432), .B1(new_n454), .B2(new_n418), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n1010), .B(new_n1021), .C1(new_n848), .C2(new_n854), .ZN(new_n1022));
  AND4_X1   g836(.A1(new_n943), .A2(new_n1015), .A3(new_n1020), .A4(new_n1022), .ZN(G57));
endmodule


