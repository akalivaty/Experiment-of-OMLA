//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n204), .A2(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT77), .ZN(new_n211));
  OAI22_X1  g010(.A1(new_n206), .A2(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT78), .B1(new_n204), .B2(G148gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(G141gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n221), .A3(new_n205), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n216), .B1(new_n215), .B2(KEYINPUT2), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n212), .A2(new_n217), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G134gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G127gat), .ZN(new_n226));
  INV_X1    g025(.A(G127gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G134gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT70), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(KEYINPUT70), .A3(G134gat), .ZN(new_n231));
  INV_X1    g030(.A(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G113gat), .ZN(new_n233));
  INV_X1    g032(.A(G113gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G120gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n230), .A2(new_n231), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n226), .A2(new_n228), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n236), .A2(new_n239), .A3(new_n237), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT79), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT1), .B1(new_n233), .B2(new_n235), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n239), .ZN(new_n244));
  INV_X1    g043(.A(new_n231), .ZN(new_n245));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(new_n229), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n242), .B(new_n244), .C1(new_n247), .C2(new_n243), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n224), .B1(new_n241), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n238), .A2(new_n240), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n212), .A2(new_n217), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n223), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n203), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n244), .B1(new_n247), .B2(new_n243), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n224), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(new_n258), .B2(new_n224), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n224), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n248), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n230), .A2(new_n231), .ZN(new_n267));
  INV_X1    g066(.A(new_n243), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n242), .B1(new_n269), .B2(new_n244), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n263), .B(new_n265), .C1(new_n266), .C2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n262), .A2(new_n271), .A3(new_n202), .ZN(new_n272));
  OAI211_X1 g071(.A(KEYINPUT81), .B(new_n203), .C1(new_n249), .C2(new_n254), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n272), .A3(KEYINPUT5), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n224), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n254), .A2(new_n260), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n271), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n203), .A2(KEYINPUT5), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n283));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n281), .A3(new_n287), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT91), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n274), .B2(new_n281), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT6), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT91), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n289), .A2(new_n296), .A3(new_n290), .A4(new_n291), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n293), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299));
  INV_X1    g098(.A(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(G218gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n299), .B1(KEYINPUT22), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G211gat), .B(G218gat), .Z(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT67), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(G169gat), .A3(G176gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n316), .A2(KEYINPUT69), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT69), .B1(new_n316), .B2(new_n317), .ZN(new_n319));
  INV_X1    g118(.A(G183gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT27), .B1(new_n320), .B2(KEYINPUT68), .ZN(new_n321));
  INV_X1    g120(.A(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G183gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n321), .B(new_n322), .C1(KEYINPUT68), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT27), .B(G183gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(G190gat), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n318), .A2(new_n319), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n311), .A2(KEYINPUT25), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n317), .A2(KEYINPUT24), .ZN(new_n337));
  NOR2_X1   g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(KEYINPUT66), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n331), .A2(new_n333), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n343), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n341), .A2(new_n311), .A3(new_n342), .A4(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n340), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G226gat), .ZN(new_n349));
  INV_X1    g148(.A(G233gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n330), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(KEYINPUT29), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n345), .A2(new_n347), .ZN(new_n354));
  INV_X1    g153(.A(new_n340), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n308), .A2(new_n310), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n315), .A2(new_n312), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n317), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n325), .A2(new_n326), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n327), .A2(new_n328), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n316), .A2(KEYINPUT69), .A3(new_n317), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n353), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n306), .B1(new_n352), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n353), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n330), .B2(new_n348), .ZN(new_n370));
  INV_X1    g169(.A(new_n351), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n320), .A2(new_n322), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT24), .A3(new_n317), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n343), .B1(new_n373), .B2(new_n336), .ZN(new_n374));
  INV_X1    g173(.A(new_n344), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n342), .A2(new_n311), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n346), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n371), .B(new_n366), .C1(new_n378), .C2(new_n340), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n370), .A2(new_n379), .A3(new_n305), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n368), .A2(KEYINPUT92), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT92), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n370), .A2(new_n379), .A3(new_n382), .A4(new_n305), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(KEYINPUT37), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT37), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n385), .A3(new_n380), .ZN(new_n386));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT76), .ZN(new_n388));
  INV_X1    g187(.A(G64gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G92gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(KEYINPUT38), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n384), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n368), .A2(new_n380), .A3(new_n392), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n385), .B1(new_n368), .B2(new_n380), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT93), .B1(new_n397), .B2(new_n392), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n370), .A2(new_n379), .A3(new_n305), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n305), .B1(new_n370), .B2(new_n379), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT37), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT93), .ZN(new_n402));
  INV_X1    g201(.A(new_n392), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n404), .A3(new_n386), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n396), .B1(KEYINPUT38), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n298), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT85), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT31), .B(G50gat), .Z(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(G22gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(KEYINPUT86), .A2(G22gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n416), .B(KEYINPUT87), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n415), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n305), .B1(new_n265), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n264), .B1(new_n306), .B2(KEYINPUT29), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(new_n253), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n418), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT89), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n249), .A2(new_n254), .A3(new_n203), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT39), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n253), .B1(new_n266), .B2(new_n270), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n202), .A3(new_n275), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(KEYINPUT89), .A3(KEYINPUT39), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n279), .A2(new_n203), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n279), .A2(new_n426), .A3(new_n203), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n287), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT40), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n289), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n433), .A2(new_n287), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT90), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n434), .A2(new_n441), .A3(new_n435), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n436), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n403), .B1(new_n399), .B2(new_n400), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n395), .A3(KEYINPUT30), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n368), .A2(new_n446), .A3(new_n380), .A4(new_n392), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(KEYINPUT88), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n423), .B1(new_n443), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(KEYINPUT83), .A2(KEYINPUT6), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n274), .A2(new_n281), .A3(new_n287), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(new_n294), .ZN(new_n456));
  INV_X1    g255(.A(new_n454), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n289), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n458), .A3(new_n448), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n456), .A2(new_n458), .A3(new_n448), .A4(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n407), .A2(new_n453), .B1(new_n463), .B2(new_n423), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n250), .B1(new_n330), .B2(new_n348), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT72), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT72), .B(new_n250), .C1(new_n330), .C2(new_n348), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n258), .B(new_n366), .C1(new_n378), .C2(new_n340), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT71), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT71), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n356), .A2(new_n472), .A3(new_n258), .A4(new_n366), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G227gat), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n469), .B(new_n474), .C1(new_n475), .C2(new_n350), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT34), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n467), .A2(new_n468), .B1(new_n471), .B2(new_n473), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n475), .A2(new_n350), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n479), .B(KEYINPUT64), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(KEYINPUT34), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G43gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT73), .ZN(new_n486));
  INV_X1    g285(.A(G71gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G99gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n486), .A2(new_n487), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n487), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(G99gat), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n469), .A2(new_n474), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n481), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT33), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(KEYINPUT32), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n480), .B1(new_n469), .B2(new_n474), .ZN(new_n501));
  INV_X1    g300(.A(new_n493), .ZN(new_n502));
  AOI21_X1  g301(.A(G99gat), .B1(new_n491), .B2(new_n492), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT74), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT74), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n505), .A3(new_n493), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(KEYINPUT33), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n501), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n484), .B1(new_n500), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT75), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n493), .B(new_n490), .C1(new_n501), .C2(new_n498), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n476), .A2(KEYINPUT34), .B1(new_n478), .B2(new_n482), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n496), .A2(KEYINPUT32), .A3(new_n507), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n511), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(KEYINPUT75), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n511), .A2(KEYINPUT36), .A3(new_n516), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n517), .A2(new_n519), .ZN(new_n523));
  INV_X1    g322(.A(new_n423), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n293), .A2(new_n295), .A3(new_n297), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT94), .B(KEYINPUT35), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n452), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n523), .A2(new_n524), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n524), .A3(new_n516), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT35), .B1(new_n463), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n464), .A2(new_n522), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n532));
  NAND2_X1  g331(.A1(G43gat), .A2(G50gat), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT95), .B(G43gat), .Z(new_n534));
  OAI211_X1 g333(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(G50gat), .ZN(new_n535));
  OR2_X1    g334(.A1(G43gat), .A2(G50gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n532), .B1(new_n536), .B2(new_n533), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G29gat), .ZN(new_n540));
  INV_X1    g339(.A(G36gat), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT14), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  MUX2_X1   g342(.A(new_n542), .B(KEYINPUT14), .S(new_n543), .Z(new_n544));
  NOR2_X1   g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n538), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT17), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT105), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(G85gat), .A3(G92gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  INV_X1    g352(.A(G85gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(KEYINPUT8), .A2(new_n553), .B1(new_n554), .B2(new_n391), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n549), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G99gat), .B(G106gat), .Z(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT106), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n558), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n546), .C1(new_n539), .C2(new_n544), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT103), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n545), .A2(new_n547), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n561), .A3(new_n562), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(G190gat), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n566), .A2(new_n572), .A3(new_n322), .A4(new_n570), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(G218gat), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(G218gat), .B1(new_n574), .B2(new_n575), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT107), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT107), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n576), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT104), .B(G134gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G162gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n583), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n579), .A2(new_n582), .A3(new_n587), .ZN(new_n588));
  OAI211_X1 g387(.A(KEYINPUT107), .B(new_n586), .C1(new_n577), .C2(new_n578), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G15gat), .B(G22gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT16), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n592), .B2(G1gat), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(G1gat), .B2(new_n591), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(G8gat), .Z(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT98), .B(G57gat), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n596), .A2(new_n389), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n389), .ZN(new_n598));
  NAND2_X1  g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n597), .B(new_n598), .C1(KEYINPUT9), .C2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n605), .A2(KEYINPUT97), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(KEYINPUT97), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n601), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT100), .B(G64gat), .Z(new_n609));
  NAND2_X1  g408(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT9), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n612), .A2(G71gat), .A3(G78gat), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n600), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n595), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT102), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT19), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n617), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G127gat), .B(G155gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n615), .A2(new_n616), .ZN(new_n624));
  XOR2_X1   g423(.A(G183gat), .B(G211gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n623), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n590), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n531), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n548), .A2(new_n595), .A3(new_n565), .ZN(new_n632));
  INV_X1    g431(.A(new_n595), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n571), .ZN(new_n634));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT18), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n633), .B(new_n571), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n635), .B(KEYINPUT13), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n637), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G113gat), .B(G141gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G197gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT11), .ZN(new_n646));
  INV_X1    g445(.A(G169gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n638), .A2(new_n649), .A3(new_n642), .A4(new_n641), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n563), .A2(new_n615), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n557), .B(KEYINPUT108), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n558), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n561), .A2(new_n659), .A3(new_n614), .A4(new_n608), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n615), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n662), .A2(KEYINPUT10), .A3(new_n561), .A4(new_n562), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n655), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n656), .A2(new_n660), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n655), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT109), .ZN(new_n670));
  INV_X1    g469(.A(G176gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G204gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n665), .A2(new_n667), .A3(new_n673), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n653), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n631), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n456), .A2(new_n458), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  INV_X1    g482(.A(new_n452), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT42), .B1(new_n685), .B2(KEYINPUT110), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n688), .ZN(new_n690));
  OAI21_X1  g489(.A(G8gat), .B1(new_n679), .B2(new_n684), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT111), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n689), .B(new_n690), .C1(new_n693), .C2(new_n694), .ZN(G1325gat));
  XNOR2_X1  g494(.A(new_n522), .B(KEYINPUT112), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n680), .A2(G15gat), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(G15gat), .B1(new_n680), .B2(new_n523), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n679), .A2(new_n524), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  NAND2_X1  g502(.A1(new_n528), .A2(new_n530), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n443), .A2(new_n452), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n394), .A2(new_n395), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n405), .A2(KEYINPUT38), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n705), .B(new_n524), .C1(new_n525), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n463), .A2(new_n423), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n522), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n590), .B1(new_n704), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n629), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n678), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n540), .A3(new_n681), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT45), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n678), .A2(new_n713), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n531), .B2(new_n590), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n711), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  INV_X1    g520(.A(new_n590), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n718), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n681), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n717), .A2(new_n727), .ZN(G1328gat));
  NOR3_X1   g527(.A1(new_n714), .A2(G36gat), .A3(new_n684), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT46), .ZN(new_n730));
  OAI21_X1  g529(.A(G36gat), .B1(new_n725), .B2(new_n684), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1329gat));
  OAI21_X1  g531(.A(new_n534), .B1(new_n725), .B2(new_n522), .ZN(new_n733));
  INV_X1    g532(.A(new_n534), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n715), .A2(new_n734), .A3(new_n523), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n534), .B1(new_n725), .B2(new_n696), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(new_n735), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g538(.A(G50gat), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n724), .B2(new_n423), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n714), .A2(G50gat), .A3(new_n524), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT113), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g543(.A(new_n677), .ZN(new_n745));
  INV_X1    g544(.A(new_n653), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n630), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT114), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n720), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n681), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n684), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  AND2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n753), .B2(new_n754), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n749), .B2(new_n696), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n523), .A2(new_n487), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n749), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1334gat));
  NOR2_X1   g561(.A1(new_n749), .A2(new_n524), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT115), .B(G78gat), .Z(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n746), .A2(new_n629), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n677), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n719), .B2(new_n723), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n726), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n712), .A2(new_n766), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n677), .A2(new_n681), .A3(new_n554), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT116), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n770), .B1(new_n776), .B2(new_n778), .ZN(G1336gat));
  NOR2_X1   g578(.A1(new_n684), .A2(G92gat), .ZN(new_n780));
  AND4_X1   g579(.A1(KEYINPUT51), .A2(new_n720), .A3(new_n722), .A4(new_n766), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n712), .B2(new_n766), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n677), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n391), .B1(new_n768), .B2(new_n452), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT118), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n768), .A2(new_n452), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G92gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n789), .A2(new_n790), .A3(new_n784), .A4(new_n783), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n783), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n775), .A2(KEYINPUT117), .A3(new_n677), .A4(new_n780), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n789), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n792), .A2(new_n797), .ZN(G1337gat));
  NOR3_X1   g597(.A1(new_n769), .A2(new_n489), .A3(new_n696), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n775), .A2(new_n677), .A3(new_n523), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(new_n489), .ZN(G1338gat));
  OAI211_X1 g600(.A(new_n677), .B(new_n423), .C1(new_n781), .C2(new_n782), .ZN(new_n802));
  INV_X1    g601(.A(G106gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n768), .B2(new_n423), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT119), .B1(new_n768), .B2(new_n423), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n804), .A2(new_n806), .B1(new_n807), .B2(new_n803), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI221_X1 g609(.A(KEYINPUT53), .B1(new_n807), .B2(new_n803), .C1(new_n804), .C2(new_n806), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1339gat));
  NOR2_X1   g611(.A1(new_n726), .A2(new_n452), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n661), .A2(new_n655), .A3(new_n663), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT54), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n664), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n661), .A2(new_n663), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n654), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n674), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n814), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n673), .B1(new_n664), .B2(new_n819), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n823), .B(KEYINPUT55), .C1(new_n664), .C2(new_n816), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n676), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n822), .A2(KEYINPUT120), .A3(new_n824), .A4(new_n676), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n653), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n639), .A2(new_n640), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n635), .B1(new_n632), .B2(new_n634), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n648), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n652), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n677), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n590), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n827), .A2(new_n828), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n722), .A3(new_n833), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n629), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n630), .A2(new_n677), .A3(new_n746), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n813), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n423), .B1(new_n517), .B2(new_n519), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n653), .ZN(new_n844));
  INV_X1    g643(.A(new_n529), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n746), .A2(new_n234), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(G1340gat));
  OAI21_X1  g647(.A(G120gat), .B1(new_n843), .B2(new_n745), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n677), .A2(new_n232), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT121), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(new_n846), .B2(new_n851), .ZN(G1341gat));
  NOR3_X1   g651(.A1(new_n843), .A2(new_n227), .A3(new_n713), .ZN(new_n853));
  INV_X1    g652(.A(new_n846), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n629), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n227), .B2(new_n855), .ZN(G1342gat));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n225), .A3(new_n722), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n843), .B2(new_n590), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n854), .A2(new_n860), .A3(new_n225), .A4(new_n722), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(G1343gat));
  NAND2_X1  g661(.A1(new_n696), .A2(new_n423), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n863), .A2(KEYINPUT123), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n840), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n863), .A2(KEYINPUT123), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n865), .A2(new_n204), .A3(new_n746), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n653), .B1(new_n825), .B2(KEYINPUT122), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n822), .A2(new_n869), .A3(new_n824), .A4(new_n676), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n834), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n837), .B1(new_n871), .B2(new_n722), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n839), .B1(new_n872), .B2(new_n713), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT57), .B1(new_n873), .B2(new_n524), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n875), .B(new_n423), .C1(new_n838), .C2(new_n839), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n522), .A2(new_n813), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n874), .A2(new_n746), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G141gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT58), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1344gat));
  AND2_X1   g683(.A1(new_n865), .A2(new_n866), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n220), .A3(new_n677), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n871), .A2(new_n722), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n722), .A2(new_n833), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(new_n825), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n629), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n875), .B(new_n423), .C1(new_n891), .C2(new_n839), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n423), .B1(new_n838), .B2(new_n839), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n892), .A2(new_n894), .A3(new_n677), .A4(new_n877), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n887), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n874), .A2(new_n677), .A3(new_n876), .A4(new_n877), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n897), .A2(new_n887), .A3(G148gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n886), .B1(new_n896), .B2(new_n898), .ZN(G1345gat));
  NAND4_X1  g698(.A1(new_n865), .A2(new_n213), .A3(new_n629), .A4(new_n866), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n874), .A2(new_n629), .A3(new_n876), .A4(new_n877), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G155gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n900), .B2(new_n902), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  NAND3_X1  g705(.A1(new_n885), .A2(new_n214), .A3(new_n722), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n908));
  OAI21_X1  g707(.A(G162gat), .B1(new_n908), .B2(new_n590), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n684), .A2(new_n681), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n842), .B(new_n911), .C1(new_n838), .C2(new_n839), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n653), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n845), .B(new_n911), .C1(new_n838), .C2(new_n839), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n746), .A2(new_n647), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(G1348gat));
  NOR3_X1   g715(.A1(new_n912), .A2(new_n671), .A3(new_n745), .ZN(new_n917));
  INV_X1    g716(.A(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n677), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n671), .B2(new_n919), .ZN(G1349gat));
  INV_X1    g719(.A(new_n911), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n835), .A2(new_n837), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n713), .ZN(new_n923));
  INV_X1    g722(.A(new_n839), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n925), .A2(KEYINPUT125), .A3(new_n842), .A4(new_n629), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n912), .B2(new_n713), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(G183gat), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n629), .A2(new_n327), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n918), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT60), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n929), .A2(new_n935), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n912), .B2(new_n590), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT61), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n918), .A2(new_n322), .A3(new_n722), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n653), .A2(G197gat), .ZN(new_n942));
  INV_X1    g741(.A(new_n893), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n697), .A2(new_n921), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n943), .A2(KEYINPUT127), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT127), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n892), .A2(new_n894), .ZN(new_n948));
  INV_X1    g747(.A(new_n944), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n948), .A2(new_n653), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(G197gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  NOR2_X1   g751(.A1(new_n949), .A2(new_n893), .ZN(new_n953));
  INV_X1    g752(.A(G204gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n954), .A3(new_n677), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n953), .A2(new_n957), .A3(new_n954), .A4(new_n677), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n948), .A2(new_n745), .A3(new_n949), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n956), .B(new_n958), .C1(new_n959), .C2(new_n954), .ZN(G1353gat));
  OAI211_X1 g759(.A(new_n300), .B(new_n629), .C1(new_n945), .C2(new_n946), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n892), .A2(new_n894), .A3(new_n629), .A4(new_n944), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  NOR4_X1   g764(.A1(new_n948), .A2(new_n301), .A3(new_n590), .A4(new_n949), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n722), .B1(new_n945), .B2(new_n946), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n301), .ZN(G1355gat));
endmodule


