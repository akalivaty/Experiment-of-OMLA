

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  NOR2_X1 U321 ( .A1(n526), .A2(n447), .ZN(n561) );
  XOR2_X1 U322 ( .A(n402), .B(n401), .Z(n515) );
  XOR2_X1 U323 ( .A(G64GAT), .B(G204GAT), .Z(n289) );
  XOR2_X1 U324 ( .A(n339), .B(n443), .Z(n290) );
  INV_X1 U325 ( .A(KEYINPUT98), .ZN(n395) );
  XNOR2_X1 U326 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U327 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U328 ( .A(n343), .B(n342), .Z(n570) );
  INV_X1 U329 ( .A(G190GAT), .ZN(n448) );
  XNOR2_X1 U330 ( .A(KEYINPUT107), .B(n472), .ZN(n496) );
  XNOR2_X1 U331 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U332 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n475) );
  XNOR2_X1 U333 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XNOR2_X1 U334 ( .A(n476), .B(n475), .ZN(G1330GAT) );
  XNOR2_X1 U335 ( .A(G127GAT), .B(KEYINPUT81), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n291), .B(KEYINPUT0), .ZN(n292) );
  XOR2_X1 U337 ( .A(n292), .B(KEYINPUT82), .Z(n294) );
  XNOR2_X1 U338 ( .A(G113GAT), .B(G134GAT), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n421) );
  XOR2_X1 U340 ( .A(KEYINPUT86), .B(G176GAT), .Z(n296) );
  XNOR2_X1 U341 ( .A(G15GAT), .B(G190GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U343 ( .A(n297), .B(G99GAT), .Z(n299) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G71GAT), .Z(n340) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(n340), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U347 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n301) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U350 ( .A(n303), .B(n302), .Z(n309) );
  XNOR2_X1 U351 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n304), .B(KEYINPUT17), .ZN(n305) );
  XOR2_X1 U353 ( .A(n305), .B(G183GAT), .Z(n307) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(KEYINPUT85), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n400) );
  XNOR2_X1 U356 ( .A(n400), .B(KEYINPUT20), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n421), .B(n310), .ZN(n526) );
  XOR2_X1 U359 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n312) );
  XNOR2_X1 U360 ( .A(G211GAT), .B(KEYINPUT79), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n328) );
  XOR2_X1 U362 ( .A(G22GAT), .B(G155GAT), .Z(n427) );
  XOR2_X1 U363 ( .A(G78GAT), .B(G64GAT), .Z(n314) );
  XNOR2_X1 U364 ( .A(G127GAT), .B(G71GAT), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U366 ( .A(n427), .B(n315), .Z(n317) );
  NAND2_X1 U367 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U369 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n319) );
  XNOR2_X1 U370 ( .A(G183GAT), .B(KEYINPUT15), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U372 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U373 ( .A(G8GAT), .B(G15GAT), .Z(n323) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(KEYINPUT68), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n346) );
  XNOR2_X1 U376 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n324), .B(KEYINPUT13), .ZN(n335) );
  XNOR2_X1 U378 ( .A(n346), .B(n335), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n574) );
  XNOR2_X1 U381 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n361) );
  XOR2_X1 U382 ( .A(KEYINPUT71), .B(KEYINPUT73), .Z(n330) );
  XNOR2_X1 U383 ( .A(KEYINPUT32), .B(KEYINPUT70), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n343) );
  XOR2_X1 U385 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n332) );
  NAND2_X1 U386 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U388 ( .A(n333), .B(KEYINPUT31), .Z(n337) );
  XNOR2_X1 U389 ( .A(G176GAT), .B(G92GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n289), .B(n334), .ZN(n391) );
  XNOR2_X1 U391 ( .A(n335), .B(n391), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U393 ( .A(G148GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n338), .B(G78GAT), .ZN(n443) );
  XOR2_X1 U395 ( .A(G99GAT), .B(G85GAT), .Z(n375) );
  XNOR2_X1 U396 ( .A(n340), .B(n375), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n290), .B(n341), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n570), .B(KEYINPUT41), .ZN(n546) );
  XOR2_X1 U399 ( .A(G29GAT), .B(G43GAT), .Z(n345) );
  XNOR2_X1 U400 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n367) );
  XNOR2_X1 U402 ( .A(n367), .B(n346), .ZN(n359) );
  XOR2_X1 U403 ( .A(KEYINPUT66), .B(G22GAT), .Z(n348) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U406 ( .A(n349), .B(KEYINPUT67), .Z(n357) );
  XOR2_X1 U407 ( .A(G141GAT), .B(G113GAT), .Z(n351) );
  XNOR2_X1 U408 ( .A(G50GAT), .B(G36GAT), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U410 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n353) );
  XNOR2_X1 U411 ( .A(G169GAT), .B(G197GAT), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n566) );
  NAND2_X1 U416 ( .A1(n546), .A2(n566), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  NOR2_X1 U418 ( .A1(n574), .A2(n362), .ZN(n380) );
  XOR2_X1 U419 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n364) );
  XNOR2_X1 U420 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n379) );
  XOR2_X1 U422 ( .A(KEYINPUT75), .B(G218GAT), .Z(n366) );
  XOR2_X1 U423 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XOR2_X1 U424 ( .A(G36GAT), .B(G190GAT), .Z(n394) );
  XNOR2_X1 U425 ( .A(n428), .B(n394), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U427 ( .A(G134GAT), .B(n367), .Z(n369) );
  NAND2_X1 U428 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U430 ( .A(n371), .B(n370), .Z(n377) );
  XOR2_X1 U431 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n373) );
  XNOR2_X1 U432 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n477) );
  NAND2_X1 U437 ( .A1(n380), .A2(n477), .ZN(n381) );
  XNOR2_X1 U438 ( .A(KEYINPUT47), .B(n381), .ZN(n387) );
  XOR2_X1 U439 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n383) );
  INV_X1 U440 ( .A(n477), .ZN(n551) );
  XNOR2_X1 U441 ( .A(KEYINPUT36), .B(n551), .ZN(n576) );
  NAND2_X1 U442 ( .A1(n574), .A2(n576), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n384) );
  NAND2_X1 U444 ( .A1(n384), .A2(n570), .ZN(n385) );
  NOR2_X1 U445 ( .A1(n566), .A2(n385), .ZN(n386) );
  NOR2_X1 U446 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U447 ( .A(KEYINPUT48), .B(n388), .ZN(n524) );
  XOR2_X1 U448 ( .A(KEYINPUT21), .B(G211GAT), .Z(n390) );
  XNOR2_X1 U449 ( .A(G197GAT), .B(G218GAT), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n442) );
  XOR2_X1 U451 ( .A(n391), .B(KEYINPUT97), .Z(n393) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n398) );
  XNOR2_X1 U454 ( .A(G8GAT), .B(n394), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n442), .B(n399), .ZN(n402) );
  INV_X1 U456 ( .A(n400), .ZN(n401) );
  INV_X1 U457 ( .A(n515), .ZN(n453) );
  NOR2_X1 U458 ( .A1(n524), .A2(n453), .ZN(n404) );
  INV_X1 U459 ( .A(KEYINPUT54), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n426) );
  XOR2_X1 U461 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n406) );
  XNOR2_X1 U462 ( .A(KEYINPUT1), .B(KEYINPUT93), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U464 ( .A(G57GAT), .B(G162GAT), .Z(n408) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(G85GAT), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n425) );
  XOR2_X1 U468 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n412) );
  XNOR2_X1 U469 ( .A(KEYINPUT92), .B(KEYINPUT95), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U471 ( .A(G148GAT), .B(KEYINPUT5), .Z(n414) );
  XNOR2_X1 U472 ( .A(G120GAT), .B(G155GAT), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U474 ( .A(n416), .B(n415), .Z(n423) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n417), .B(KEYINPUT2), .ZN(n432) );
  XOR2_X1 U477 ( .A(n432), .B(G1GAT), .Z(n419) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n513) );
  NOR2_X1 U483 ( .A1(n426), .A2(n513), .ZN(n565) );
  XOR2_X1 U484 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n430) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U487 ( .A(n431), .B(KEYINPUT89), .Z(n437) );
  XOR2_X1 U488 ( .A(KEYINPUT88), .B(n432), .Z(n434) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U491 ( .A(G204GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U493 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n439) );
  XNOR2_X1 U494 ( .A(KEYINPUT22), .B(KEYINPUT90), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U496 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n461) );
  AND2_X1 U499 ( .A1(n565), .A2(n461), .ZN(n446) );
  XNOR2_X1 U500 ( .A(KEYINPUT55), .B(n446), .ZN(n447) );
  NAND2_X1 U501 ( .A1(n561), .A2(n551), .ZN(n451) );
  XOR2_X1 U502 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n449) );
  XOR2_X1 U503 ( .A(KEYINPUT37), .B(KEYINPUT106), .Z(n470) );
  INV_X1 U504 ( .A(n526), .ZN(n517) );
  XNOR2_X1 U505 ( .A(n461), .B(KEYINPUT65), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n452), .B(KEYINPUT28), .ZN(n529) );
  XOR2_X1 U507 ( .A(KEYINPUT27), .B(n453), .Z(n458) );
  NAND2_X1 U508 ( .A1(n513), .A2(n458), .ZN(n523) );
  NOR2_X1 U509 ( .A1(n529), .A2(n523), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n454), .B(KEYINPUT99), .ZN(n455) );
  NOR2_X1 U511 ( .A1(n517), .A2(n455), .ZN(n467) );
  XNOR2_X1 U512 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n457) );
  NOR2_X1 U513 ( .A1(n517), .A2(n461), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n564) );
  NAND2_X1 U515 ( .A1(n564), .A2(n458), .ZN(n459) );
  XNOR2_X1 U516 ( .A(KEYINPUT101), .B(n459), .ZN(n464) );
  NAND2_X1 U517 ( .A1(n517), .A2(n515), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U519 ( .A(KEYINPUT25), .B(n462), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n513), .A2(n465), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n479) );
  NOR2_X1 U523 ( .A1(n479), .A2(n574), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n468), .A2(n576), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n470), .B(n469), .ZN(n512) );
  NAND2_X1 U526 ( .A1(n566), .A2(n570), .ZN(n482) );
  NOR2_X1 U527 ( .A1(n512), .A2(n482), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT38), .B(n471), .Z(n472) );
  NAND2_X1 U529 ( .A1(n496), .A2(n515), .ZN(n474) );
  XNOR2_X1 U530 ( .A(G36GAT), .B(KEYINPUT108), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n474), .B(n473), .ZN(G1329GAT) );
  NAND2_X1 U532 ( .A1(n496), .A2(n517), .ZN(n476) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n485) );
  NAND2_X1 U534 ( .A1(n477), .A2(n574), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(n478), .Z(n481) );
  INV_X1 U536 ( .A(n479), .ZN(n480) );
  NAND2_X1 U537 ( .A1(n481), .A2(n480), .ZN(n499) );
  NOR2_X1 U538 ( .A1(n482), .A2(n499), .ZN(n483) );
  XNOR2_X1 U539 ( .A(KEYINPUT102), .B(n483), .ZN(n491) );
  NAND2_X1 U540 ( .A1(n513), .A2(n491), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  XOR2_X1 U542 ( .A(G8GAT), .B(KEYINPUT103), .Z(n487) );
  NAND2_X1 U543 ( .A1(n515), .A2(n491), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U546 ( .A1(n517), .A2(n491), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(n490), .ZN(G1326GAT) );
  XOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT105), .Z(n493) );
  NAND2_X1 U550 ( .A1(n529), .A2(n491), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(G1327GAT) );
  XOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U553 ( .A1(n513), .A2(n496), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n496), .A2(n529), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n497), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U557 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n501) );
  INV_X1 U558 ( .A(n566), .ZN(n498) );
  XOR2_X1 U559 ( .A(KEYINPUT109), .B(n546), .Z(n558) );
  NAND2_X1 U560 ( .A1(n498), .A2(n558), .ZN(n511) );
  NOR2_X1 U561 ( .A1(n499), .A2(n511), .ZN(n506) );
  NAND2_X1 U562 ( .A1(n513), .A2(n506), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1332GAT) );
  NAND2_X1 U564 ( .A1(n506), .A2(n515), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n504) );
  NAND2_X1 U567 ( .A1(n506), .A2(n517), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U569 ( .A(G71GAT), .B(n505), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U571 ( .A1(n506), .A2(n529), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n510) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT113), .Z(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NOR2_X1 U575 ( .A1(n512), .A2(n511), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n513), .A2(n519), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n519), .A2(n515), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U580 ( .A1(n519), .A2(n517), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n521) );
  NAND2_X1 U583 ( .A1(n519), .A2(n529), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(G106GAT), .B(n522), .Z(G1339GAT) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(KEYINPUT118), .ZN(n531) );
  NOR2_X1 U587 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U588 ( .A(KEYINPUT116), .B(n525), .Z(n544) );
  NOR2_X1 U589 ( .A1(n544), .A2(n526), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(KEYINPUT117), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n566), .A2(n539), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U595 ( .A1(n539), .A2(n558), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U597 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(KEYINPUT121), .ZN(n538) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n536) );
  NAND2_X1 U600 ( .A1(n539), .A2(n574), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U604 ( .A1(n539), .A2(n551), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  INV_X1 U607 ( .A(n564), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n566), .A2(n552), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U612 ( .A1(n552), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n574), .A2(n552), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n566), .A2(n561), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n556) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(n557), .Z(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT125), .Z(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n574), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  AND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n577) );
  NAND2_X1 U632 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  INV_X1 U636 ( .A(n570), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n577), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n577), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

