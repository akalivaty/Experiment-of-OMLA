//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287;
  OR3_X1    g0000(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n201));
  OAI21_X1  g0001(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(KEYINPUT65), .B(G50), .ZN(new_n205));
  AND3_X1   g0005(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT66), .Z(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n203), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n212), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT67), .Z(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT68), .Z(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n218), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT69), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT70), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  AND2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G222), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n254), .B1(new_n204), .B2(new_n252), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n258), .A2(new_n262), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(G226), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G200), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n213), .ZN(new_n271));
  XOR2_X1   g0071(.A(KEYINPUT8), .B(G58), .Z(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n214), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n214), .B1(new_n203), .B2(new_n205), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n271), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G13), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G1), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(G1), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n271), .B1(new_n285), .B2(G20), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(G50), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT9), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n259), .A2(G190), .A3(new_n267), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n280), .A2(KEYINPUT9), .A3(new_n287), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n269), .A2(new_n290), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n294), .A2(KEYINPUT72), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n296), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(KEYINPUT72), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n268), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n288), .C1(G179), .C2(new_n268), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n283), .A2(G77), .ZN(new_n306));
  INV_X1    g0106(.A(new_n271), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT15), .B(G87), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n274), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n309), .A2(new_n310), .B1(G20), .B2(G77), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n272), .A2(new_n276), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n307), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI211_X1 g0113(.A(new_n306), .B(new_n313), .C1(G77), .C2(new_n286), .ZN(new_n314));
  INV_X1    g0114(.A(G238), .ZN(new_n315));
  INV_X1    g0115(.A(G107), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n255), .A2(new_n315), .B1(new_n316), .B2(new_n252), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n249), .A2(new_n251), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n318), .A2(new_n232), .A3(G1698), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n258), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n265), .B1(new_n266), .B2(G244), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n314), .B1(new_n322), .B2(new_n303), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(G200), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n314), .B(new_n327), .C1(new_n328), .C2(new_n322), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n302), .A2(new_n305), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT73), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n282), .ZN(new_n334));
  INV_X1    g0134(.A(G68), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G20), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT75), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  XOR2_X1   g0137(.A(new_n337), .B(KEYINPUT12), .Z(new_n338));
  NAND2_X1  g0138(.A1(new_n286), .A2(G68), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT76), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n336), .B1(new_n274), .B2(new_n204), .C1(new_n277), .C2(new_n216), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n271), .ZN(new_n343));
  XOR2_X1   g0143(.A(new_n343), .B(KEYINPUT11), .Z(new_n344));
  NOR2_X1   g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n265), .ZN(new_n346));
  INV_X1    g0146(.A(new_n266), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n315), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n252), .A2(G226), .A3(new_n253), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n348), .B1(new_n352), .B2(new_n258), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n353), .A2(new_n354), .ZN(new_n357));
  OAI21_X1  g0157(.A(G200), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n355), .B(G190), .C1(new_n359), .C2(new_n353), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n345), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(G169), .B1(new_n356), .B2(new_n357), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT14), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(G169), .C1(new_n356), .C2(new_n357), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n355), .B(G179), .C1(new_n359), .C2(new_n353), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n345), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n333), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n273), .B1(new_n285), .B2(G20), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n281), .A2(new_n214), .A3(G1), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n271), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n371), .A2(new_n373), .B1(new_n372), .B2(new_n273), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G58), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n335), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n203), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n276), .A2(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT77), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT77), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n250), .A3(G33), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n383), .A3(new_n249), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n214), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G68), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n384), .B2(new_n214), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT78), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n384), .A2(new_n214), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT7), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT78), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(G68), .A4(new_n386), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n380), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n307), .B1(new_n394), .B2(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT7), .B1(new_n252), .B2(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n318), .A2(new_n385), .A3(new_n214), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n397), .A2(G68), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n396), .B1(new_n399), .B2(new_n380), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n375), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(G226), .A2(G1698), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n381), .A2(new_n383), .A3(new_n249), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT79), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n381), .A2(new_n383), .A3(new_n253), .A4(new_n249), .ZN(new_n406));
  INV_X1    g0206(.A(G87), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n406), .A2(new_n256), .B1(new_n248), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n258), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n265), .B1(new_n266), .B2(G232), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n303), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n410), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n403), .B(KEYINPUT79), .ZN(new_n413));
  INV_X1    g0213(.A(new_n408), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(new_n415), .B2(new_n258), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n411), .B1(G179), .B2(new_n416), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n401), .A2(KEYINPUT18), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n389), .A2(new_n393), .ZN(new_n420));
  INV_X1    g0220(.A(new_n380), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(KEYINPUT16), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(new_n400), .A3(new_n271), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n374), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n416), .A2(G179), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n303), .B2(new_n416), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n419), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT80), .B1(new_n418), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT81), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n409), .A2(new_n328), .A3(new_n410), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n416), .B2(G200), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n429), .B1(new_n401), .B2(new_n431), .ZN(new_n432));
  AND4_X1   g0232(.A1(new_n429), .A2(new_n423), .A3(new_n374), .A4(new_n431), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT17), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT17), .B1(new_n401), .B2(new_n431), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT18), .B1(new_n401), .B2(new_n417), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n424), .A2(new_n419), .A3(new_n426), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT80), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n428), .A2(new_n434), .A3(new_n436), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n331), .A2(new_n332), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n370), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(G1), .B(G13), .C1(new_n248), .C2(new_n260), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n383), .A2(new_n249), .ZN(new_n445));
  NOR2_X1   g0245(.A1(G257), .A2(G1698), .ZN(new_n446));
  INV_X1    g0246(.A(G264), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(G1698), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n381), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n318), .A2(G303), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n444), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n285), .A2(G45), .ZN(new_n452));
  OR2_X1    g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(G274), .A3(new_n444), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT5), .B(G41), .ZN(new_n457));
  INV_X1    g0257(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n444), .ZN(new_n460));
  INV_X1    g0260(.A(G270), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT83), .B1(new_n451), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n455), .A2(new_n258), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n258), .A2(new_n264), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n464), .A2(G270), .B1(new_n465), .B2(new_n455), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n447), .A2(G1698), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(G257), .B2(G1698), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n450), .B1(new_n384), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n258), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT83), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  INV_X1    g0273(.A(G97), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n473), .B(new_n214), .C1(G33), .C2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G20), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n271), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT20), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n475), .A2(KEYINPUT20), .A3(new_n271), .A4(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n283), .A2(G116), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n248), .A2(G1), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n372), .A2(new_n271), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(G116), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n303), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n463), .A2(KEYINPUT21), .A3(new_n472), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n486), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(G179), .A3(new_n470), .A4(new_n466), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n463), .A2(new_n472), .A3(new_n487), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n491), .A2(KEYINPUT84), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n488), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n489), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n463), .A2(G200), .A3(new_n472), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n463), .A2(new_n472), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n498), .C1(new_n499), .C2(new_n328), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n494), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n316), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n474), .A2(new_n316), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n502), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n397), .A2(G107), .A3(new_n398), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n307), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n485), .A2(G97), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(G97), .B2(new_n283), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n464), .A2(G257), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n456), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n318), .A2(new_n253), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT4), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n381), .A2(new_n383), .A3(G244), .A4(new_n249), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(G1698), .ZN(new_n520));
  AND2_X1   g0320(.A1(KEYINPUT4), .A2(G244), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n249), .A2(new_n251), .A3(new_n521), .A4(new_n253), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT82), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n522), .A2(KEYINPUT82), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n517), .A2(new_n520), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n515), .B1(new_n525), .B2(new_n258), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n324), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n513), .B(new_n527), .C1(G169), .C2(new_n526), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n381), .A2(new_n383), .A3(new_n214), .A4(new_n249), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT22), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n529), .A2(new_n530), .A3(new_n407), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n214), .A2(G87), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n318), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G20), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n214), .B2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n316), .A2(KEYINPUT23), .A3(G20), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  OR3_X1    g0340(.A1(new_n531), .A2(new_n540), .A3(KEYINPUT24), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT24), .B1(new_n531), .B2(new_n540), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n307), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n485), .A2(G107), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT25), .B1(new_n372), .B2(new_n316), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n372), .A2(KEYINPUT25), .A3(new_n316), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G257), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G1698), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(G250), .B2(G1698), .ZN(new_n551));
  INV_X1    g0351(.A(G294), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n384), .A2(new_n551), .B1(new_n248), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n258), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n464), .A2(G264), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n456), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n328), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(G200), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n526), .A2(G190), .ZN(new_n560));
  INV_X1    g0360(.A(G200), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n512), .C1(new_n561), .C2(new_n526), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n528), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n554), .A2(new_n555), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n324), .A3(new_n456), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n556), .A2(new_n303), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n565), .B(new_n566), .C1(new_n543), .C2(new_n547), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n452), .A2(G250), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n444), .B1(G274), .B2(new_n458), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n445), .A2(G238), .A3(new_n253), .A4(new_n381), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n445), .A2(G244), .A3(G1698), .A4(new_n381), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(new_n534), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n570), .B1(new_n573), .B2(new_n258), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n324), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n529), .A2(new_n335), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  AND4_X1   g0377(.A1(new_n577), .A2(new_n214), .A3(G33), .A4(G97), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n407), .A2(new_n474), .A3(new_n316), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n351), .A2(new_n214), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n578), .B1(new_n581), .B2(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n271), .B1(new_n576), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n308), .A2(new_n372), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n485), .A2(new_n309), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n575), .B(new_n586), .C1(new_n574), .C2(G169), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n485), .A2(G87), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n583), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n574), .B2(G190), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n534), .B1(new_n519), .B2(new_n253), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n406), .A2(new_n315), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n258), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n569), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n567), .A2(new_n587), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n563), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n443), .A2(new_n501), .A3(new_n598), .ZN(G372));
  INV_X1    g0399(.A(KEYINPUT85), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(KEYINPUT85), .B(new_n258), .C1(new_n591), .C2(new_n592), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n570), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n575), .B(new_n586), .C1(new_n603), .C2(G169), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n590), .B1(new_n603), .B2(new_n561), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT86), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT86), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT26), .ZN(new_n611));
  INV_X1    g0411(.A(new_n528), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n563), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n493), .A2(new_n492), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n567), .A2(new_n488), .A3(new_n615), .A4(new_n490), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n604), .ZN(new_n618));
  INV_X1    g0418(.A(new_n526), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n512), .B1(new_n619), .B2(new_n303), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n620), .A2(new_n587), .A3(new_n596), .A4(new_n527), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n621), .B2(KEYINPUT26), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n613), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n443), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n434), .A2(new_n436), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n367), .A2(new_n368), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n345), .A2(new_n358), .A3(new_n360), .ZN(new_n627));
  INV_X1    g0427(.A(new_n326), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n625), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT87), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n418), .B2(new_n427), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT87), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n302), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n305), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n624), .A2(new_n637), .ZN(G369));
  OR3_X1    g0438(.A1(new_n334), .A2(KEYINPUT27), .A3(G20), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT27), .B1(new_n334), .B2(G20), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n489), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n501), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n644), .ZN(new_n647));
  XOR2_X1   g0447(.A(KEYINPUT88), .B(G330), .Z(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n567), .A2(new_n643), .ZN(new_n651));
  INV_X1    g0451(.A(new_n643), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n559), .B1(new_n548), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n651), .B1(new_n653), .B2(new_n567), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n643), .B1(new_n494), .B2(new_n496), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(G399));
  INV_X1    g0458(.A(new_n209), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n579), .A2(G116), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G1), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n217), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n661), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT29), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n604), .B1(new_n621), .B2(KEYINPUT26), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n608), .B1(new_n604), .B2(new_n605), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n612), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n668), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n491), .A2(KEYINPUT84), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n496), .A3(new_n567), .A4(new_n615), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT93), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT93), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n494), .A2(new_n676), .A3(new_n496), .A4(new_n567), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n610), .A2(new_n675), .A3(new_n614), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n652), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT94), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT94), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n679), .A2(new_n682), .A3(new_n652), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n667), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n623), .A2(new_n652), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT95), .B1(new_n685), .B2(KEYINPUT29), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n598), .A2(new_n501), .A3(new_n652), .ZN(new_n688));
  OR2_X1    g0488(.A1(KEYINPUT91), .A2(KEYINPUT30), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n526), .A2(new_n564), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT91), .B1(KEYINPUT90), .B2(KEYINPUT30), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT89), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n466), .A2(new_n470), .A3(new_n694), .A4(G179), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n466), .A2(new_n470), .A3(G179), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n594), .B1(KEYINPUT89), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n691), .A2(new_n693), .A3(new_n695), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(KEYINPUT89), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n574), .A3(new_n695), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n692), .B1(new_n690), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n603), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n556), .A2(new_n324), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n499), .A3(new_n619), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n698), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n643), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n688), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n648), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT92), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n713), .A3(new_n648), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT95), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n682), .B1(new_n679), .B2(new_n652), .ZN(new_n718));
  AOI211_X1 g0518(.A(KEYINPUT94), .B(new_n643), .C1(new_n672), .C2(new_n678), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n717), .B(KEYINPUT29), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n687), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n666), .B1(new_n722), .B2(G1), .ZN(G364));
  NOR2_X1   g0523(.A1(new_n281), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n285), .B1(new_n724), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n660), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n650), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n648), .B2(new_n647), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n213), .B1(G20), .B2(new_n303), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n324), .A2(new_n561), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n214), .A2(G190), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G317), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT33), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(KEYINPUT33), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G329), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G179), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n739), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n214), .A2(new_n328), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n324), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n743), .B1(G322), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n214), .B1(new_n741), .B2(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G294), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n561), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n744), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G303), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n733), .A2(new_n745), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n732), .A2(new_n744), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n252), .B(new_n757), .C1(G326), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n733), .A2(new_n752), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT96), .Z(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G283), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n748), .A2(new_n751), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n252), .B1(new_n749), .B2(new_n474), .C1(new_n758), .C2(new_n216), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n734), .A2(new_n335), .B1(new_n755), .B2(new_n204), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n376), .A2(new_n746), .B1(new_n753), .B2(new_n407), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n762), .A2(G107), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n742), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n768), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n731), .B1(new_n764), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n730), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n217), .A2(new_n261), .ZN(new_n780));
  INV_X1    g0580(.A(new_n384), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n659), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n780), .B(new_n782), .C1(new_n246), .C2(new_n261), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n659), .A2(new_n318), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G355), .B1(new_n476), .B2(new_n659), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n779), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n727), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n774), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n777), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n647), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n729), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  NAND2_X1  g0592(.A1(new_n628), .A2(new_n652), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n329), .B1(new_n314), .B2(new_n652), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n326), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n685), .B(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n727), .B1(new_n799), .B2(new_n716), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n716), .B2(new_n799), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n762), .A2(G87), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n756), .B2(new_n742), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT98), .Z(new_n804));
  INV_X1    g0604(.A(new_n755), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n759), .A2(G303), .B1(new_n805), .B2(G116), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n316), .B2(new_n753), .C1(new_n807), .C2(new_n734), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n318), .B1(new_n749), .B2(new_n474), .C1(new_n552), .C2(new_n746), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G143), .A2(new_n747), .B1(new_n805), .B2(G159), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n811), .B1(new_n812), .B2(new_n758), .C1(new_n275), .C2(new_n734), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n762), .A2(G68), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n753), .A2(new_n216), .B1(new_n742), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n384), .B(new_n817), .C1(G58), .C2(new_n750), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n730), .B1(new_n810), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n731), .A2(new_n776), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT97), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n787), .B1(new_n823), .B2(new_n204), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n820), .B(new_n824), .C1(new_n798), .C2(new_n776), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n801), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G384));
  NOR2_X1   g0627(.A1(new_n724), .A2(new_n285), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n720), .B1(new_n684), .B2(new_n686), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n636), .B1(new_n829), .B2(new_n443), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT101), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT39), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n395), .B1(KEYINPUT16), .B2(new_n394), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n374), .ZN(new_n834));
  INV_X1    g0634(.A(new_n641), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n441), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n425), .B(new_n641), .C1(new_n303), .C2(new_n416), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n423), .A2(new_n374), .A3(new_n431), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT81), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n401), .A2(new_n429), .A3(new_n431), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n424), .A2(new_n839), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n842), .A2(new_n843), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n838), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n401), .A2(new_n641), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n634), .B2(new_n625), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n847), .A2(new_n841), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n848), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n832), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n367), .A2(new_n368), .A3(new_n652), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT100), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n437), .A2(new_n439), .A3(new_n438), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n439), .B1(new_n437), .B2(new_n438), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n435), .B1(new_n844), .B2(KEYINPUT17), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n836), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n845), .A2(new_n848), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n838), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n857), .A2(new_n859), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n345), .A2(new_n652), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n626), .A2(new_n627), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n367), .A2(new_n872), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n623), .A2(new_n652), .A3(new_n798), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n793), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n871), .A2(new_n879), .B1(new_n634), .B2(new_n641), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n870), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n831), .B(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n876), .A2(new_n710), .A3(new_n798), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n838), .B2(new_n849), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n850), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  INV_X1    g0688(.A(new_n851), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n437), .A2(KEYINPUT87), .A3(new_n438), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT87), .B1(new_n437), .B2(new_n438), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n889), .B1(new_n892), .B2(new_n864), .ZN(new_n893));
  INV_X1    g0693(.A(new_n855), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n860), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n868), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n884), .A2(new_n888), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n887), .A2(new_n888), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n443), .A2(new_n710), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n648), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n828), .B1(new_n883), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n883), .B2(new_n902), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n664), .A2(new_n204), .A3(new_n377), .ZN(new_n905));
  INV_X1    g0705(.A(new_n205), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n335), .ZN(new_n907));
  OAI211_X1 g0707(.A(G1), .B(new_n281), .C1(new_n905), .C2(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n506), .A2(KEYINPUT35), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n506), .A2(KEYINPUT35), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(G116), .A3(new_n215), .A4(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n904), .A2(new_n908), .A3(new_n913), .ZN(G367));
  INV_X1    g0714(.A(new_n782), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n778), .B1(new_n209), .B2(new_n308), .C1(new_n915), .C2(new_n238), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n753), .A2(new_n376), .B1(new_n761), .B2(new_n204), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n742), .A2(new_n812), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(G143), .B2(new_n759), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n252), .C1(new_n275), .C2(new_n746), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n734), .A2(new_n770), .B1(new_n755), .B2(new_n205), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n749), .A2(new_n335), .ZN(new_n922));
  OR4_X1    g0722(.A1(new_n917), .A2(new_n920), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n753), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(G116), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT46), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n758), .A2(new_n756), .B1(new_n746), .B2(new_n754), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT107), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n734), .A2(new_n552), .B1(new_n761), .B2(new_n474), .ZN(new_n932));
  XNOR2_X1  g0732(.A(KEYINPUT108), .B(G317), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n755), .A2(new_n807), .B1(new_n742), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n384), .C1(new_n316), .C2(new_n749), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n923), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT47), .Z(new_n938));
  OAI211_X1 g0738(.A(new_n727), .B(new_n916), .C1(new_n938), .C2(new_n731), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n589), .A2(new_n643), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n604), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n610), .B2(new_n940), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n939), .B1(new_n942), .B2(new_n777), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n528), .B(new_n562), .C1(new_n512), .C2(new_n652), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n528), .B2(new_n652), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT102), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n654), .A3(new_n656), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT42), .Z(new_n949));
  OAI21_X1  g0749(.A(new_n528), .B1(new_n946), .B2(new_n567), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n652), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT43), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n942), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n942), .A2(new_n953), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n655), .A2(new_n946), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n956), .B2(new_n957), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n960), .B2(KEYINPUT103), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(KEYINPUT103), .B2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(new_n657), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n946), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT105), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT104), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n964), .B2(new_n965), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(KEYINPUT105), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n946), .A2(new_n963), .A3(KEYINPUT104), .A4(KEYINPUT44), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n967), .A2(new_n969), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n947), .A2(new_n657), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT45), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n650), .A2(KEYINPUT106), .A3(new_n654), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n975), .B(new_n976), .Z(new_n977));
  XNOR2_X1  g0777(.A(new_n654), .B(new_n656), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n649), .B(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n722), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(new_n721), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n660), .B(KEYINPUT41), .Z(new_n984));
  OAI21_X1  g0784(.A(new_n725), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n943), .B1(new_n962), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(G387));
  NAND2_X1  g0787(.A1(new_n721), .A2(new_n979), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n981), .A2(new_n660), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n979), .A2(new_n725), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT109), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT109), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n654), .A2(new_n789), .ZN(new_n994));
  INV_X1    g0794(.A(new_n662), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n784), .A2(new_n995), .B1(new_n316), .B2(new_n659), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT110), .Z(new_n997));
  OR2_X1    g0797(.A1(new_n235), .A2(new_n261), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n272), .A2(new_n216), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT50), .Z(new_n1000));
  AOI211_X1 g0800(.A(G45), .B(new_n995), .C1(G68), .C2(G77), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n915), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n997), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n753), .A2(new_n204), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G50), .B2(new_n747), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n750), .A2(new_n309), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n781), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n742), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n759), .A2(G159), .B1(new_n1008), .B2(G150), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n335), .B2(new_n755), .C1(new_n273), .C2(new_n734), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1007), .B(new_n1010), .C1(G97), .C2(new_n762), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n924), .A2(G294), .B1(new_n750), .B2(G283), .ZN(new_n1012));
  XOR2_X1   g0812(.A(KEYINPUT111), .B(G322), .Z(new_n1013));
  AOI22_X1  g0813(.A1(new_n759), .A2(new_n1013), .B1(new_n735), .B2(G311), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n754), .B2(new_n755), .C1(new_n746), .C2(new_n933), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT48), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n1016), .B2(new_n1015), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT49), .ZN(new_n1019));
  INV_X1    g0819(.A(G326), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n384), .B1(new_n742), .B2(new_n1020), .C1(new_n476), .C2(new_n761), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT112), .Z(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n1018), .B2(KEYINPUT49), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1011), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n727), .B1(new_n779), .B2(new_n1003), .C1(new_n1024), .C2(new_n731), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT113), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n992), .A2(new_n993), .B1(new_n994), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n989), .A2(new_n1027), .ZN(G393));
  AOI22_X1  g0828(.A1(G68), .A2(new_n924), .B1(new_n1008), .B2(G143), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n735), .A2(new_n906), .B1(new_n805), .B2(new_n272), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n384), .B1(G77), .B2(new_n750), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n802), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n758), .A2(new_n275), .B1(new_n746), .B2(new_n770), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT51), .Z(new_n1034));
  OAI22_X1  g0834(.A1(new_n758), .A2(new_n736), .B1(new_n746), .B2(new_n756), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT52), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n769), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G283), .A2(new_n924), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n252), .B1(new_n805), .B2(G294), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n735), .A2(G303), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n750), .A2(G116), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1032), .A2(new_n1034), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n730), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n243), .A2(new_n915), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n778), .B1(new_n474), .B2(new_n209), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1046), .B(new_n727), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n946), .B2(new_n777), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n975), .B(new_n655), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1050), .B1(new_n1051), .B2(new_n726), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n722), .B2(new_n980), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n660), .B1(new_n977), .B2(new_n981), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(G390));
  AND2_X1   g0855(.A1(new_n710), .A2(new_n798), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1056), .A2(G330), .A3(new_n876), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n859), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n850), .B2(new_n856), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n718), .A2(new_n719), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n797), .B1(new_n1061), .B2(new_n793), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n876), .B(KEYINPUT114), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n878), .A2(new_n793), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n859), .B1(new_n1065), .B2(new_n876), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n857), .B2(new_n869), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1058), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n850), .A2(new_n886), .A3(new_n832), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT39), .B1(new_n895), .B2(new_n868), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1069), .A2(new_n1070), .B1(new_n859), .B2(new_n879), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n710), .A2(new_n713), .A3(new_n648), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n713), .B1(new_n710), .B2(new_n648), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n798), .B(new_n876), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(KEYINPUT115), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT115), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n715), .A2(new_n1076), .A3(new_n798), .A4(new_n876), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n681), .A2(new_n683), .A3(new_n793), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n796), .A3(new_n1063), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n859), .B1(new_n895), .B2(new_n868), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1071), .A2(new_n1078), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1068), .A2(new_n1083), .A3(new_n726), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n775), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n727), .B1(new_n822), .B2(new_n272), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT117), .Z(new_n1087));
  OAI22_X1  g0887(.A1(new_n758), .A2(new_n807), .B1(new_n734), .B2(new_n316), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n252), .B(new_n1088), .C1(G87), .C2(new_n924), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n750), .A2(G77), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n755), .A2(new_n474), .B1(new_n742), .B2(new_n552), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G116), .B2(new_n747), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1089), .A2(new_n815), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n252), .B1(new_n746), .B2(new_n816), .ZN(new_n1094));
  INV_X1    g0894(.A(G128), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n758), .A2(new_n1095), .B1(new_n734), .B2(new_n812), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(G159), .C2(new_n750), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n753), .A2(new_n275), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT53), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n205), .A2(new_n761), .B1(new_n755), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G125), .B2(new_n1008), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1097), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1093), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1085), .B(new_n1087), .C1(new_n731), .C2(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1084), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n899), .A2(G330), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n830), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n876), .B(KEYINPUT114), .Z(new_n1109));
  NAND2_X1  g0909(.A1(new_n1056), .A2(G330), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(new_n1110), .B1(new_n1079), .B2(new_n796), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n798), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n712), .B2(new_n714), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1057), .B1(new_n1113), .B2(new_n876), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1078), .A2(new_n1111), .B1(new_n1114), .B2(new_n1065), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n1083), .A3(new_n1068), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1068), .A2(new_n1083), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n660), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT116), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1106), .B1(new_n1122), .B2(new_n1123), .ZN(G378));
  INV_X1    g0924(.A(KEYINPUT121), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n302), .A2(new_n305), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n288), .A2(new_n835), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n898), .B2(G330), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n897), .B1(new_n850), .B2(new_n856), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n884), .B1(new_n867), .B2(new_n868), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n1132), .C1(new_n1133), .C2(KEYINPUT40), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1130), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n881), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT119), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n881), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n898), .A2(G330), .A3(new_n1130), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1138), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1108), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n1118), .B2(new_n1115), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1140), .A2(new_n1139), .A3(new_n1141), .A4(KEYINPUT119), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT120), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT57), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1148), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1145), .A2(new_n1152), .A3(KEYINPUT57), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n660), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1150), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1143), .A2(new_n726), .A3(new_n1146), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n727), .B1(new_n821), .B2(new_n906), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n758), .A2(new_n1158), .B1(new_n734), .B2(new_n816), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n805), .A2(G137), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n1095), .B2(new_n746), .C1(new_n753), .C2(new_n1100), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1159), .B(new_n1161), .C1(G150), .C2(new_n750), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n733), .A2(new_n752), .A3(G159), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G33), .B(G41), .C1(new_n1008), .C2(G124), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n734), .A2(new_n474), .B1(new_n755), .B2(new_n308), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n758), .A2(new_n476), .B1(new_n746), .B2(new_n316), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n761), .A2(new_n376), .B1(new_n742), .B2(new_n807), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n922), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n384), .A2(new_n260), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT118), .B1(new_n1173), .B2(new_n1004), .ZN(new_n1174));
  OR3_X1    g0974(.A1(new_n1173), .A2(new_n1004), .A3(KEYINPUT118), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1173), .B(new_n216), .C1(G33), .C2(G41), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1168), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1157), .B1(new_n1181), .B2(new_n730), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1130), .B2(new_n776), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1156), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1125), .B1(new_n1155), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT120), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1187), .A2(new_n660), .A3(new_n1188), .A4(new_n1153), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1184), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(KEYINPUT121), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(G375));
  AOI22_X1  g0993(.A1(G97), .A2(new_n924), .B1(new_n747), .B2(G283), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n252), .B1(new_n759), .B2(G294), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1006), .A3(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G116), .A2(new_n735), .B1(new_n805), .B2(G107), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n754), .B2(new_n742), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G77), .C2(new_n762), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G132), .A2(new_n759), .B1(new_n747), .B2(G137), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n734), .B2(new_n1100), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n376), .A2(new_n761), .B1(new_n755), .B2(new_n275), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n753), .A2(new_n770), .B1(new_n742), .B2(new_n1095), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n781), .B1(new_n216), .B2(new_n749), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n730), .B1(new_n1199), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n787), .B1(new_n823), .B2(new_n335), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n1063), .C2(new_n776), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n1115), .B2(new_n725), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1116), .A2(new_n984), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1210), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT122), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT122), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(G381));
  NAND3_X1  g1017(.A1(new_n989), .A2(new_n791), .A3(new_n1027), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(G390), .A2(new_n1218), .A3(G384), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n986), .A2(new_n1215), .A3(new_n1216), .A4(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT123), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1120), .A2(new_n1106), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1192), .A3(new_n1222), .ZN(G407));
  NAND2_X1  g1023(.A1(new_n1192), .A2(new_n1222), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G407), .B(G213), .C1(G343), .C2(new_n1224), .ZN(G409));
  NAND3_X1  g1025(.A1(new_n642), .A2(G213), .A3(G2897), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1116), .A2(new_n661), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT125), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT60), .B1(new_n1212), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  AOI211_X1 g1030(.A(KEYINPUT125), .B(new_n1230), .C1(new_n1108), .C2(new_n1115), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1227), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT126), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT126), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n1227), .C1(new_n1229), .C2(new_n1231), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1210), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n826), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(G384), .A3(new_n1210), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1226), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G384), .B1(new_n1236), .B2(new_n1210), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n826), .B(new_n1209), .C1(new_n1233), .C2(new_n1235), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1226), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1240), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1189), .A2(G378), .A3(new_n1190), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1152), .A2(new_n726), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1183), .B(new_n1247), .C1(new_n1147), .C2(new_n984), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1222), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT124), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1248), .A2(new_n1222), .A3(KEYINPUT124), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1246), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n642), .A2(G213), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT61), .B1(new_n1245), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT62), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1253), .A2(new_n1257), .A3(new_n1254), .A4(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1253), .A2(new_n1254), .A3(new_n1258), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1256), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(new_n791), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(G390), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(G390), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1264), .A2(new_n986), .A3(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n986), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1262), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  OR2_X1    g1071(.A1(new_n1260), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1260), .A2(new_n1271), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1268), .A3(new_n1256), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1270), .A2(new_n1274), .ZN(G405));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1185), .A2(new_n1191), .A3(new_n1222), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1277), .A2(new_n1258), .A3(new_n1246), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1258), .B1(new_n1277), .B2(new_n1246), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1246), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1258), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1277), .A2(new_n1258), .A3(new_n1246), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(KEYINPUT127), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1280), .A2(new_n1285), .A3(new_n1269), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1268), .B(new_n1276), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(G402));
endmodule


