

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783;

  XNOR2_X1 U372 ( .A(n630), .B(n629), .ZN(n650) );
  AND2_X1 U373 ( .A1(n525), .A2(n526), .ZN(n628) );
  OR2_X1 U374 ( .A1(n572), .A2(n559), .ZN(n522) );
  NOR2_X2 U375 ( .A1(G953), .A2(G237), .ZN(n541) );
  AND2_X2 U376 ( .A1(n668), .A2(n520), .ZN(n376) );
  XNOR2_X2 U377 ( .A(n385), .B(n435), .ZN(n701) );
  INV_X1 U378 ( .A(G953), .ZN(n758) );
  XOR2_X1 U379 ( .A(n666), .B(n667), .Z(n351) );
  XNOR2_X1 U380 ( .A(n538), .B(n537), .ZN(n606) );
  AND2_X2 U381 ( .A1(n460), .A2(n657), .ZN(n450) );
  XNOR2_X2 U382 ( .A(G137), .B(n487), .ZN(n764) );
  INV_X2 U383 ( .A(n509), .ZN(n511) );
  XNOR2_X2 U384 ( .A(G113), .B(KEYINPUT95), .ZN(n509) );
  AND2_X1 U385 ( .A1(n699), .A2(n711), .ZN(n366) );
  XNOR2_X1 U386 ( .A(n446), .B(n560), .ZN(n681) );
  INV_X1 U387 ( .A(KEYINPUT10), .ZN(n464) );
  NAND2_X1 U388 ( .A1(n387), .A2(G210), .ZN(n356) );
  AND2_X1 U389 ( .A1(n391), .A2(n389), .ZN(n367) );
  AND2_X1 U390 ( .A1(n438), .A2(n641), .ZN(n437) );
  NAND2_X1 U391 ( .A1(n569), .A2(n366), .ZN(n571) );
  NOR2_X1 U392 ( .A1(n558), .A2(n436), .ZN(n634) );
  NOR2_X1 U393 ( .A1(n605), .A2(n426), .ZN(n568) );
  OR2_X1 U394 ( .A1(n377), .A2(n400), .ZN(n399) );
  NOR2_X1 U395 ( .A1(G902), .A2(n741), .ZN(n537) );
  XNOR2_X1 U396 ( .A(n536), .B(n535), .ZN(n741) );
  XNOR2_X1 U397 ( .A(n479), .B(KEYINPUT98), .ZN(n480) );
  INV_X1 U398 ( .A(n748), .ZN(n354) );
  XNOR2_X1 U399 ( .A(n464), .B(KEYINPUT79), .ZN(n465) );
  XNOR2_X1 U400 ( .A(G119), .B(G128), .ZN(n468) );
  XNOR2_X2 U401 ( .A(n511), .B(n510), .ZN(n513) );
  XNOR2_X1 U402 ( .A(n353), .B(n352), .ZN(G51) );
  INV_X1 U403 ( .A(KEYINPUT56), .ZN(n352) );
  NAND2_X1 U404 ( .A1(n355), .A2(n354), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n356), .B(n351), .ZN(n355) );
  XNOR2_X1 U406 ( .A(n754), .B(n396), .ZN(n357) );
  BUF_X1 U407 ( .A(n767), .Z(n358) );
  XNOR2_X1 U408 ( .A(n754), .B(n396), .ZN(n395) );
  BUF_X1 U409 ( .A(n749), .Z(n359) );
  BUF_X1 U410 ( .A(n549), .Z(n360) );
  NAND2_X1 U411 ( .A1(n401), .A2(n399), .ZN(n385) );
  NAND2_X2 U412 ( .A1(n448), .A2(n454), .ZN(n386) );
  INV_X1 U413 ( .A(n430), .ZN(n361) );
  XNOR2_X2 U414 ( .A(n549), .B(n548), .ZN(n754) );
  XNOR2_X2 U415 ( .A(n513), .B(n512), .ZN(n549) );
  NOR2_X1 U416 ( .A1(G902), .A2(G237), .ZN(n521) );
  INV_X1 U417 ( .A(n634), .ZN(n422) );
  INV_X1 U418 ( .A(KEYINPUT90), .ZN(n405) );
  XNOR2_X1 U419 ( .A(KEYINPUT66), .B(G101), .ZN(n492) );
  XNOR2_X1 U420 ( .A(n373), .B(KEYINPUT102), .ZN(n607) );
  INV_X1 U421 ( .A(KEYINPUT118), .ZN(n441) );
  XNOR2_X1 U422 ( .A(n421), .B(n420), .ZN(n438) );
  NAND2_X1 U423 ( .A1(n690), .A2(n677), .ZN(n373) );
  AND2_X1 U424 ( .A1(n708), .A2(n572), .ZN(n462) );
  XNOR2_X1 U425 ( .A(G134), .B(KEYINPUT69), .ZN(n486) );
  XOR2_X1 U426 ( .A(G131), .B(G140), .Z(n539) );
  XNOR2_X1 U427 ( .A(G146), .B(n764), .ZN(n508) );
  INV_X1 U428 ( .A(KEYINPUT2), .ZN(n453) );
  INV_X1 U429 ( .A(n459), .ZN(n457) );
  NAND2_X1 U430 ( .A1(n364), .A2(n656), .ZN(n402) );
  XNOR2_X1 U431 ( .A(n372), .B(KEYINPUT0), .ZN(n586) );
  NAND2_X1 U432 ( .A1(n681), .A2(n567), .ZN(n372) );
  NOR2_X1 U433 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U434 ( .A(G137), .B(G110), .ZN(n469) );
  XOR2_X1 U435 ( .A(KEYINPUT24), .B(G140), .Z(n470) );
  INV_X1 U436 ( .A(KEYINPUT23), .ZN(n467) );
  XOR2_X1 U437 ( .A(KEYINPUT82), .B(KEYINPUT8), .Z(n475) );
  XNOR2_X1 U438 ( .A(n419), .B(n418), .ZN(n417) );
  XNOR2_X1 U439 ( .A(G104), .B(G122), .ZN(n419) );
  XNOR2_X1 U440 ( .A(G113), .B(G143), .ZN(n418) );
  XNOR2_X1 U441 ( .A(n415), .B(KEYINPUT104), .ZN(n414) );
  INV_X1 U442 ( .A(KEYINPUT103), .ZN(n415) );
  XNOR2_X1 U443 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n413) );
  NAND2_X1 U444 ( .A1(n698), .A2(n699), .ZN(n440) );
  NAND2_X1 U445 ( .A1(n603), .A2(n463), .ZN(n716) );
  NOR2_X1 U446 ( .A1(n382), .A2(n383), .ZN(n622) );
  OR2_X1 U447 ( .A1(n572), .A2(n621), .ZN(n383) );
  NOR2_X1 U448 ( .A1(n394), .A2(KEYINPUT65), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n545), .B(n546), .ZN(n428) );
  XNOR2_X1 U450 ( .A(n572), .B(KEYINPUT6), .ZN(n635) );
  INV_X1 U451 ( .A(KEYINPUT76), .ZN(n420) );
  INV_X1 U452 ( .A(KEYINPUT86), .ZN(n380) );
  NOR2_X1 U453 ( .A1(n713), .A2(n463), .ZN(n714) );
  XOR2_X1 U454 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n515) );
  NOR2_X1 U455 ( .A1(n776), .A2(KEYINPUT44), .ZN(n594) );
  INV_X1 U456 ( .A(KEYINPUT38), .ZN(n435) );
  XNOR2_X1 U457 ( .A(n522), .B(n404), .ZN(n523) );
  XNOR2_X1 U458 ( .A(KEYINPUT30), .B(KEYINPUT117), .ZN(n404) );
  OR2_X1 U459 ( .A1(n462), .A2(KEYINPUT65), .ZN(n432) );
  INV_X1 U460 ( .A(KEYINPUT16), .ZN(n547) );
  XNOR2_X1 U461 ( .A(n508), .B(n409), .ZN(n498) );
  XNOR2_X1 U462 ( .A(n488), .B(n490), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n489), .B(KEYINPUT80), .ZN(n490) );
  NOR2_X1 U464 ( .A1(n459), .A2(n453), .ZN(n452) );
  AND2_X1 U465 ( .A1(n456), .A2(n455), .ZN(n454) );
  NAND2_X1 U466 ( .A1(n653), .A2(KEYINPUT2), .ZN(n461) );
  NAND2_X1 U467 ( .A1(G234), .A2(G237), .ZN(n501) );
  XNOR2_X1 U468 ( .A(n425), .B(KEYINPUT109), .ZN(n676) );
  NAND2_X1 U469 ( .A1(n427), .A2(n426), .ZN(n425) );
  BUF_X2 U470 ( .A(n581), .Z(n708) );
  XNOR2_X1 U471 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U472 ( .A(n363), .B(n471), .ZN(n472) );
  XNOR2_X1 U473 ( .A(n416), .B(n412), .ZN(n543) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n417), .B(n542), .ZN(n416) );
  AND2_X1 U476 ( .A1(n662), .A2(G953), .ZN(n748) );
  XNOR2_X1 U477 ( .A(n583), .B(KEYINPUT92), .ZN(n584) );
  NAND2_X1 U478 ( .A1(n648), .A2(n436), .ZN(n649) );
  NAND2_X1 U479 ( .A1(n682), .A2(n729), .ZN(n627) );
  XNOR2_X1 U480 ( .A(n604), .B(n374), .ZN(n690) );
  XNOR2_X1 U481 ( .A(n375), .B(KEYINPUT31), .ZN(n374) );
  INV_X1 U482 ( .A(KEYINPUT101), .ZN(n375) );
  NAND2_X1 U483 ( .A1(n430), .A2(n390), .ZN(n389) );
  NOR2_X1 U484 ( .A1(n597), .A2(n463), .ZN(n598) );
  OR2_X1 U485 ( .A1(n638), .A2(n676), .ZN(n362) );
  XOR2_X1 U486 ( .A(n468), .B(n467), .Z(n363) );
  AND2_X1 U487 ( .A1(n557), .A2(G210), .ZN(n364) );
  XNOR2_X1 U488 ( .A(n544), .B(n428), .ZN(n605) );
  INV_X1 U489 ( .A(n605), .ZN(n427) );
  AND2_X1 U490 ( .A1(G227), .A2(n758), .ZN(n365) );
  AND2_X1 U491 ( .A1(n461), .A2(n460), .ZN(n368) );
  INV_X1 U492 ( .A(n572), .ZN(n463) );
  AND2_X1 U493 ( .A1(n431), .A2(n394), .ZN(n369) );
  INV_X1 U494 ( .A(KEYINPUT113), .ZN(n394) );
  XOR2_X1 U495 ( .A(KEYINPUT84), .B(KEYINPUT48), .Z(n370) );
  XNOR2_X1 U496 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n371) );
  NAND2_X1 U497 ( .A1(n447), .A2(n700), .ZN(n446) );
  XNOR2_X2 U498 ( .A(n376), .B(G472), .ZN(n572) );
  XNOR2_X1 U499 ( .A(n357), .B(n555), .ZN(n377) );
  XNOR2_X1 U500 ( .A(n395), .B(n555), .ZN(n665) );
  AND2_X1 U501 ( .A1(n433), .A2(n369), .ZN(n378) );
  XNOR2_X2 U502 ( .A(n627), .B(KEYINPUT42), .ZN(n781) );
  XNOR2_X1 U503 ( .A(n594), .B(KEYINPUT67), .ZN(n379) );
  XNOR2_X1 U504 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U505 ( .A(n380), .B(n694), .ZN(n641) );
  BUF_X1 U506 ( .A(n681), .Z(n381) );
  NAND2_X1 U507 ( .A1(n619), .A2(n711), .ZN(n382) );
  NAND2_X1 U508 ( .A1(n361), .A2(n708), .ZN(n612) );
  AND2_X1 U509 ( .A1(n432), .A2(n619), .ZN(n431) );
  NAND2_X1 U510 ( .A1(n577), .A2(n434), .ZN(n433) );
  BUF_X1 U511 ( .A(n446), .Z(n384) );
  NAND2_X1 U512 ( .A1(n401), .A2(n399), .ZN(n447) );
  NAND2_X1 U513 ( .A1(n448), .A2(n454), .ZN(n387) );
  XNOR2_X2 U514 ( .A(n571), .B(n570), .ZN(n577) );
  NAND2_X1 U515 ( .A1(n433), .A2(n431), .ZN(n392) );
  NAND2_X1 U516 ( .A1(n378), .A2(n388), .ZN(n393) );
  NAND2_X1 U517 ( .A1(n430), .A2(n429), .ZN(n388) );
  NAND2_X1 U518 ( .A1(n392), .A2(KEYINPUT113), .ZN(n391) );
  NOR2_X2 U519 ( .A1(n579), .A2(n779), .ZN(n406) );
  NAND2_X1 U520 ( .A1(n393), .A2(n367), .ZN(n579) );
  XNOR2_X1 U521 ( .A(n397), .B(n553), .ZN(n396) );
  XNOR2_X1 U522 ( .A(n552), .B(n554), .ZN(n397) );
  AND2_X2 U523 ( .A1(n398), .A2(n402), .ZN(n401) );
  NAND2_X1 U524 ( .A1(n665), .A2(n364), .ZN(n398) );
  OR2_X1 U525 ( .A1(n364), .A2(n656), .ZN(n400) );
  NAND2_X1 U526 ( .A1(n628), .A2(n701), .ZN(n630) );
  XNOR2_X1 U527 ( .A(n403), .B(n371), .ZN(n439) );
  NAND2_X1 U528 ( .A1(n782), .A2(n781), .ZN(n403) );
  XNOR2_X1 U529 ( .A(n411), .B(n370), .ZN(n410) );
  AND2_X2 U530 ( .A1(n410), .A2(n652), .ZN(n654) );
  XNOR2_X2 U531 ( .A(n406), .B(n405), .ZN(n596) );
  XNOR2_X1 U532 ( .A(n532), .B(n407), .ZN(n534) );
  XNOR2_X1 U533 ( .A(n530), .B(n408), .ZN(n407) );
  INV_X1 U534 ( .A(n531), .ZN(n408) );
  XNOR2_X2 U535 ( .A(n654), .B(KEYINPUT83), .ZN(n767) );
  NAND2_X1 U536 ( .A1(n437), .A2(n439), .ZN(n411) );
  NAND2_X1 U537 ( .A1(n423), .A2(n422), .ZN(n421) );
  XNOR2_X1 U538 ( .A(n424), .B(n633), .ZN(n423) );
  NAND2_X1 U539 ( .A1(n682), .A2(n632), .ZN(n424) );
  INV_X1 U540 ( .A(n606), .ZN(n426) );
  INV_X1 U541 ( .A(KEYINPUT65), .ZN(n429) );
  INV_X1 U542 ( .A(n577), .ZN(n430) );
  AND2_X1 U543 ( .A1(n462), .A2(KEYINPUT65), .ZN(n434) );
  INV_X1 U544 ( .A(n385), .ZN(n436) );
  NAND2_X1 U545 ( .A1(n442), .A2(n617), .ZN(n618) );
  XNOR2_X2 U546 ( .A(n440), .B(n626), .ZN(n729) );
  XNOR2_X2 U547 ( .A(n625), .B(n441), .ZN(n698) );
  NAND2_X1 U548 ( .A1(n444), .A2(n443), .ZN(n442) );
  NAND2_X1 U549 ( .A1(n596), .A2(n595), .ZN(n443) );
  NAND2_X1 U550 ( .A1(n445), .A2(n379), .ZN(n444) );
  INV_X1 U551 ( .A(n596), .ZN(n445) );
  NOR2_X1 U552 ( .A1(n642), .A2(n384), .ZN(n639) );
  AND2_X2 U553 ( .A1(n449), .A2(n458), .ZN(n448) );
  NAND2_X1 U554 ( .A1(n450), .A2(n461), .ZN(n449) );
  NAND2_X1 U555 ( .A1(n655), .A2(n749), .ZN(n460) );
  NAND2_X1 U556 ( .A1(n451), .A2(n655), .ZN(n456) );
  AND2_X1 U557 ( .A1(n749), .A2(n457), .ZN(n451) );
  NAND2_X1 U558 ( .A1(n653), .A2(n452), .ZN(n458) );
  NAND2_X1 U559 ( .A1(n556), .A2(n657), .ZN(n455) );
  NAND2_X1 U560 ( .A1(n656), .A2(KEYINPUT64), .ZN(n459) );
  BUF_X1 U561 ( .A(n386), .Z(n744) );
  INV_X1 U562 ( .A(KEYINPUT97), .ZN(n489) );
  BUF_X1 U563 ( .A(n754), .Z(n755) );
  XNOR2_X1 U564 ( .A(n588), .B(KEYINPUT75), .ZN(n589) );
  BUF_X1 U565 ( .A(n579), .Z(n573) );
  XOR2_X2 U566 ( .A(G146), .B(G125), .Z(n554) );
  XNOR2_X1 U567 ( .A(n554), .B(n465), .ZN(n466) );
  XNOR2_X1 U568 ( .A(n466), .B(KEYINPUT72), .ZN(n473) );
  XNOR2_X1 U569 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U570 ( .A1(G234), .A2(n758), .ZN(n474) );
  XNOR2_X1 U571 ( .A(n475), .B(n474), .ZN(n527) );
  NAND2_X1 U572 ( .A1(G221), .A2(n527), .ZN(n476) );
  XNOR2_X1 U573 ( .A(n477), .B(n476), .ZN(n745) );
  NOR2_X1 U574 ( .A1(G902), .A2(n745), .ZN(n481) );
  XNOR2_X1 U575 ( .A(KEYINPUT15), .B(G902), .ZN(n556) );
  NAND2_X1 U576 ( .A1(G234), .A2(n556), .ZN(n478) );
  XNOR2_X1 U577 ( .A(KEYINPUT20), .B(n478), .ZN(n484) );
  NAND2_X1 U578 ( .A1(G217), .A2(n484), .ZN(n479) );
  XNOR2_X1 U579 ( .A(n481), .B(n480), .ZN(n483) );
  INV_X1 U580 ( .A(KEYINPUT25), .ZN(n482) );
  XNOR2_X2 U581 ( .A(n483), .B(n482), .ZN(n619) );
  INV_X1 U582 ( .A(n619), .ZN(n602) );
  AND2_X1 U583 ( .A1(n484), .A2(G221), .ZN(n485) );
  XNOR2_X1 U584 ( .A(n485), .B(KEYINPUT21), .ZN(n711) );
  NAND2_X1 U585 ( .A1(n602), .A2(n711), .ZN(n707) );
  INV_X1 U586 ( .A(n486), .ZN(n487) );
  XNOR2_X1 U587 ( .A(n539), .B(n365), .ZN(n488) );
  XNOR2_X2 U588 ( .A(G143), .B(G128), .ZN(n531) );
  XNOR2_X1 U589 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n491) );
  XNOR2_X1 U590 ( .A(n531), .B(n491), .ZN(n763) );
  XNOR2_X1 U591 ( .A(n763), .B(n492), .ZN(n507) );
  INV_X1 U592 ( .A(KEYINPUT94), .ZN(n493) );
  XNOR2_X1 U593 ( .A(n493), .B(G110), .ZN(n495) );
  XNOR2_X1 U594 ( .A(G107), .B(G104), .ZN(n494) );
  XNOR2_X1 U595 ( .A(n495), .B(n494), .ZN(n756) );
  INV_X1 U596 ( .A(KEYINPUT73), .ZN(n496) );
  XNOR2_X1 U597 ( .A(n756), .B(n496), .ZN(n497) );
  XNOR2_X1 U598 ( .A(n507), .B(n497), .ZN(n555) );
  XNOR2_X1 U599 ( .A(n498), .B(n555), .ZN(n735) );
  NOR2_X1 U600 ( .A1(n735), .A2(G902), .ZN(n500) );
  XNOR2_X1 U601 ( .A(KEYINPUT70), .B(G469), .ZN(n499) );
  XNOR2_X2 U602 ( .A(n500), .B(n499), .ZN(n623) );
  NOR2_X1 U603 ( .A1(n707), .A2(n623), .ZN(n526) );
  XNOR2_X1 U604 ( .A(n501), .B(KEYINPUT14), .ZN(n724) );
  INV_X1 U605 ( .A(n724), .ZN(n504) );
  NAND2_X1 U606 ( .A1(G953), .A2(G902), .ZN(n561) );
  NOR2_X1 U607 ( .A1(n504), .A2(n561), .ZN(n502) );
  XOR2_X1 U608 ( .A(KEYINPUT114), .B(n502), .Z(n503) );
  NOR2_X1 U609 ( .A1(G900), .A2(n503), .ZN(n506) );
  NAND2_X1 U610 ( .A1(n758), .A2(G952), .ZN(n565) );
  NOR2_X1 U611 ( .A1(n504), .A2(n565), .ZN(n505) );
  NOR2_X1 U612 ( .A1(n506), .A2(n505), .ZN(n621) );
  INV_X1 U613 ( .A(n621), .ZN(n524) );
  XNOR2_X1 U614 ( .A(n508), .B(n507), .ZN(n519) );
  XNOR2_X2 U615 ( .A(G119), .B(G116), .ZN(n510) );
  XOR2_X1 U616 ( .A(KEYINPUT71), .B(KEYINPUT3), .Z(n512) );
  NAND2_X1 U617 ( .A1(n541), .A2(G210), .ZN(n514) );
  XNOR2_X1 U618 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U619 ( .A(n516), .B(G131), .Z(n517) );
  XNOR2_X1 U620 ( .A(n360), .B(n517), .ZN(n518) );
  XNOR2_X1 U621 ( .A(n519), .B(n518), .ZN(n668) );
  INV_X1 U622 ( .A(G902), .ZN(n520) );
  XNOR2_X1 U623 ( .A(KEYINPUT77), .B(n521), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n557), .A2(G214), .ZN(n700) );
  AND2_X1 U625 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U626 ( .A(KEYINPUT108), .B(G478), .ZN(n538) );
  NAND2_X1 U627 ( .A1(G217), .A2(n527), .ZN(n536) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n529) );
  XNOR2_X1 U629 ( .A(G134), .B(G107), .ZN(n528) );
  XNOR2_X1 U630 ( .A(n529), .B(n528), .ZN(n532) );
  XOR2_X1 U631 ( .A(G122), .B(G116), .Z(n530) );
  XNOR2_X1 U632 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n533) );
  XNOR2_X1 U633 ( .A(n534), .B(n533), .ZN(n535) );
  INV_X1 U634 ( .A(G475), .ZN(n546) );
  XNOR2_X1 U635 ( .A(KEYINPUT13), .B(KEYINPUT105), .ZN(n545) );
  XOR2_X1 U636 ( .A(KEYINPUT10), .B(n554), .Z(n540) );
  XNOR2_X1 U637 ( .A(n540), .B(n539), .ZN(n766) );
  NAND2_X1 U638 ( .A1(G214), .A2(n541), .ZN(n542) );
  XNOR2_X1 U639 ( .A(n766), .B(n543), .ZN(n659) );
  NOR2_X1 U640 ( .A1(G902), .A2(n659), .ZN(n544) );
  NOR2_X1 U641 ( .A1(n606), .A2(n427), .ZN(n591) );
  NAND2_X1 U642 ( .A1(n628), .A2(n591), .ZN(n558) );
  XNOR2_X1 U643 ( .A(n547), .B(G122), .ZN(n548) );
  XOR2_X1 U644 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n551) );
  XNOR2_X1 U645 ( .A(KEYINPUT96), .B(KEYINPUT93), .ZN(n550) );
  XNOR2_X1 U646 ( .A(n551), .B(n550), .ZN(n553) );
  AND2_X1 U647 ( .A1(n758), .A2(G224), .ZN(n552) );
  INV_X1 U648 ( .A(n556), .ZN(n656) );
  XOR2_X1 U649 ( .A(G143), .B(n634), .Z(G45) );
  INV_X1 U650 ( .A(n700), .ZN(n559) );
  XNOR2_X1 U651 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n560) );
  INV_X1 U652 ( .A(G898), .ZN(n563) );
  INV_X1 U653 ( .A(n561), .ZN(n562) );
  NAND2_X1 U654 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U655 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U656 ( .A1(n724), .A2(n566), .ZN(n567) );
  INV_X1 U657 ( .A(n586), .ZN(n569) );
  XNOR2_X1 U658 ( .A(n568), .B(KEYINPUT110), .ZN(n699) );
  INV_X1 U659 ( .A(KEYINPUT22), .ZN(n570) );
  XNOR2_X1 U660 ( .A(n623), .B(KEYINPUT1), .ZN(n581) );
  XOR2_X1 U661 ( .A(n573), .B(G110), .Z(G12) );
  XNOR2_X1 U662 ( .A(KEYINPUT111), .B(n619), .ZN(n710) );
  NOR2_X1 U663 ( .A1(n710), .A2(n708), .ZN(n574) );
  XOR2_X1 U664 ( .A(KEYINPUT112), .B(n574), .Z(n575) );
  NOR2_X1 U665 ( .A1(n575), .A2(n635), .ZN(n576) );
  AND2_X1 U666 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U667 ( .A(n578), .B(KEYINPUT32), .ZN(n779) );
  INV_X1 U668 ( .A(n711), .ZN(n580) );
  NOR2_X2 U669 ( .A1(n581), .A2(n580), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n635), .A2(n601), .ZN(n582) );
  NOR2_X1 U671 ( .A1(n582), .A2(n619), .ZN(n585) );
  XNOR2_X1 U672 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n583) );
  XNOR2_X1 U673 ( .A(n585), .B(n584), .ZN(n730) );
  BUF_X1 U674 ( .A(n586), .Z(n587) );
  NOR2_X1 U675 ( .A1(n730), .A2(n587), .ZN(n590) );
  XNOR2_X1 U676 ( .A(KEYINPUT34), .B(KEYINPUT81), .ZN(n588) );
  XNOR2_X1 U677 ( .A(n590), .B(n589), .ZN(n592) );
  NAND2_X1 U678 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X2 U679 ( .A(n593), .B(KEYINPUT35), .ZN(n776) );
  INV_X1 U680 ( .A(KEYINPUT44), .ZN(n595) );
  INV_X1 U681 ( .A(n587), .ZN(n599) );
  OR2_X1 U682 ( .A1(n623), .A2(n707), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U684 ( .A(KEYINPUT100), .B(n600), .ZN(n677) );
  AND2_X1 U685 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U686 ( .A1(n587), .A2(n716), .ZN(n604) );
  NAND2_X1 U687 ( .A1(n606), .A2(n605), .ZN(n687) );
  INV_X1 U688 ( .A(n687), .ZN(n638) );
  NAND2_X1 U689 ( .A1(n607), .A2(n362), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n776), .A2(KEYINPUT44), .ZN(n609) );
  INV_X1 U691 ( .A(KEYINPUT89), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n612), .A2(n635), .ZN(n613) );
  XNOR2_X1 U694 ( .A(n613), .B(KEYINPUT88), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n614), .A2(n710), .ZN(n674) );
  INV_X1 U696 ( .A(n674), .ZN(n615) );
  XNOR2_X2 U697 ( .A(n618), .B(KEYINPUT45), .ZN(n749) );
  NAND2_X1 U698 ( .A1(n619), .A2(n711), .ZN(n620) );
  NOR2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n636) );
  XOR2_X1 U700 ( .A(KEYINPUT28), .B(n622), .Z(n624) );
  NOR2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n682) );
  XOR2_X1 U702 ( .A(KEYINPUT119), .B(KEYINPUT41), .Z(n626) );
  NAND2_X1 U703 ( .A1(n701), .A2(n700), .ZN(n625) );
  XOR2_X1 U704 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n629) );
  NAND2_X1 U705 ( .A1(n650), .A2(n638), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT40), .ZN(n782) );
  INV_X1 U707 ( .A(KEYINPUT47), .ZN(n633) );
  AND2_X1 U708 ( .A1(n381), .A2(n362), .ZN(n632) );
  AND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n642) );
  XOR2_X1 U711 ( .A(KEYINPUT36), .B(n639), .Z(n640) );
  NOR2_X1 U712 ( .A1(n708), .A2(n640), .ZN(n694) );
  INV_X1 U713 ( .A(n708), .ZN(n645) );
  INV_X1 U714 ( .A(n642), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n643), .A2(n700), .ZN(n644) );
  NOR2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n647) );
  XNOR2_X1 U717 ( .A(KEYINPUT115), .B(KEYINPUT43), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(n648) );
  XOR2_X1 U719 ( .A(KEYINPUT116), .B(n649), .Z(n777) );
  NAND2_X1 U720 ( .A1(n650), .A2(n676), .ZN(n697) );
  INV_X1 U721 ( .A(n697), .ZN(n651) );
  NOR2_X1 U722 ( .A1(n777), .A2(n651), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n749), .A2(n654), .ZN(n653) );
  NOR2_X2 U724 ( .A1(n767), .A2(KEYINPUT2), .ZN(n655) );
  INV_X1 U725 ( .A(KEYINPUT64), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n386), .A2(G475), .ZN(n661) );
  XOR2_X1 U727 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(n660), .ZN(n663) );
  INV_X1 U730 ( .A(G952), .ZN(n662) );
  NOR2_X2 U731 ( .A1(n663), .A2(n748), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n664), .B(KEYINPUT60), .ZN(G60) );
  BUF_X1 U733 ( .A(n377), .Z(n666) );
  XOR2_X1 U734 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n667) );
  NAND2_X1 U735 ( .A1(n386), .A2(G472), .ZN(n670) );
  XOR2_X1 U736 ( .A(KEYINPUT62), .B(n668), .Z(n669) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X2 U738 ( .A1(n671), .A2(n748), .ZN(n673) );
  XNOR2_X1 U739 ( .A(KEYINPUT91), .B(KEYINPUT63), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n673), .B(n672), .ZN(G57) );
  XNOR2_X1 U741 ( .A(G101), .B(n674), .ZN(G3) );
  NOR2_X1 U742 ( .A1(n677), .A2(n687), .ZN(n675) );
  XOR2_X1 U743 ( .A(G104), .B(n675), .Z(G6) );
  INV_X1 U744 ( .A(n676), .ZN(n691) );
  NOR2_X1 U745 ( .A1(n677), .A2(n691), .ZN(n679) );
  XNOR2_X1 U746 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U748 ( .A(G107), .B(n680), .ZN(G9) );
  NAND2_X1 U749 ( .A1(n682), .A2(n381), .ZN(n685) );
  NOR2_X1 U750 ( .A1(n685), .A2(n691), .ZN(n684) );
  XNOR2_X1 U751 ( .A(G128), .B(KEYINPUT29), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n684), .B(n683), .ZN(G30) );
  NOR2_X1 U753 ( .A1(n685), .A2(n687), .ZN(n686) );
  XOR2_X1 U754 ( .A(G146), .B(n686), .Z(G48) );
  NOR2_X1 U755 ( .A1(n687), .A2(n690), .ZN(n688) );
  XOR2_X1 U756 ( .A(KEYINPUT120), .B(n688), .Z(n689) );
  XNOR2_X1 U757 ( .A(G113), .B(n689), .ZN(G15) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n693) );
  XNOR2_X1 U759 ( .A(G116), .B(KEYINPUT121), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n693), .B(n692), .ZN(G18) );
  XNOR2_X1 U761 ( .A(n694), .B(KEYINPUT37), .ZN(n695) );
  XNOR2_X1 U762 ( .A(n695), .B(KEYINPUT122), .ZN(n696) );
  XNOR2_X1 U763 ( .A(G125), .B(n696), .ZN(G27) );
  XNOR2_X1 U764 ( .A(G134), .B(n697), .ZN(G36) );
  AND2_X1 U765 ( .A1(n698), .A2(n362), .ZN(n705) );
  INV_X1 U766 ( .A(n699), .ZN(n703) );
  NOR2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U769 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U770 ( .A1(n730), .A2(n706), .ZN(n722) );
  NAND2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U772 ( .A(n709), .B(KEYINPUT50), .ZN(n715) );
  NOR2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U774 ( .A(KEYINPUT49), .B(n712), .Z(n713) );
  NAND2_X1 U775 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U776 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U777 ( .A(KEYINPUT51), .B(n718), .Z(n719) );
  NAND2_X1 U778 ( .A1(n729), .A2(n719), .ZN(n720) );
  XOR2_X1 U779 ( .A(KEYINPUT124), .B(n720), .Z(n721) );
  NOR2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U781 ( .A(KEYINPUT52), .B(n723), .ZN(n726) );
  NAND2_X1 U782 ( .A1(n724), .A2(G952), .ZN(n725) );
  NOR2_X1 U783 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U784 ( .A1(n727), .A2(G953), .ZN(n728) );
  NAND2_X1 U785 ( .A1(n368), .A2(n728), .ZN(n733) );
  INV_X1 U786 ( .A(n729), .ZN(n731) );
  NOR2_X1 U787 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U788 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U789 ( .A(KEYINPUT53), .B(n734), .ZN(G75) );
  XOR2_X1 U790 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n737) );
  XNOR2_X1 U791 ( .A(n735), .B(KEYINPUT125), .ZN(n736) );
  XNOR2_X1 U792 ( .A(n737), .B(n736), .ZN(n739) );
  NAND2_X1 U793 ( .A1(n387), .A2(G469), .ZN(n738) );
  XOR2_X1 U794 ( .A(n739), .B(n738), .Z(n740) );
  NOR2_X1 U795 ( .A1(n748), .A2(n740), .ZN(G54) );
  NAND2_X1 U796 ( .A1(n744), .A2(G478), .ZN(n742) );
  XNOR2_X1 U797 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U798 ( .A1(n748), .A2(n743), .ZN(G63) );
  NAND2_X1 U799 ( .A1(n744), .A2(G217), .ZN(n746) );
  XNOR2_X1 U800 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U801 ( .A1(n748), .A2(n747), .ZN(G66) );
  NAND2_X1 U802 ( .A1(n359), .A2(n758), .ZN(n753) );
  NAND2_X1 U803 ( .A1(G953), .A2(G224), .ZN(n750) );
  XNOR2_X1 U804 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U805 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U806 ( .A1(n753), .A2(n752), .ZN(n762) );
  XNOR2_X1 U807 ( .A(n755), .B(G101), .ZN(n757) );
  XNOR2_X1 U808 ( .A(n757), .B(n756), .ZN(n760) );
  NOR2_X1 U809 ( .A1(G898), .A2(n758), .ZN(n759) );
  NOR2_X1 U810 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U811 ( .A(n762), .B(n761), .ZN(G69) );
  XNOR2_X1 U812 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U813 ( .A(n766), .B(n765), .ZN(n771) );
  INV_X1 U814 ( .A(n771), .ZN(n768) );
  XNOR2_X1 U815 ( .A(n768), .B(n358), .ZN(n769) );
  NOR2_X1 U816 ( .A1(G953), .A2(n769), .ZN(n770) );
  XNOR2_X1 U817 ( .A(KEYINPUT127), .B(n770), .ZN(n775) );
  XNOR2_X1 U818 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U819 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U820 ( .A1(n773), .A2(G953), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n775), .A2(n774), .ZN(G72) );
  XOR2_X1 U822 ( .A(n776), .B(G122), .Z(G24) );
  XNOR2_X1 U823 ( .A(G140), .B(KEYINPUT123), .ZN(n778) );
  XNOR2_X1 U824 ( .A(n778), .B(n777), .ZN(G42) );
  INV_X1 U825 ( .A(n779), .ZN(n780) );
  XNOR2_X1 U826 ( .A(G119), .B(n780), .ZN(G21) );
  XNOR2_X1 U827 ( .A(G137), .B(n781), .ZN(G39) );
  BUF_X1 U828 ( .A(n782), .Z(n783) );
  XNOR2_X1 U829 ( .A(G131), .B(n783), .ZN(G33) );
endmodule

