//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(KEYINPUT64), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n209), .B1(new_n210), .B2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G13), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n212), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n205), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n210), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G20), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n216), .B(new_n226), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n219), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  AOI21_X1  g0049(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT67), .ZN(new_n253));
  INV_X1    g0053(.A(G223), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n251), .A2(G222), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n259), .B2(KEYINPUT66), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(KEYINPUT66), .B2(new_n257), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n250), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G274), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n250), .A2(new_n268), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(G226), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G200), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT68), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n227), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G1), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n283), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n288), .A2(new_n291), .B1(new_n202), .B2(new_n287), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT9), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n274), .B(new_n294), .C1(new_n295), .C2(new_n273), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(new_n275), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n280), .A2(new_n298), .B1(new_n277), .B2(new_n258), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT15), .B(G87), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(new_n278), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n283), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n288), .A2(G77), .A3(new_n289), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n302), .B(new_n303), .C1(G77), .C2(new_n286), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n270), .B1(G244), .B2(new_n271), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n251), .A2(G232), .A3(new_n256), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n206), .B2(new_n251), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT67), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n252), .B(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n309), .B2(G238), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n305), .B1(new_n310), .B2(new_n264), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n304), .B1(new_n312), .B2(G190), .ZN(new_n313));
  INV_X1    g0113(.A(G200), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n312), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n317), .A2(new_n304), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n251), .A2(G232), .A3(G1698), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n251), .A2(G226), .A3(new_n256), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n250), .ZN(new_n327));
  INV_X1    g0127(.A(new_n265), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n268), .B1(new_n271), .B2(G238), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT13), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n327), .A2(new_n332), .A3(new_n329), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(G190), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT70), .B1(new_n277), .B2(G68), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n298), .B2(new_n202), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n275), .A2(KEYINPUT70), .A3(G50), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n336), .B(new_n337), .C1(new_n279), .C2(new_n258), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(KEYINPUT11), .A3(new_n283), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT12), .B1(new_n286), .B2(G68), .ZN(new_n340));
  OR3_X1    g0140(.A1(new_n286), .A2(KEYINPUT12), .A3(G68), .ZN(new_n341));
  INV_X1    g0141(.A(G68), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n285), .B2(G20), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n340), .A2(new_n341), .B1(new_n288), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT11), .B1(new_n338), .B2(new_n283), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n334), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n331), .A2(new_n333), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT69), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(G200), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n327), .A2(new_n332), .A3(new_n329), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n332), .B1(new_n327), .B2(new_n329), .ZN(new_n353));
  OAI21_X1  g0153(.A(G200), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT69), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n348), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n352), .A2(new_n353), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT14), .B1(new_n357), .B2(new_n316), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n349), .A2(new_n359), .A3(G169), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT71), .B1(new_n357), .B2(G179), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT71), .ZN(new_n362));
  NOR4_X1   g0162(.A1(new_n352), .A2(new_n353), .A3(new_n362), .A4(new_n319), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n358), .B(new_n360), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n346), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(new_n339), .A3(new_n344), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n356), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n273), .A2(new_n316), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n293), .C1(G179), .C2(new_n273), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n297), .A2(new_n322), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n251), .B2(G20), .ZN(new_n372));
  INV_X1    g0172(.A(G33), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT3), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G33), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(KEYINPUT7), .A3(new_n277), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G68), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n218), .A2(new_n342), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n381), .B2(new_n201), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n275), .A2(G159), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n380), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n342), .B1(new_n372), .B2(new_n378), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(new_n384), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n389), .A3(new_n283), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n280), .B1(new_n285), .B2(G20), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n288), .B1(new_n287), .B2(new_n280), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n374), .A2(new_n376), .A3(G226), .A4(G1698), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G87), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n374), .A2(new_n376), .A3(G223), .A4(new_n256), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n251), .A2(KEYINPUT72), .A3(G223), .A4(new_n256), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n264), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n271), .A2(G232), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n265), .B2(new_n269), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n316), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n401), .B2(new_n264), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n399), .A2(new_n400), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT73), .B(new_n250), .C1(new_n408), .C2(new_n396), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n404), .A2(G179), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n393), .A2(KEYINPUT18), .A3(new_n405), .A4(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT74), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n411), .A2(new_n405), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n415), .A2(KEYINPUT74), .A3(KEYINPUT18), .A4(new_n393), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n393), .A2(new_n405), .A3(new_n411), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n390), .A2(new_n392), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n314), .B1(new_n402), .B2(new_n404), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n409), .A2(new_n407), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n404), .A2(G190), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT17), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT17), .B1(new_n421), .B2(new_n425), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n420), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(KEYINPUT75), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(KEYINPUT75), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n370), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n267), .A2(G1), .ZN(new_n433));
  AND2_X1   g0233(.A1(KEYINPUT5), .A2(G41), .ZN(new_n434));
  NOR2_X1   g0234(.A1(KEYINPUT5), .A2(G41), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n265), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT5), .B(G41), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(new_n433), .B1(new_n228), .B2(new_n263), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(G270), .B2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n374), .A2(new_n376), .A3(G264), .A4(G1698), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n374), .A2(new_n376), .A3(G257), .A4(new_n256), .ZN(new_n442));
  INV_X1    g0242(.A(G303), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n251), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n250), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n314), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n285), .A2(G33), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n288), .A2(G116), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G116), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n287), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n282), .A2(new_n227), .B1(G20), .B2(new_n449), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n277), .C1(G33), .C2(new_n205), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n451), .A2(KEYINPUT20), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT20), .B1(new_n451), .B2(new_n453), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n448), .B(new_n450), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  OR3_X1    g0256(.A1(new_n446), .A2(KEYINPUT82), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT82), .B1(new_n446), .B2(new_n456), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n440), .A2(new_n445), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n295), .C2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n445), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n265), .A2(new_n436), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n436), .A2(new_n264), .ZN(new_n463));
  INV_X1    g0263(.A(G270), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n456), .B(G169), .C1(new_n461), .C2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT21), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n459), .A2(KEYINPUT21), .A3(G169), .A4(new_n456), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n456), .A2(G179), .A3(new_n445), .A4(new_n440), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n460), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n251), .A2(new_n277), .A3(G68), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT19), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n277), .B1(new_n325), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(G87), .B2(new_n207), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n278), .B2(new_n205), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n479), .A2(new_n283), .B1(new_n287), .B2(new_n300), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n282), .A2(new_n227), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n481), .A2(new_n286), .A3(new_n447), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G87), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n285), .A2(G45), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n264), .A2(G250), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n265), .B2(new_n484), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n251), .A2(G244), .A3(G1698), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n251), .A2(G238), .A3(new_n256), .ZN(new_n488));
  AND2_X1   g0288(.A1(G33), .A2(G116), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n486), .B1(new_n491), .B2(new_n250), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n480), .B(new_n483), .C1(new_n492), .C2(new_n314), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n493), .A2(KEYINPUT81), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n493), .A2(KEYINPUT81), .B1(G190), .B2(new_n492), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n479), .A2(new_n283), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n300), .A2(new_n287), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n481), .A2(new_n286), .A3(new_n447), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n498), .C1(new_n499), .C2(new_n300), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n492), .A2(new_n319), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(new_n501), .C1(G169), .C2(new_n492), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n374), .A2(new_n376), .A3(new_n277), .A4(G87), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT22), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(KEYINPUT22), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n251), .A2(new_n277), .A3(G87), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT84), .B1(new_n277), .B2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(KEYINPUT85), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT84), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT85), .B1(new_n513), .B2(new_n511), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n206), .A2(G20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n489), .A2(new_n277), .B1(new_n517), .B2(KEYINPUT23), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n512), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n509), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT24), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n481), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n512), .A2(new_n516), .A3(new_n518), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n508), .B2(new_n506), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT24), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n482), .A2(G107), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT86), .ZN(new_n527));
  OR3_X1    g0327(.A1(new_n286), .A2(KEYINPUT25), .A3(G107), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT25), .B1(new_n286), .B2(G107), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n528), .B(new_n529), .C1(new_n499), .C2(new_n206), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT86), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n522), .A2(new_n525), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n374), .A2(new_n376), .A3(G257), .A4(G1698), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n374), .A2(new_n376), .A3(G250), .A4(new_n256), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G294), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n250), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n439), .A2(G264), .ZN(new_n539));
  AND4_X1   g0339(.A1(new_n295), .A2(new_n538), .A3(new_n462), .A4(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n537), .A2(new_n250), .B1(new_n439), .B2(G264), .ZN(new_n541));
  AOI21_X1  g0341(.A(G200), .B1(new_n541), .B2(new_n462), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n533), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n530), .A2(new_n532), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n283), .B1(new_n524), .B2(KEYINPUT24), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n520), .A2(new_n521), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n541), .A2(new_n319), .A3(new_n462), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n541), .A2(new_n462), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n316), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n473), .A2(new_n503), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT80), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n374), .A2(new_n376), .A3(G244), .A4(new_n256), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT4), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n377), .A2(KEYINPUT76), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT76), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n251), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n557), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(G250), .A2(G1698), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n374), .A2(new_n376), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT77), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n251), .A2(KEYINPUT77), .A3(new_n564), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n452), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n250), .B1(new_n563), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT79), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n463), .B2(new_n220), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n436), .A2(KEYINPUT79), .A3(G257), .A4(new_n264), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n462), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(G179), .ZN(new_n577));
  OAI211_X1 g0377(.A(KEYINPUT78), .B(new_n250), .C1(new_n563), .C2(new_n569), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n572), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT76), .B1(new_n377), .B2(new_n558), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n251), .A2(new_n560), .A3(new_n561), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n580), .A2(new_n581), .B1(new_n556), .B2(new_n555), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n567), .A2(new_n568), .A3(new_n452), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n264), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n316), .B1(new_n584), .B2(new_n576), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT6), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n586), .A2(new_n205), .A3(G107), .ZN(new_n587));
  XNOR2_X1  g0387(.A(G97), .B(G107), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n589), .A2(new_n277), .B1(new_n258), .B2(new_n298), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n206), .B1(new_n372), .B2(new_n378), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n283), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n286), .A2(G97), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n482), .B2(G97), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n585), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n554), .B1(new_n579), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n462), .A2(new_n575), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT79), .B1(new_n439), .B2(G257), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n572), .A2(new_n578), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G200), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n584), .A2(new_n576), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n595), .B1(new_n603), .B2(G190), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n570), .A2(new_n600), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(new_n316), .B1(new_n592), .B2(new_n594), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n572), .A2(new_n577), .A3(new_n578), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(KEYINPUT80), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n597), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n553), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n432), .A2(new_n612), .ZN(G372));
  INV_X1    g0413(.A(new_n502), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n494), .B2(new_n495), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n607), .A2(KEYINPUT80), .A3(new_n608), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT80), .B1(new_n607), .B2(new_n608), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n615), .B(KEYINPUT26), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n492), .A2(G169), .ZN(new_n619));
  AOI211_X1 g0419(.A(G179), .B(new_n486), .C1(new_n491), .C2(new_n250), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n491), .A2(new_n250), .ZN(new_n622));
  INV_X1    g0422(.A(new_n486), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n314), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n497), .A2(new_n498), .A3(new_n483), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n492), .A2(G190), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n621), .A2(new_n500), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(new_n608), .A3(new_n607), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT88), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n607), .A2(new_n608), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n622), .A2(new_n623), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  INV_X1    g0435(.A(new_n625), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n627), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n502), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n631), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT88), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n618), .A2(new_n632), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n502), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n616), .A2(new_n617), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n540), .A2(new_n542), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n637), .B(new_n502), .C1(new_n547), .C2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n472), .B2(new_n551), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n644), .A2(new_n647), .A3(KEYINPUT87), .A4(new_n605), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n550), .A2(new_n548), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n533), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n628), .B(new_n543), .C1(new_n651), .C2(new_n471), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n649), .B1(new_n610), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n643), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n432), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n369), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n321), .A2(new_n356), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n358), .A2(new_n360), .ZN(new_n659));
  INV_X1    g0459(.A(new_n363), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n362), .B1(new_n349), .B2(new_n319), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n347), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n428), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n419), .A2(new_n412), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n657), .B1(new_n666), .B2(new_n297), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n656), .A2(new_n667), .ZN(G369));
  NAND3_X1  g0468(.A1(new_n285), .A2(new_n277), .A3(G13), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT89), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n675), .A2(new_n456), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n471), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n473), .B2(new_n676), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n551), .A2(new_n675), .ZN(new_n680));
  INV_X1    g0480(.A(new_n675), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n543), .B1(new_n533), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n680), .B1(new_n682), .B2(new_n551), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n472), .A2(new_n675), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n680), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(G399));
  NOR3_X1   g0487(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT90), .Z(new_n689));
  INV_X1    g0489(.A(new_n214), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n692), .A3(G1), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n232), .B2(new_n692), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT91), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n675), .B1(new_n643), .B2(new_n654), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n601), .A2(new_n549), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n459), .A2(new_n634), .A3(new_n319), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n440), .A2(G179), .A3(new_n445), .ZN(new_n705));
  INV_X1    g0505(.A(new_n541), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n634), .A3(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n707), .A2(KEYINPUT30), .A3(new_n603), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT30), .B1(new_n707), .B2(new_n603), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n675), .B1(new_n704), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n700), .B(KEYINPUT92), .ZN(new_n715));
  INV_X1    g0515(.A(new_n703), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n681), .B1(new_n717), .B2(new_n710), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT31), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n553), .A2(new_n611), .A3(new_n681), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n714), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT93), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n644), .A2(new_n647), .A3(new_n723), .A4(new_n605), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT93), .B1(new_n610), .B2(new_n652), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n597), .A2(new_n609), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n631), .A3(new_n615), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n614), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n724), .A2(new_n725), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n681), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n699), .A2(new_n722), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n696), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(new_n678), .A2(G330), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT94), .ZN(new_n736));
  INV_X1    g0536(.A(new_n679), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n212), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n285), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n691), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n736), .A2(new_n737), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n214), .A2(G355), .A3(new_n251), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G116), .B2(new_n214), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n245), .A2(new_n267), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n251), .B(new_n690), .C1(new_n267), .C2(new_n233), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n227), .B1(G20), .B2(new_n316), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n742), .ZN(new_n756));
  INV_X1    g0556(.A(new_n751), .ZN(new_n757));
  INV_X1    g0557(.A(new_n752), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n277), .A2(new_n295), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n319), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n277), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n760), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n761), .A2(new_n218), .B1(new_n763), .B2(new_n258), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n277), .A2(new_n319), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(G190), .A3(G200), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(KEYINPUT95), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(KEYINPUT95), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n764), .B1(new_n770), .B2(G50), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT96), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n277), .B1(new_n773), .B2(G190), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT98), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT98), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n205), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n314), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n762), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G87), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n759), .A2(new_n779), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n251), .B1(new_n780), .B2(new_n206), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n762), .A2(new_n773), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT97), .B(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n765), .A2(new_n295), .A3(G200), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n342), .B2(new_n788), .ZN(new_n789));
  NOR4_X1   g0589(.A1(new_n772), .A2(new_n778), .A3(new_n783), .A4(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT99), .B(G326), .Z(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n769), .A2(new_n791), .B1(new_n792), .B2(new_n777), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(KEYINPUT100), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(KEYINPUT100), .ZN(new_n795));
  INV_X1    g0595(.A(new_n761), .ZN(new_n796));
  INV_X1    g0596(.A(new_n784), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G322), .A2(new_n796), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n798), .B1(new_n799), .B2(new_n780), .C1(new_n800), .C2(new_n763), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT33), .B(G317), .Z(new_n802));
  OAI221_X1 g0602(.A(new_n377), .B1(new_n782), .B2(new_n443), .C1(new_n788), .C2(new_n802), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n794), .A2(new_n795), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n790), .A2(new_n804), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n756), .B1(new_n678), .B2(new_n757), .C1(new_n758), .C2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n743), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NOR2_X1   g0608(.A1(new_n321), .A2(new_n675), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n675), .A2(new_n304), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n315), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(new_n811), .B2(new_n321), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n697), .B(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n741), .B1(new_n813), .B2(new_n722), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n722), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n752), .A2(new_n749), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n742), .B1(new_n258), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n769), .A2(new_n443), .ZN(new_n818));
  INV_X1    g0618(.A(new_n782), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G107), .A2(new_n819), .B1(new_n797), .B2(G311), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n762), .A2(new_n779), .A3(G87), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n792), .C2(new_n761), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n377), .B1(new_n763), .B2(new_n449), .C1(new_n788), .C2(new_n799), .ZN(new_n823));
  NOR4_X1   g0623(.A1(new_n818), .A2(new_n822), .A3(new_n778), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n251), .B1(new_n782), .B2(new_n202), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n780), .A2(new_n342), .B1(new_n784), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n777), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n825), .B(new_n827), .C1(new_n828), .C2(G58), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT101), .ZN(new_n830));
  INV_X1    g0630(.A(new_n763), .ZN(new_n831));
  INV_X1    g0631(.A(new_n785), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G143), .A2(new_n796), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G150), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n834), .B2(new_n788), .C1(new_n769), .C2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT34), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n824), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n817), .B1(new_n758), .B2(new_n838), .C1(new_n812), .C2(new_n750), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n815), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  XOR2_X1   g0641(.A(new_n589), .B(KEYINPUT102), .Z(new_n842));
  INV_X1    g0642(.A(KEYINPUT35), .ZN(new_n843));
  OAI211_X1 g0643(.A(G116), .B(new_n230), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n843), .B2(new_n842), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT36), .ZN(new_n846));
  OR3_X1    g0646(.A1(new_n232), .A2(new_n258), .A3(new_n381), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n202), .A2(G68), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n285), .B(G13), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n699), .A2(new_n731), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n432), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n667), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n364), .A2(new_n366), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n355), .A2(new_n351), .ZN(new_n855));
  INV_X1    g0655(.A(new_n348), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(KEYINPUT103), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n681), .A2(new_n347), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n364), .A2(new_n860), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n862), .B(new_n857), .C1(new_n663), .C2(KEYINPUT103), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n648), .A2(new_n653), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n681), .B(new_n812), .C1(new_n865), .C2(new_n642), .ZN(new_n866));
  INV_X1    g0666(.A(new_n809), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n673), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n390), .A2(KEYINPUT104), .A3(new_n392), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT104), .B1(new_n390), .B2(new_n392), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n420), .B2(new_n428), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n415), .B1(new_n870), .B2(new_n871), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n421), .A2(new_n425), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n393), .A2(new_n869), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n417), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(KEYINPUT37), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n874), .A2(new_n881), .A3(KEYINPUT38), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(KEYINPUT37), .B2(new_n877), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n885), .B2(new_n873), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n868), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n419), .A2(new_n412), .A3(new_n673), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n854), .A2(new_n675), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n885), .A2(new_n873), .A3(new_n883), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n428), .A2(new_n665), .ZN(new_n894));
  INV_X1    g0694(.A(new_n879), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n880), .B(KEYINPUT37), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n892), .B1(new_n893), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n882), .A2(new_n886), .A3(KEYINPUT39), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n888), .B(new_n889), .C1(new_n891), .C2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n853), .B(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(G330), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(new_n884), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n879), .B1(new_n428), .B2(new_n665), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n883), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n882), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n861), .A2(new_n812), .A3(new_n863), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n721), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT40), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n721), .A2(new_n887), .A3(new_n914), .A4(new_n911), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n432), .A2(new_n721), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n904), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n917), .B2(new_n916), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n903), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n285), .B2(new_n738), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n903), .A2(new_n919), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n850), .B1(new_n921), .B2(new_n922), .ZN(G367));
  INV_X1    g0723(.A(KEYINPUT107), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT106), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n675), .A2(new_n595), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n644), .A2(new_n605), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n607), .A2(new_n608), .A3(new_n675), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n683), .A3(new_n685), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT42), .Z(new_n931));
  AOI21_X1  g0731(.A(new_n726), .B1(new_n929), .B2(new_n651), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n675), .B1(new_n932), .B2(KEYINPUT105), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(KEYINPUT105), .B2(new_n932), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n925), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n675), .A2(new_n625), .ZN(new_n936));
  MUX2_X1   g0736(.A(new_n614), .B(new_n628), .S(new_n936), .Z(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT43), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n931), .A2(new_n934), .A3(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n935), .B2(new_n938), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n929), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n684), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n924), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n929), .A2(new_n686), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n929), .A2(new_n686), .ZN(new_n949));
  XOR2_X1   g0749(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n948), .A2(new_n684), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n684), .B1(new_n948), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n683), .B(new_n685), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(new_n679), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n732), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n691), .B(KEYINPUT41), .Z(new_n958));
  OAI21_X1  g0758(.A(new_n739), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n942), .A2(new_n945), .ZN(new_n960));
  OAI211_X1 g0760(.A(KEYINPUT107), .B(new_n944), .C1(new_n939), .C2(new_n941), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n946), .A2(new_n959), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n690), .A2(new_n251), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n241), .ZN(new_n964));
  INV_X1    g0764(.A(new_n300), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n754), .B1(new_n690), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n742), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n788), .A2(new_n792), .ZN(new_n968));
  INV_X1    g0768(.A(G317), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n782), .A2(new_n449), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n377), .B1(new_n969), .B2(new_n784), .C1(new_n970), .C2(KEYINPUT46), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n968), .B(new_n971), .C1(KEYINPUT46), .C2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n763), .A2(new_n799), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n780), .A2(new_n205), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(G303), .C2(new_n796), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n770), .A2(G311), .B1(G107), .B2(new_n828), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n972), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n770), .A2(G143), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n780), .A2(new_n258), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n763), .A2(new_n202), .B1(new_n784), .B2(new_n835), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(G150), .C2(new_n796), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n828), .A2(G68), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n251), .B1(new_n782), .B2(new_n218), .ZN(new_n983));
  INV_X1    g0783(.A(new_n788), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n983), .B1(new_n984), .B2(new_n832), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n978), .A2(new_n981), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n977), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT47), .Z(new_n988));
  OAI221_X1 g0788(.A(new_n967), .B1(new_n757), .B2(new_n937), .C1(new_n988), .C2(new_n758), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n962), .A2(new_n989), .ZN(G387));
  NAND2_X1  g0790(.A1(new_n956), .A2(new_n740), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n683), .A2(new_n757), .ZN(new_n992));
  OR3_X1    g0792(.A1(new_n238), .A2(new_n267), .A3(new_n251), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT50), .B1(new_n280), .B2(G50), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n994), .B(new_n267), .C1(new_n342), .C2(new_n258), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n280), .A2(KEYINPUT50), .A3(G50), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n377), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n689), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n690), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n753), .B1(new_n206), .B2(new_n214), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n828), .A2(new_n965), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n280), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n377), .B(new_n974), .C1(new_n1002), .C2(new_n984), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n782), .A2(new_n258), .B1(new_n763), .B2(new_n342), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n761), .A2(new_n202), .B1(new_n784), .B2(new_n834), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1001), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G159), .B2(new_n770), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G317), .A2(new_n796), .B1(new_n831), .B2(G303), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n800), .B2(new_n788), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G322), .B2(new_n770), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT48), .Z(new_n1012));
  OAI22_X1  g0812(.A1(new_n777), .A2(new_n799), .B1(new_n792), .B2(new_n782), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT109), .Z(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n377), .B1(new_n780), .B2(new_n449), .C1(new_n791), .C2(new_n784), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1016), .B2(KEYINPUT49), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1008), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n741), .B1(new_n999), .B2(new_n1000), .C1(new_n1020), .C2(new_n758), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n733), .A2(new_n956), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n691), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n733), .A2(new_n956), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n991), .B1(new_n992), .B2(new_n1021), .C1(new_n1023), .C2(new_n1024), .ZN(G393));
  OAI21_X1  g0825(.A(new_n753), .B1(new_n205), .B2(new_n214), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n248), .B2(new_n963), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1027), .A2(new_n742), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT110), .ZN(new_n1029));
  INV_X1    g0829(.A(G159), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n769), .A2(new_n834), .B1(new_n1030), .B2(new_n761), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT51), .Z(new_n1032));
  AOI22_X1  g0832(.A1(new_n984), .A2(G50), .B1(new_n831), .B2(new_n1002), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT111), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G68), .A2(new_n819), .B1(new_n797), .B2(G143), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1035), .A2(new_n251), .A3(new_n821), .A4(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n777), .A2(new_n258), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1032), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n769), .A2(new_n969), .B1(new_n800), .B2(new_n761), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT52), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n377), .B1(new_n780), .B2(new_n206), .C1(new_n788), .C2(new_n443), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G283), .A2(new_n819), .B1(new_n797), .B2(G322), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n792), .B2(new_n763), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(G116), .C2(new_n828), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1040), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1029), .B1(new_n1047), .B2(new_n758), .C1(new_n929), .C2(new_n757), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n954), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(new_n1049), .B2(new_n739), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1022), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n692), .B1(new_n1051), .B2(new_n954), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1022), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(G390));
  NAND2_X1  g0855(.A1(new_n866), .A2(new_n867), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n720), .B1(new_n718), .B2(KEYINPUT31), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n712), .A2(new_n713), .ZN(new_n1058));
  OAI211_X1 g0858(.A(G330), .B(new_n812), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1059), .A2(new_n864), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n864), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n721), .A2(G330), .A3(new_n812), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1056), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n857), .A2(new_n659), .A3(new_n662), .A4(new_n859), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT103), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n367), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n859), .B1(new_n367), .B2(KEYINPUT103), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1067), .A2(new_n1068), .A3(KEYINPUT113), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT113), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n861), .B2(new_n863), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1059), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n811), .A2(new_n321), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n729), .A2(new_n681), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT112), .B1(new_n1075), .B2(new_n867), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1075), .A2(KEYINPUT112), .A3(new_n867), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1073), .B(new_n1062), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1064), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n432), .A2(new_n721), .A3(G330), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n852), .A2(new_n667), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n901), .B1(new_n868), .B2(new_n890), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1077), .A2(new_n1076), .A3(new_n1072), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n909), .A2(new_n891), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT114), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(KEYINPUT114), .B(new_n1083), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1062), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1063), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1082), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1089), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1075), .A2(new_n867), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT112), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1075), .A2(KEYINPUT112), .A3(new_n867), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1085), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT114), .B1(new_n1101), .B2(new_n1083), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1063), .B1(new_n1093), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1091), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n852), .A2(new_n667), .A3(new_n1080), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n1064), .B2(new_n1078), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1092), .A2(new_n691), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1091), .B1(new_n1109), .B2(new_n1063), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n740), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n901), .A2(new_n749), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n742), .B1(new_n280), .B2(new_n816), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n770), .A2(G283), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n377), .B1(new_n782), .B2(new_n781), .C1(new_n206), .C2(new_n788), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n342), .A2(new_n780), .B1(new_n763), .B2(new_n205), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n761), .A2(new_n449), .B1(new_n784), .B2(new_n792), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1038), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n797), .A2(G125), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1119), .B1(new_n826), .B2(new_n761), .C1(new_n763), .C2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n782), .A2(new_n834), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT53), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n835), .B2(new_n788), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n251), .B1(new_n202), .B2(new_n780), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1121), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n770), .A2(G128), .B1(G159), .B2(new_n828), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1114), .A2(new_n1118), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1112), .B(new_n1113), .C1(new_n758), .C2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1108), .A2(new_n1111), .A3(new_n1130), .ZN(G378));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n297), .A2(new_n369), .ZN(new_n1133));
  XOR2_X1   g0933(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n869), .A2(new_n293), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT116), .Z(new_n1137));
  INV_X1    g0937(.A(new_n1134), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n297), .A2(new_n369), .A3(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1135), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1137), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n904), .B(new_n1142), .C1(new_n915), .C2(new_n913), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1142), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n916), .B2(G330), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n902), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n721), .A2(new_n911), .A3(new_n914), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1147), .A2(new_n887), .B1(new_n912), .B2(KEYINPUT40), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1142), .B1(new_n1148), .B2(new_n904), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n902), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n916), .A2(G330), .A3(new_n1144), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1132), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1090), .A2(new_n1091), .A3(new_n1082), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n1105), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n902), .A2(KEYINPUT118), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1149), .A2(new_n1151), .A3(KEYINPUT118), .A4(new_n902), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1107), .B2(new_n1081), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1155), .B(new_n691), .C1(KEYINPUT57), .C2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n816), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n741), .B1(G50), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(G33), .A2(G41), .ZN(new_n1164));
  AOI211_X1 g0964(.A(G50), .B(new_n1164), .C1(new_n377), .C2(new_n266), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n770), .A2(G116), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n780), .A2(new_n218), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n266), .B(new_n377), .C1(new_n784), .C2(new_n799), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(new_n965), .C2(new_n831), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n258), .A2(new_n782), .B1(new_n761), .B2(new_n206), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G97), .B2(new_n984), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1166), .A2(new_n1169), .A3(new_n982), .A4(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT58), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1165), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT115), .ZN(new_n1175));
  INV_X1    g0975(.A(G124), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1164), .B1(new_n784), .B2(new_n1176), .C1(new_n780), .C2(new_n785), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n763), .A2(new_n835), .ZN(new_n1178));
  INV_X1    g0978(.A(G128), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1179), .A2(new_n761), .B1(new_n782), .B2(new_n1120), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G132), .C2(new_n984), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n770), .A2(G125), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n834), .C2(new_n777), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1177), .B1(new_n1183), .B2(KEYINPUT59), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(KEYINPUT59), .B2(new_n1183), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1175), .B(new_n1185), .C1(new_n1173), .C2(new_n1172), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1163), .B1(new_n1186), .B2(new_n752), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1144), .B2(new_n750), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT117), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1159), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n740), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1161), .A2(new_n1191), .ZN(G375));
  INV_X1    g0992(.A(new_n1079), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1105), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n958), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1195), .A3(new_n1082), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n739), .B(KEYINPUT119), .Z(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1072), .A2(new_n749), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n741), .B1(G68), .B2(new_n1162), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n761), .A2(new_n835), .B1(new_n763), .B2(new_n834), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n782), .A2(new_n1030), .B1(new_n784), .B2(new_n1179), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n788), .A2(new_n1120), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n251), .B1(new_n780), .B2(new_n218), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n202), .B2(new_n777), .C1(new_n826), .C2(new_n769), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n769), .A2(new_n792), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n251), .B(new_n979), .C1(G116), .C2(new_n984), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n761), .A2(new_n799), .B1(new_n763), .B2(new_n206), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n782), .A2(new_n205), .B1(new_n784), .B2(new_n443), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1001), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1206), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1200), .B1(new_n1213), .B2(new_n752), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1079), .A2(new_n1198), .B1(new_n1199), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1196), .A2(new_n1215), .ZN(G381));
  XOR2_X1   g1016(.A(G375), .B(KEYINPUT121), .Z(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(G378), .ZN(new_n1218));
  OR2_X1    g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1219), .A2(KEYINPUT120), .A3(G384), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(G381), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n962), .A2(new_n1054), .A3(new_n989), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT120), .B1(new_n1219), .B2(G384), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1218), .A2(new_n1224), .ZN(G407));
  OAI21_X1  g1025(.A(new_n1218), .B1(new_n674), .B2(new_n1224), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(G213), .ZN(G409));
  NAND2_X1  g1027(.A1(new_n1082), .A2(KEYINPUT60), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1194), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1193), .A2(KEYINPUT60), .A3(new_n1105), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n691), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1215), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n840), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1231), .A2(G384), .A3(new_n1215), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n674), .A2(G213), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(G2897), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(G2897), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1233), .A2(new_n1234), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G378), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1197), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1242));
  OR3_X1    g1042(.A1(new_n1242), .A2(KEYINPUT122), .A3(new_n1189), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT122), .B1(new_n1242), .B2(new_n1189), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1105), .B1(new_n1110), .B2(new_n1079), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1246), .A2(new_n958), .A3(new_n1159), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1241), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1153), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n691), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1107), .A2(new_n1081), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1251), .B2(new_n1190), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G378), .B(new_n1191), .C1(new_n1250), .C2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1236), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  OR3_X1    g1054(.A1(new_n1240), .A2(new_n1254), .A3(KEYINPUT123), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(G393), .B(new_n807), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1054), .B1(new_n962), .B2(new_n989), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1256), .B1(new_n1222), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(G390), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n962), .A2(new_n1054), .A3(new_n989), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1256), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1258), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1236), .B(new_n1235), .C1(new_n1248), .C2(new_n1253), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1265), .B1(new_n1266), .B2(KEYINPUT63), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1235), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1254), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT123), .B1(new_n1240), .B2(new_n1254), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1255), .A2(new_n1267), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1269), .A2(KEYINPUT62), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1266), .A2(new_n1275), .ZN(new_n1276));
  XOR2_X1   g1076(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1240), .B2(new_n1254), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1274), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1273), .B1(new_n1279), .B2(new_n1263), .ZN(G405));
  NOR2_X1   g1080(.A1(new_n1263), .A2(KEYINPUT126), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1258), .A2(new_n1262), .A3(KEYINPUT126), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1253), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1161), .B2(new_n1191), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1233), .A2(KEYINPUT125), .A3(new_n1234), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1284), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1288), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1283), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G375), .A2(new_n1241), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n1253), .A3(new_n1288), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1258), .A2(new_n1262), .A3(KEYINPUT126), .ZN(new_n1295));
  AND4_X1   g1095(.A1(new_n1283), .A2(new_n1294), .A3(new_n1291), .A4(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1282), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1291), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT127), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1289), .A2(new_n1283), .A3(new_n1291), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1301), .A3(new_n1281), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1297), .A2(new_n1302), .ZN(G402));
endmodule


