

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U556 ( .A1(n693), .A2(n692), .ZN(n694) );
  AND2_X1 U557 ( .A1(n575), .A2(G2105), .ZN(n927) );
  NOR2_X2 U558 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U559 ( .A1(n550), .A2(KEYINPUT109), .ZN(n549) );
  AND2_X1 U560 ( .A1(n546), .A2(n540), .ZN(n539) );
  AND2_X1 U561 ( .A1(n695), .A2(n696), .ZN(n536) );
  NOR2_X1 U562 ( .A1(n666), .A2(n981), .ZN(n668) );
  NAND2_X2 U563 ( .A1(n569), .A2(n566), .ZN(n580) );
  NAND2_X1 U564 ( .A1(n559), .A2(n556), .ZN(n683) );
  NAND2_X1 U565 ( .A1(n558), .A2(n557), .ZN(n556) );
  AND2_X1 U566 ( .A1(n561), .A2(n560), .ZN(n559) );
  NOR2_X1 U567 ( .A1(n1021), .A2(n563), .ZN(n557) );
  NAND2_X1 U568 ( .A1(n562), .A2(n1012), .ZN(n564) );
  INV_X1 U569 ( .A(n683), .ZN(n562) );
  NAND2_X1 U570 ( .A1(n534), .A2(n531), .ZN(n711) );
  XNOR2_X1 U571 ( .A(n533), .B(n532), .ZN(n531) );
  XNOR2_X1 U572 ( .A(n706), .B(KEYINPUT31), .ZN(n532) );
  XNOR2_X1 U573 ( .A(n654), .B(KEYINPUT64), .ZN(n666) );
  NAND2_X1 U574 ( .A1(KEYINPUT33), .A2(n544), .ZN(n542) );
  AND2_X1 U575 ( .A1(n730), .A2(KEYINPUT105), .ZN(n547) );
  NAND2_X1 U576 ( .A1(n545), .A2(n544), .ZN(n543) );
  INV_X1 U577 ( .A(n571), .ZN(n545) );
  INV_X1 U578 ( .A(KEYINPUT105), .ZN(n544) );
  INV_X1 U579 ( .A(n784), .ZN(n552) );
  AND2_X1 U580 ( .A1(n568), .A2(n567), .ZN(n566) );
  NAND2_X1 U581 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n568) );
  XNOR2_X1 U582 ( .A(n587), .B(n586), .ZN(n588) );
  INV_X1 U583 ( .A(KEYINPUT68), .ZN(n586) );
  XNOR2_X1 U584 ( .A(n584), .B(KEYINPUT23), .ZN(n589) );
  NAND2_X1 U585 ( .A1(n583), .A2(G101), .ZN(n584) );
  INV_X1 U586 ( .A(KEYINPUT65), .ZN(n563) );
  NAND2_X1 U587 ( .A1(n1021), .A2(n563), .ZN(n560) );
  NAND2_X1 U588 ( .A1(n564), .A2(n682), .ZN(n685) );
  NAND2_X1 U589 ( .A1(n526), .A2(n524), .ZN(n533) );
  XNOR2_X1 U590 ( .A(n722), .B(n721), .ZN(n736) );
  NAND2_X1 U591 ( .A1(n543), .A2(n541), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n731), .A2(n547), .ZN(n546) );
  NAND2_X1 U593 ( .A1(n571), .A2(n542), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n538), .A2(n528), .ZN(n537) );
  NOR2_X1 U595 ( .A1(KEYINPUT17), .A2(G2104), .ZN(n565) );
  NAND2_X1 U596 ( .A1(G2105), .A2(KEYINPUT17), .ZN(n567) );
  AND2_X1 U597 ( .A1(n572), .A2(G2104), .ZN(n583) );
  AND2_X1 U598 ( .A1(n784), .A2(n786), .ZN(n554) );
  NAND2_X1 U599 ( .A1(n552), .A2(KEYINPUT109), .ZN(n551) );
  NOR2_X1 U600 ( .A1(G651), .A2(n627), .ZN(n834) );
  AND2_X1 U601 ( .A1(n582), .A2(n581), .ZN(n591) );
  XNOR2_X1 U602 ( .A(KEYINPUT100), .B(n705), .ZN(n524) );
  AND2_X1 U603 ( .A1(n553), .A2(n530), .ZN(n525) );
  AND2_X2 U604 ( .A1(G2105), .A2(G2104), .ZN(n585) );
  OR2_X1 U605 ( .A1(G168), .A2(n703), .ZN(n526) );
  OR2_X1 U606 ( .A1(G301), .A2(n704), .ZN(n527) );
  AND2_X1 U607 ( .A1(n571), .A2(n544), .ZN(n528) );
  OR2_X1 U608 ( .A1(n726), .A2(n725), .ZN(n529) );
  AND2_X1 U609 ( .A1(n800), .A2(n551), .ZN(n530) );
  NAND2_X1 U610 ( .A1(n535), .A2(n527), .ZN(n534) );
  XNOR2_X1 U611 ( .A(n536), .B(KEYINPUT29), .ZN(n535) );
  NAND2_X1 U612 ( .A1(n539), .A2(n537), .ZN(n548) );
  INV_X1 U613 ( .A(n731), .ZN(n538) );
  NOR2_X2 U614 ( .A1(n548), .A2(n741), .ZN(n742) );
  NAND2_X1 U615 ( .A1(n525), .A2(n549), .ZN(n555) );
  INV_X1 U616 ( .A(n785), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n785), .A2(n554), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n555), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U619 ( .A(n671), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n671), .A2(n563), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n565), .A2(n572), .ZN(n569) );
  NAND2_X1 U622 ( .A1(n580), .A2(G137), .ZN(n582) );
  XNOR2_X2 U623 ( .A(n592), .B(KEYINPUT67), .ZN(G160) );
  OR2_X1 U624 ( .A1(n732), .A2(n713), .ZN(n570) );
  AND2_X1 U625 ( .A1(n1003), .A2(n570), .ZN(n571) );
  INV_X1 U626 ( .A(n713), .ZN(n728) );
  INV_X1 U627 ( .A(G2105), .ZN(n572) );
  INV_X1 U628 ( .A(G2104), .ZN(n575) );
  INV_X1 U629 ( .A(KEYINPUT109), .ZN(n786) );
  NAND2_X1 U630 ( .A1(G138), .A2(n580), .ZN(n574) );
  BUF_X1 U631 ( .A(n583), .Z(n923) );
  NAND2_X1 U632 ( .A1(G102), .A2(n923), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U634 ( .A1(G126), .A2(n927), .ZN(n577) );
  NAND2_X1 U635 ( .A1(G114), .A2(n585), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U637 ( .A1(n579), .A2(n578), .ZN(G164) );
  NAND2_X1 U638 ( .A1(G125), .A2(n927), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G113), .A2(n585), .ZN(n587) );
  NAND2_X1 U640 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U641 ( .A(G543), .B(KEYINPUT0), .Z(n627) );
  NAND2_X1 U642 ( .A1(G53), .A2(n834), .ZN(n602) );
  INV_X1 U643 ( .A(G651), .ZN(n597) );
  NOR2_X1 U644 ( .A1(G543), .A2(n597), .ZN(n593) );
  XOR2_X1 U645 ( .A(KEYINPUT1), .B(n593), .Z(n830) );
  NAND2_X1 U646 ( .A1(n830), .A2(G65), .ZN(n596) );
  NOR2_X1 U647 ( .A1(G543), .A2(G651), .ZN(n594) );
  XNOR2_X1 U648 ( .A(n594), .B(KEYINPUT66), .ZN(n828) );
  NAND2_X1 U649 ( .A1(G91), .A2(n828), .ZN(n595) );
  NAND2_X1 U650 ( .A1(n596), .A2(n595), .ZN(n600) );
  NOR2_X1 U651 ( .A1(n627), .A2(n597), .ZN(n833) );
  NAND2_X1 U652 ( .A1(G78), .A2(n833), .ZN(n598) );
  XNOR2_X1 U653 ( .A(KEYINPUT71), .B(n598), .ZN(n599) );
  NOR2_X1 U654 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U655 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U656 ( .A(n603), .B(KEYINPUT72), .ZN(G299) );
  NAND2_X1 U657 ( .A1(n833), .A2(G77), .ZN(n604) );
  XNOR2_X1 U658 ( .A(n604), .B(KEYINPUT70), .ZN(n606) );
  NAND2_X1 U659 ( .A1(G90), .A2(n828), .ZN(n605) );
  NAND2_X1 U660 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U661 ( .A(KEYINPUT9), .B(n607), .ZN(n611) );
  NAND2_X1 U662 ( .A1(G64), .A2(n830), .ZN(n609) );
  NAND2_X1 U663 ( .A1(G52), .A2(n834), .ZN(n608) );
  AND2_X1 U664 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U665 ( .A1(n611), .A2(n610), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G89), .A2(n828), .ZN(n612) );
  XNOR2_X1 U667 ( .A(n612), .B(KEYINPUT4), .ZN(n614) );
  NAND2_X1 U668 ( .A1(G76), .A2(n833), .ZN(n613) );
  NAND2_X1 U669 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U670 ( .A(n615), .B(KEYINPUT5), .ZN(n620) );
  NAND2_X1 U671 ( .A1(G63), .A2(n830), .ZN(n617) );
  NAND2_X1 U672 ( .A1(G51), .A2(n834), .ZN(n616) );
  NAND2_X1 U673 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U674 ( .A(KEYINPUT6), .B(n618), .Z(n619) );
  NAND2_X1 U675 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U676 ( .A(n621), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U677 ( .A1(G651), .A2(G74), .ZN(n622) );
  XOR2_X1 U678 ( .A(KEYINPUT79), .B(n622), .Z(n624) );
  NAND2_X1 U679 ( .A1(n834), .A2(G49), .ZN(n623) );
  NAND2_X1 U680 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U681 ( .A(KEYINPUT80), .B(n625), .ZN(n626) );
  NOR2_X1 U682 ( .A1(n830), .A2(n626), .ZN(n629) );
  NAND2_X1 U683 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U684 ( .A1(n629), .A2(n628), .ZN(G288) );
  XOR2_X1 U685 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U686 ( .A1(n833), .A2(G75), .ZN(n631) );
  NAND2_X1 U687 ( .A1(G88), .A2(n828), .ZN(n630) );
  NAND2_X1 U688 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U689 ( .A1(G62), .A2(n830), .ZN(n633) );
  NAND2_X1 U690 ( .A1(G50), .A2(n834), .ZN(n632) );
  NAND2_X1 U691 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U692 ( .A1(n635), .A2(n634), .ZN(G166) );
  INV_X1 U693 ( .A(G166), .ZN(G303) );
  NAND2_X1 U694 ( .A1(n830), .A2(G61), .ZN(n637) );
  NAND2_X1 U695 ( .A1(G86), .A2(n828), .ZN(n636) );
  NAND2_X1 U696 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U697 ( .A1(n834), .A2(G48), .ZN(n638) );
  XOR2_X1 U698 ( .A(KEYINPUT82), .B(n638), .Z(n639) );
  NOR2_X1 U699 ( .A1(n640), .A2(n639), .ZN(n644) );
  XOR2_X1 U700 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n642) );
  NAND2_X1 U701 ( .A1(G73), .A2(n833), .ZN(n641) );
  XNOR2_X1 U702 ( .A(n642), .B(n641), .ZN(n643) );
  NAND2_X1 U703 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U704 ( .A(KEYINPUT83), .B(n645), .Z(G305) );
  NAND2_X1 U705 ( .A1(G72), .A2(n833), .ZN(n647) );
  NAND2_X1 U706 ( .A1(G47), .A2(n834), .ZN(n646) );
  NAND2_X1 U707 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U708 ( .A1(G85), .A2(n828), .ZN(n648) );
  XNOR2_X1 U709 ( .A(KEYINPUT69), .B(n648), .ZN(n649) );
  NOR2_X1 U710 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U711 ( .A1(n830), .A2(G60), .ZN(n651) );
  NAND2_X1 U712 ( .A1(n652), .A2(n651), .ZN(G290) );
  NOR2_X1 U713 ( .A1(G164), .A2(G1384), .ZN(n749) );
  NAND2_X1 U714 ( .A1(G160), .A2(G40), .ZN(n748) );
  XNOR2_X1 U715 ( .A(n748), .B(KEYINPUT93), .ZN(n653) );
  NAND2_X1 U716 ( .A1(n749), .A2(n653), .ZN(n654) );
  INV_X1 U717 ( .A(n666), .ZN(n655) );
  INV_X2 U718 ( .A(n655), .ZN(n697) );
  NOR2_X1 U719 ( .A1(n697), .A2(G2084), .ZN(n700) );
  NAND2_X1 U720 ( .A1(n700), .A2(G8), .ZN(n710) );
  NAND2_X1 U721 ( .A1(n697), .A2(G8), .ZN(n713) );
  NOR2_X1 U722 ( .A1(G1966), .A2(n713), .ZN(n708) );
  NAND2_X1 U723 ( .A1(G81), .A2(n828), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n656), .B(KEYINPUT12), .ZN(n658) );
  NAND2_X1 U725 ( .A1(G68), .A2(n833), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT13), .B(n659), .Z(n663) );
  NAND2_X1 U728 ( .A1(G56), .A2(n830), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n660), .B(KEYINPUT73), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT14), .ZN(n662) );
  NOR2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n834), .A2(G43), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n1021) );
  XNOR2_X1 U734 ( .A(G1996), .B(KEYINPUT97), .ZN(n981) );
  XOR2_X1 U735 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n697), .A2(G1341), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n833), .A2(G79), .ZN(n673) );
  NAND2_X1 U740 ( .A1(G92), .A2(n828), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n677) );
  NAND2_X1 U742 ( .A1(G66), .A2(n830), .ZN(n675) );
  NAND2_X1 U743 ( .A1(G54), .A2(n834), .ZN(n674) );
  NAND2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U746 ( .A(KEYINPUT15), .B(n678), .Z(n1012) );
  INV_X1 U747 ( .A(n1012), .ZN(n813) );
  INV_X1 U748 ( .A(G2067), .ZN(n760) );
  NOR2_X1 U749 ( .A1(n697), .A2(n760), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n679), .B(KEYINPUT99), .ZN(n681) );
  NAND2_X1 U751 ( .A1(n697), .A2(G1348), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U753 ( .A1(n813), .A2(n683), .ZN(n684) );
  NAND2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n691) );
  XOR2_X1 U755 ( .A(KEYINPUT95), .B(KEYINPUT27), .Z(n687) );
  NAND2_X1 U756 ( .A1(G2072), .A2(n655), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n687), .B(n686), .ZN(n689) );
  XOR2_X1 U758 ( .A(G1956), .B(KEYINPUT96), .Z(n1044) );
  NOR2_X1 U759 ( .A1(n1044), .A2(n655), .ZN(n688) );
  NOR2_X1 U760 ( .A1(n689), .A2(n688), .ZN(n693) );
  INV_X1 U761 ( .A(G299), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n690) );
  NAND2_X1 U763 ( .A1(n691), .A2(n690), .ZN(n696) );
  XOR2_X1 U764 ( .A(n694), .B(KEYINPUT28), .Z(n695) );
  XOR2_X1 U765 ( .A(G2078), .B(KEYINPUT25), .Z(n983) );
  NAND2_X1 U766 ( .A1(n983), .A2(n655), .ZN(n699) );
  NAND2_X1 U767 ( .A1(n697), .A2(G1961), .ZN(n698) );
  NAND2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n704) );
  XOR2_X1 U769 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n706) );
  NOR2_X1 U770 ( .A1(n708), .A2(n700), .ZN(n701) );
  NAND2_X1 U771 ( .A1(G8), .A2(n701), .ZN(n702) );
  XNOR2_X1 U772 ( .A(KEYINPUT30), .B(n702), .ZN(n703) );
  NAND2_X1 U773 ( .A1(G301), .A2(n704), .ZN(n705) );
  INV_X1 U774 ( .A(n711), .ZN(n707) );
  NOR2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n735) );
  NAND2_X1 U777 ( .A1(G1976), .A2(G288), .ZN(n1007) );
  AND2_X1 U778 ( .A1(n735), .A2(n1007), .ZN(n723) );
  NAND2_X1 U779 ( .A1(n711), .A2(G286), .ZN(n720) );
  INV_X1 U780 ( .A(G8), .ZN(n718) );
  NOR2_X1 U781 ( .A1(n697), .A2(G2090), .ZN(n712) );
  XNOR2_X1 U782 ( .A(KEYINPUT103), .B(n712), .ZN(n716) );
  NOR2_X1 U783 ( .A1(G1971), .A2(n713), .ZN(n714) );
  NOR2_X1 U784 ( .A1(G166), .A2(n714), .ZN(n715) );
  NAND2_X1 U785 ( .A1(n716), .A2(n715), .ZN(n717) );
  OR2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U787 ( .A1(n720), .A2(n719), .ZN(n722) );
  XOR2_X1 U788 ( .A(KEYINPUT104), .B(KEYINPUT32), .Z(n721) );
  NAND2_X1 U789 ( .A1(n723), .A2(n736), .ZN(n727) );
  INV_X1 U790 ( .A(n1007), .ZN(n726) );
  NOR2_X1 U791 ( .A1(G1976), .A2(G288), .ZN(n1006) );
  NOR2_X1 U792 ( .A1(G1971), .A2(G303), .ZN(n724) );
  NOR2_X1 U793 ( .A1(n1006), .A2(n724), .ZN(n725) );
  NAND2_X1 U794 ( .A1(n727), .A2(n529), .ZN(n729) );
  NAND2_X1 U795 ( .A1(n729), .A2(n728), .ZN(n731) );
  INV_X1 U796 ( .A(KEYINPUT33), .ZN(n730) );
  XOR2_X1 U797 ( .A(G1981), .B(G305), .Z(n1003) );
  NAND2_X1 U798 ( .A1(n1006), .A2(KEYINPUT33), .ZN(n732) );
  NOR2_X1 U799 ( .A1(G2090), .A2(G303), .ZN(n733) );
  NAND2_X1 U800 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U801 ( .A(n734), .B(KEYINPUT106), .ZN(n738) );
  NAND2_X1 U802 ( .A1(n735), .A2(n736), .ZN(n737) );
  NAND2_X1 U803 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U804 ( .A1(n739), .A2(n713), .ZN(n740) );
  XNOR2_X1 U805 ( .A(KEYINPUT107), .B(n740), .ZN(n741) );
  XNOR2_X1 U806 ( .A(n742), .B(KEYINPUT108), .ZN(n747) );
  NOR2_X1 U807 ( .A1(G1981), .A2(G305), .ZN(n743) );
  XOR2_X1 U808 ( .A(n743), .B(KEYINPUT24), .Z(n744) );
  NOR2_X1 U809 ( .A1(n713), .A2(n744), .ZN(n745) );
  XOR2_X1 U810 ( .A(KEYINPUT94), .B(n745), .Z(n746) );
  NAND2_X1 U811 ( .A1(n747), .A2(n746), .ZN(n785) );
  NOR2_X1 U812 ( .A1(n749), .A2(n748), .ZN(n798) );
  INV_X1 U813 ( .A(n798), .ZN(n761) );
  NAND2_X1 U814 ( .A1(G128), .A2(n927), .ZN(n751) );
  NAND2_X1 U815 ( .A1(G116), .A2(n585), .ZN(n750) );
  NAND2_X1 U816 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U817 ( .A(n752), .B(KEYINPUT35), .ZN(n758) );
  NAND2_X1 U818 ( .A1(n580), .A2(G140), .ZN(n753) );
  XOR2_X1 U819 ( .A(KEYINPUT87), .B(n753), .Z(n755) );
  NAND2_X1 U820 ( .A1(n923), .A2(G104), .ZN(n754) );
  NAND2_X1 U821 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U822 ( .A(KEYINPUT34), .B(n756), .Z(n757) );
  NAND2_X1 U823 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U824 ( .A(n759), .B(KEYINPUT36), .ZN(n939) );
  XNOR2_X1 U825 ( .A(n760), .B(KEYINPUT37), .ZN(n795) );
  NAND2_X1 U826 ( .A1(n939), .A2(n795), .ZN(n972) );
  NOR2_X1 U827 ( .A1(n761), .A2(n972), .ZN(n792) );
  XOR2_X1 U828 ( .A(KEYINPUT38), .B(KEYINPUT88), .Z(n763) );
  NAND2_X1 U829 ( .A1(G105), .A2(n923), .ZN(n762) );
  XNOR2_X1 U830 ( .A(n763), .B(n762), .ZN(n767) );
  NAND2_X1 U831 ( .A1(G129), .A2(n927), .ZN(n765) );
  NAND2_X1 U832 ( .A1(G117), .A2(n585), .ZN(n764) );
  NAND2_X1 U833 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U834 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U835 ( .A(KEYINPUT89), .B(n768), .Z(n770) );
  NAND2_X1 U836 ( .A1(n580), .A2(G141), .ZN(n769) );
  NAND2_X1 U837 ( .A1(n770), .A2(n769), .ZN(n933) );
  NAND2_X1 U838 ( .A1(G1996), .A2(n933), .ZN(n771) );
  XNOR2_X1 U839 ( .A(n771), .B(KEYINPUT90), .ZN(n779) );
  NAND2_X1 U840 ( .A1(G119), .A2(n927), .ZN(n773) );
  NAND2_X1 U841 ( .A1(G107), .A2(n585), .ZN(n772) );
  NAND2_X1 U842 ( .A1(n773), .A2(n772), .ZN(n777) );
  NAND2_X1 U843 ( .A1(G131), .A2(n580), .ZN(n775) );
  NAND2_X1 U844 ( .A1(G95), .A2(n923), .ZN(n774) );
  NAND2_X1 U845 ( .A1(n775), .A2(n774), .ZN(n776) );
  OR2_X1 U846 ( .A1(n777), .A2(n776), .ZN(n919) );
  NAND2_X1 U847 ( .A1(G1991), .A2(n919), .ZN(n778) );
  NAND2_X1 U848 ( .A1(n779), .A2(n778), .ZN(n954) );
  NAND2_X1 U849 ( .A1(n798), .A2(n954), .ZN(n780) );
  XNOR2_X1 U850 ( .A(KEYINPUT91), .B(n780), .ZN(n789) );
  NOR2_X1 U851 ( .A1(n792), .A2(n789), .ZN(n781) );
  XNOR2_X1 U852 ( .A(KEYINPUT92), .B(n781), .ZN(n783) );
  XNOR2_X1 U853 ( .A(G1986), .B(G290), .ZN(n1011) );
  NAND2_X1 U854 ( .A1(n798), .A2(n1011), .ZN(n782) );
  AND2_X1 U855 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U856 ( .A1(G1996), .A2(n933), .ZN(n957) );
  NOR2_X1 U857 ( .A1(G1991), .A2(n919), .ZN(n965) );
  NOR2_X1 U858 ( .A1(G1986), .A2(G290), .ZN(n787) );
  NOR2_X1 U859 ( .A1(n965), .A2(n787), .ZN(n788) );
  NOR2_X1 U860 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U861 ( .A1(n957), .A2(n790), .ZN(n791) );
  XNOR2_X1 U862 ( .A(KEYINPUT39), .B(n791), .ZN(n794) );
  INV_X1 U863 ( .A(n792), .ZN(n793) );
  NAND2_X1 U864 ( .A1(n794), .A2(n793), .ZN(n797) );
  NOR2_X1 U865 ( .A1(n939), .A2(n795), .ZN(n955) );
  INV_X1 U866 ( .A(n955), .ZN(n796) );
  NAND2_X1 U867 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U868 ( .A1(n799), .A2(n798), .ZN(n800) );
  AND2_X1 U869 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U870 ( .A1(G123), .A2(n927), .ZN(n801) );
  XNOR2_X1 U871 ( .A(n801), .B(KEYINPUT18), .ZN(n808) );
  NAND2_X1 U872 ( .A1(G135), .A2(n580), .ZN(n803) );
  NAND2_X1 U873 ( .A1(G111), .A2(n585), .ZN(n802) );
  NAND2_X1 U874 ( .A1(n803), .A2(n802), .ZN(n806) );
  NAND2_X1 U875 ( .A1(G99), .A2(n923), .ZN(n804) );
  XNOR2_X1 U876 ( .A(KEYINPUT77), .B(n804), .ZN(n805) );
  NOR2_X1 U877 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U878 ( .A1(n808), .A2(n807), .ZN(n962) );
  XNOR2_X1 U879 ( .A(G2096), .B(n962), .ZN(n809) );
  OR2_X1 U880 ( .A1(G2100), .A2(n809), .ZN(G156) );
  INV_X1 U881 ( .A(G57), .ZN(G237) );
  NAND2_X1 U882 ( .A1(G7), .A2(G661), .ZN(n810) );
  XNOR2_X1 U883 ( .A(n810), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U884 ( .A(G223), .ZN(n865) );
  NAND2_X1 U885 ( .A1(n865), .A2(G567), .ZN(n811) );
  XOR2_X1 U886 ( .A(KEYINPUT11), .B(n811), .Z(G234) );
  INV_X1 U887 ( .A(G860), .ZN(n827) );
  OR2_X1 U888 ( .A1(n1021), .A2(n827), .ZN(G153) );
  NAND2_X1 U889 ( .A1(G301), .A2(G868), .ZN(n812) );
  XNOR2_X1 U890 ( .A(n812), .B(KEYINPUT74), .ZN(n815) );
  INV_X1 U891 ( .A(G868), .ZN(n817) );
  NAND2_X1 U892 ( .A1(n817), .A2(n813), .ZN(n814) );
  NAND2_X1 U893 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U894 ( .A(KEYINPUT75), .B(n816), .Z(G284) );
  NOR2_X1 U895 ( .A1(G299), .A2(G868), .ZN(n819) );
  NOR2_X1 U896 ( .A1(G286), .A2(n817), .ZN(n818) );
  NOR2_X1 U897 ( .A1(n819), .A2(n818), .ZN(G297) );
  NAND2_X1 U898 ( .A1(n827), .A2(G559), .ZN(n820) );
  NAND2_X1 U899 ( .A1(n820), .A2(n1012), .ZN(n821) );
  XNOR2_X1 U900 ( .A(n821), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U901 ( .A1(G868), .A2(n1021), .ZN(n824) );
  NAND2_X1 U902 ( .A1(G868), .A2(n1012), .ZN(n822) );
  NOR2_X1 U903 ( .A1(G559), .A2(n822), .ZN(n823) );
  NOR2_X1 U904 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U905 ( .A(KEYINPUT76), .B(n825), .ZN(G282) );
  NAND2_X1 U906 ( .A1(G559), .A2(n1012), .ZN(n826) );
  XOR2_X1 U907 ( .A(n1021), .B(n826), .Z(n846) );
  NAND2_X1 U908 ( .A1(n827), .A2(n846), .ZN(n839) );
  NAND2_X1 U909 ( .A1(G93), .A2(n828), .ZN(n829) );
  XNOR2_X1 U910 ( .A(n829), .B(KEYINPUT78), .ZN(n832) );
  NAND2_X1 U911 ( .A1(G67), .A2(n830), .ZN(n831) );
  NAND2_X1 U912 ( .A1(n832), .A2(n831), .ZN(n838) );
  NAND2_X1 U913 ( .A1(G80), .A2(n833), .ZN(n836) );
  NAND2_X1 U914 ( .A1(G55), .A2(n834), .ZN(n835) );
  NAND2_X1 U915 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U916 ( .A1(n838), .A2(n837), .ZN(n848) );
  XOR2_X1 U917 ( .A(n839), .B(n848), .Z(G145) );
  XNOR2_X1 U918 ( .A(G299), .B(G305), .ZN(n845) );
  XNOR2_X1 U919 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n841) );
  XNOR2_X1 U920 ( .A(G288), .B(G166), .ZN(n840) );
  XNOR2_X1 U921 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U922 ( .A(n848), .B(n842), .ZN(n843) );
  XNOR2_X1 U923 ( .A(n843), .B(G290), .ZN(n844) );
  XNOR2_X1 U924 ( .A(n845), .B(n844), .ZN(n942) );
  XNOR2_X1 U925 ( .A(n846), .B(n942), .ZN(n847) );
  NAND2_X1 U926 ( .A1(n847), .A2(G868), .ZN(n850) );
  OR2_X1 U927 ( .A1(G868), .A2(n848), .ZN(n849) );
  NAND2_X1 U928 ( .A1(n850), .A2(n849), .ZN(G295) );
  NAND2_X1 U929 ( .A1(G2084), .A2(G2078), .ZN(n851) );
  XOR2_X1 U930 ( .A(KEYINPUT20), .B(n851), .Z(n852) );
  NAND2_X1 U931 ( .A1(G2090), .A2(n852), .ZN(n853) );
  XNOR2_X1 U932 ( .A(KEYINPUT21), .B(n853), .ZN(n854) );
  NAND2_X1 U933 ( .A1(n854), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U934 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U935 ( .A1(G120), .A2(G69), .ZN(n855) );
  NOR2_X1 U936 ( .A1(G237), .A2(n855), .ZN(n856) );
  XNOR2_X1 U937 ( .A(KEYINPUT86), .B(n856), .ZN(n857) );
  NAND2_X1 U938 ( .A1(n857), .A2(G108), .ZN(n869) );
  NAND2_X1 U939 ( .A1(n869), .A2(G567), .ZN(n863) );
  XOR2_X1 U940 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n859) );
  NAND2_X1 U941 ( .A1(G132), .A2(G82), .ZN(n858) );
  XNOR2_X1 U942 ( .A(n859), .B(n858), .ZN(n860) );
  NOR2_X1 U943 ( .A1(n860), .A2(G218), .ZN(n861) );
  NAND2_X1 U944 ( .A1(G96), .A2(n861), .ZN(n870) );
  NAND2_X1 U945 ( .A1(n870), .A2(G2106), .ZN(n862) );
  NAND2_X1 U946 ( .A1(n863), .A2(n862), .ZN(n953) );
  NAND2_X1 U947 ( .A1(G661), .A2(G483), .ZN(n864) );
  NOR2_X1 U948 ( .A1(n953), .A2(n864), .ZN(n868) );
  NAND2_X1 U949 ( .A1(n868), .A2(G36), .ZN(G176) );
  NAND2_X1 U950 ( .A1(G2106), .A2(n865), .ZN(G217) );
  AND2_X1 U951 ( .A1(G15), .A2(G2), .ZN(n866) );
  NAND2_X1 U952 ( .A1(G661), .A2(n866), .ZN(G259) );
  NAND2_X1 U953 ( .A1(G3), .A2(G1), .ZN(n867) );
  NAND2_X1 U954 ( .A1(n868), .A2(n867), .ZN(G188) );
  INV_X1 U956 ( .A(G132), .ZN(G219) );
  INV_X1 U957 ( .A(G120), .ZN(G236) );
  INV_X1 U958 ( .A(G108), .ZN(G238) );
  INV_X1 U959 ( .A(G96), .ZN(G221) );
  INV_X1 U960 ( .A(G82), .ZN(G220) );
  INV_X1 U961 ( .A(G69), .ZN(G235) );
  NOR2_X1 U962 ( .A1(n870), .A2(n869), .ZN(G325) );
  INV_X1 U963 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U964 ( .A(G1341), .B(G2454), .ZN(n871) );
  XNOR2_X1 U965 ( .A(n871), .B(G2430), .ZN(n872) );
  XNOR2_X1 U966 ( .A(n872), .B(G1348), .ZN(n878) );
  XOR2_X1 U967 ( .A(G2443), .B(G2427), .Z(n874) );
  XNOR2_X1 U968 ( .A(G2438), .B(G2446), .ZN(n873) );
  XNOR2_X1 U969 ( .A(n874), .B(n873), .ZN(n876) );
  XOR2_X1 U970 ( .A(G2451), .B(G2435), .Z(n875) );
  XNOR2_X1 U971 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U972 ( .A(n878), .B(n877), .ZN(n879) );
  NAND2_X1 U973 ( .A1(n879), .A2(G14), .ZN(n880) );
  XOR2_X1 U974 ( .A(KEYINPUT110), .B(n880), .Z(G401) );
  XOR2_X1 U975 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n882) );
  XNOR2_X1 U976 ( .A(G2678), .B(KEYINPUT111), .ZN(n881) );
  XNOR2_X1 U977 ( .A(n882), .B(n881), .ZN(n886) );
  XOR2_X1 U978 ( .A(KEYINPUT42), .B(G2072), .Z(n884) );
  XNOR2_X1 U979 ( .A(G2067), .B(G2090), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U981 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U982 ( .A(G2096), .B(G2100), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n888), .B(n887), .ZN(n890) );
  XOR2_X1 U984 ( .A(G2084), .B(G2078), .Z(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(G227) );
  XOR2_X1 U986 ( .A(G1956), .B(G1971), .Z(n892) );
  XNOR2_X1 U987 ( .A(G1986), .B(G1976), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U989 ( .A(G1966), .B(G1981), .Z(n894) );
  XNOR2_X1 U990 ( .A(G1996), .B(G1991), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U992 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U993 ( .A(KEYINPUT113), .B(G2474), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n900) );
  XOR2_X1 U995 ( .A(G1961), .B(KEYINPUT41), .Z(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(G229) );
  NAND2_X1 U997 ( .A1(n927), .A2(G124), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(KEYINPUT44), .ZN(n903) );
  NAND2_X1 U999 ( .A1(G112), .A2(n585), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(G136), .A2(n580), .ZN(n905) );
  NAND2_X1 U1002 ( .A1(G100), .A2(n923), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(G162) );
  XNOR2_X1 U1005 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n962), .B(KEYINPUT117), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n922) );
  NAND2_X1 U1008 ( .A1(G142), .A2(n580), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(G106), .A2(n923), .ZN(n910) );
  NAND2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1011 ( .A(KEYINPUT45), .B(n912), .Z(n918) );
  NAND2_X1 U1012 ( .A1(n585), .A2(G118), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n913), .B(KEYINPUT114), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(G130), .A2(n927), .ZN(n914) );
  NAND2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1016 ( .A(n916), .B(KEYINPUT115), .Z(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n922), .B(n921), .ZN(n935) );
  NAND2_X1 U1020 ( .A1(G139), .A2(n580), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(G103), .A2(n923), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(KEYINPUT116), .B(n926), .ZN(n932) );
  NAND2_X1 U1024 ( .A1(G127), .A2(n927), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(G115), .A2(n585), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT47), .B(n930), .Z(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n968) );
  XNOR2_X1 U1029 ( .A(n933), .B(n968), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(n935), .B(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(n936), .B(G162), .Z(n938) );
  XNOR2_X1 U1032 ( .A(G164), .B(G160), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(n938), .B(n937), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(n940), .B(n939), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(G37), .A2(n941), .ZN(G395) );
  INV_X1 U1036 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1037 ( .A(KEYINPUT118), .B(n942), .Z(n944) );
  XNOR2_X1 U1038 ( .A(G171), .B(n1012), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n944), .B(n943), .ZN(n946) );
  XOR2_X1 U1040 ( .A(n1021), .B(G286), .Z(n945) );
  XNOR2_X1 U1041 ( .A(n946), .B(n945), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(G37), .A2(n947), .ZN(G397) );
  OR2_X1 U1043 ( .A1(n953), .A2(G401), .ZN(n950) );
  NOR2_X1 U1044 ( .A1(G227), .A2(G229), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT49), .B(n948), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(G395), .A2(G397), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(G225) );
  INV_X1 U1049 ( .A(G225), .ZN(G308) );
  INV_X1 U1050 ( .A(n953), .ZN(G319) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n967) );
  XOR2_X1 U1052 ( .A(G160), .B(G2084), .Z(n961) );
  XOR2_X1 U1053 ( .A(G2090), .B(G162), .Z(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1055 ( .A(KEYINPUT119), .B(n958), .Z(n959) );
  XNOR2_X1 U1056 ( .A(KEYINPUT51), .B(n959), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n975) );
  XOR2_X1 U1061 ( .A(G2072), .B(n968), .Z(n970) );
  XOR2_X1 U1062 ( .A(G164), .B(G2078), .Z(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n971), .B(KEYINPUT50), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(KEYINPUT52), .B(n976), .ZN(n977) );
  INV_X1 U1068 ( .A(KEYINPUT55), .ZN(n999) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n999), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n978), .A2(G29), .ZN(n1061) );
  XNOR2_X1 U1071 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(n979), .B(G34), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G2084), .B(n980), .ZN(n997) );
  XNOR2_X1 U1074 ( .A(G2090), .B(G35), .ZN(n995) );
  XNOR2_X1 U1075 ( .A(G32), .B(n981), .ZN(n987) );
  XOR2_X1 U1076 ( .A(G1991), .B(G25), .Z(n982) );
  NAND2_X1 U1077 ( .A1(n982), .A2(G28), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(G27), .B(n983), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G2067), .B(G26), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(G2072), .B(G33), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1084 ( .A(KEYINPUT120), .B(n990), .Z(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(KEYINPUT53), .B(n993), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n999), .B(n998), .ZN(n1001) );
  INV_X1 U1090 ( .A(G29), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(G11), .A2(n1002), .ZN(n1059) );
  XNOR2_X1 U1093 ( .A(G16), .B(KEYINPUT56), .ZN(n1027) );
  XNOR2_X1 U1094 ( .A(G168), .B(G1966), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1005), .B(KEYINPUT57), .ZN(n1025) );
  XNOR2_X1 U1097 ( .A(G171), .B(G1961), .ZN(n1020) );
  INV_X1 U1098 ( .A(n1006), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(G1971), .B(KEYINPUT122), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(n1009), .B(G303), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G1348), .B(n1012), .Z(n1014) );
  XNOR2_X1 U1104 ( .A(G299), .B(G1956), .ZN(n1013) );
  NOR2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(G1341), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1057) );
  INV_X1 U1113 ( .A(G16), .ZN(n1055) );
  XNOR2_X1 U1114 ( .A(G1986), .B(KEYINPUT126), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(n1028), .B(G24), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(G1976), .B(G23), .ZN(n1030) );
  XNOR2_X1 U1117 ( .A(G22), .B(G1971), .ZN(n1029) );
  NOR2_X1 U1118 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1119 ( .A(n1031), .B(KEYINPUT125), .ZN(n1032) );
  NOR2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1121 ( .A(KEYINPUT58), .B(n1034), .ZN(n1038) );
  XNOR2_X1 U1122 ( .A(G1966), .B(G21), .ZN(n1036) );
  XNOR2_X1 U1123 ( .A(G5), .B(G1961), .ZN(n1035) );
  NOR2_X1 U1124 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1125 ( .A1(n1038), .A2(n1037), .ZN(n1051) );
  XOR2_X1 U1126 ( .A(KEYINPUT124), .B(G4), .Z(n1040) );
  XNOR2_X1 U1127 ( .A(G1348), .B(KEYINPUT59), .ZN(n1039) );
  XNOR2_X1 U1128 ( .A(n1040), .B(n1039), .ZN(n1043) );
  XOR2_X1 U1129 ( .A(KEYINPUT123), .B(G1981), .Z(n1041) );
  XNOR2_X1 U1130 ( .A(G6), .B(n1041), .ZN(n1042) );
  NOR2_X1 U1131 ( .A1(n1043), .A2(n1042), .ZN(n1048) );
  XOR2_X1 U1132 ( .A(n1044), .B(G20), .Z(n1046) );
  XNOR2_X1 U1133 ( .A(G19), .B(G1341), .ZN(n1045) );
  NOR2_X1 U1134 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NAND2_X1 U1135 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  XNOR2_X1 U1136 ( .A(KEYINPUT60), .B(n1049), .ZN(n1050) );
  NOR2_X1 U1137 ( .A1(n1051), .A2(n1050), .ZN(n1052) );
  XOR2_X1 U1138 ( .A(n1052), .B(KEYINPUT127), .Z(n1053) );
  XNOR2_X1 U1139 ( .A(KEYINPUT61), .B(n1053), .ZN(n1054) );
  NAND2_X1 U1140 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  NAND2_X1 U1141 ( .A1(n1057), .A2(n1056), .ZN(n1058) );
  NOR2_X1 U1142 ( .A1(n1059), .A2(n1058), .ZN(n1060) );
  NAND2_X1 U1143 ( .A1(n1061), .A2(n1060), .ZN(n1062) );
  XOR2_X1 U1144 ( .A(KEYINPUT62), .B(n1062), .Z(G311) );
  INV_X1 U1145 ( .A(G311), .ZN(G150) );
endmodule

