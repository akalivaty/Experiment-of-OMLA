

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  INV_X1 U323 ( .A(n473), .ZN(n519) );
  XNOR2_X2 U324 ( .A(n437), .B(n436), .ZN(n576) );
  XNOR2_X1 U325 ( .A(n353), .B(n301), .ZN(n302) );
  XNOR2_X1 U326 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U327 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n359) );
  XNOR2_X1 U328 ( .A(n306), .B(n305), .ZN(n307) );
  INV_X1 U329 ( .A(n443), .ZN(n305) );
  XNOR2_X1 U330 ( .A(n295), .B(n426), .ZN(n397) );
  XOR2_X1 U331 ( .A(KEYINPUT38), .B(n452), .Z(n503) );
  XOR2_X1 U332 ( .A(n347), .B(n346), .Z(n528) );
  XNOR2_X1 U333 ( .A(n385), .B(n384), .ZN(n572) );
  XOR2_X1 U334 ( .A(KEYINPUT102), .B(n504), .Z(n291) );
  NOR2_X1 U335 ( .A1(n477), .A2(n476), .ZN(n292) );
  XOR2_X1 U336 ( .A(KEYINPUT37), .B(KEYINPUT101), .Z(n293) );
  XOR2_X1 U337 ( .A(G211GAT), .B(KEYINPUT82), .Z(n294) );
  XOR2_X1 U338 ( .A(n447), .B(n396), .Z(n295) );
  INV_X1 U339 ( .A(KEYINPUT9), .ZN(n299) );
  XNOR2_X1 U340 ( .A(n300), .B(n299), .ZN(n301) );
  INV_X1 U341 ( .A(KEYINPUT24), .ZN(n386) );
  XNOR2_X1 U342 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n457) );
  XNOR2_X1 U343 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U344 ( .A(n389), .B(n388), .ZN(n393) );
  INV_X1 U345 ( .A(KEYINPUT93), .ZN(n403) );
  XNOR2_X1 U346 ( .A(n308), .B(n307), .ZN(n310) );
  XNOR2_X1 U347 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U348 ( .A(KEYINPUT48), .B(KEYINPUT109), .ZN(n471) );
  XNOR2_X1 U349 ( .A(n367), .B(n366), .ZN(n371) );
  XNOR2_X1 U350 ( .A(n398), .B(n397), .ZN(n400) );
  XNOR2_X1 U351 ( .A(n472), .B(n471), .ZN(n527) );
  XOR2_X1 U352 ( .A(n400), .B(n399), .Z(n477) );
  XNOR2_X1 U353 ( .A(n418), .B(n293), .ZN(n517) );
  AND2_X1 U354 ( .A1(n517), .A2(n492), .ZN(n452) );
  INV_X1 U355 ( .A(G43GAT), .ZN(n486) );
  XNOR2_X1 U356 ( .A(n483), .B(G183GAT), .ZN(n484) );
  XNOR2_X1 U357 ( .A(n486), .B(KEYINPUT40), .ZN(n487) );
  XNOR2_X1 U358 ( .A(n485), .B(n484), .ZN(G1350GAT) );
  XNOR2_X1 U359 ( .A(n488), .B(n487), .ZN(G1330GAT) );
  XOR2_X1 U360 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n297) );
  XNOR2_X1 U361 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n296) );
  XOR2_X1 U362 ( .A(n297), .B(n296), .Z(n312) );
  XOR2_X1 U363 ( .A(G134GAT), .B(KEYINPUT75), .Z(n374) );
  XNOR2_X1 U364 ( .A(G36GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U365 ( .A(n298), .B(G218GAT), .ZN(n353) );
  NAND2_X1 U366 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XOR2_X1 U367 ( .A(n374), .B(n302), .Z(n308) );
  XOR2_X1 U368 ( .A(G29GAT), .B(G43GAT), .Z(n304) );
  XNOR2_X1 U369 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n303) );
  XNOR2_X1 U370 ( .A(n304), .B(n303), .ZN(n430) );
  XOR2_X1 U371 ( .A(G50GAT), .B(G162GAT), .Z(n399) );
  XNOR2_X1 U372 ( .A(n430), .B(n399), .ZN(n306) );
  XOR2_X1 U373 ( .A(G99GAT), .B(G85GAT), .Z(n443) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(G92GAT), .ZN(n309) );
  XNOR2_X1 U375 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U376 ( .A(n312), .B(n311), .ZN(n464) );
  XNOR2_X1 U377 ( .A(KEYINPUT36), .B(KEYINPUT100), .ZN(n313) );
  XNOR2_X1 U378 ( .A(n464), .B(n313), .ZN(n585) );
  XOR2_X1 U379 ( .A(G155GAT), .B(G71GAT), .Z(n315) );
  XNOR2_X1 U380 ( .A(G22GAT), .B(G127GAT), .ZN(n314) );
  XNOR2_X1 U381 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U382 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n317) );
  XNOR2_X1 U383 ( .A(G64GAT), .B(KEYINPUT76), .ZN(n316) );
  XNOR2_X1 U384 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U385 ( .A(n319), .B(n318), .ZN(n329) );
  XOR2_X1 U386 ( .A(KEYINPUT13), .B(G57GAT), .Z(n438) );
  XOR2_X1 U387 ( .A(G8GAT), .B(G183GAT), .Z(n350) );
  XOR2_X1 U388 ( .A(n438), .B(n350), .Z(n321) );
  XNOR2_X1 U389 ( .A(G78GAT), .B(G211GAT), .ZN(n320) );
  XNOR2_X1 U390 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U391 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n323) );
  NAND2_X1 U392 ( .A1(G231GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U393 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U394 ( .A(n325), .B(n324), .Z(n327) );
  XOR2_X1 U395 ( .A(G15GAT), .B(G1GAT), .Z(n425) );
  XNOR2_X1 U396 ( .A(n425), .B(KEYINPUT77), .ZN(n326) );
  XNOR2_X1 U397 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U398 ( .A(n329), .B(n328), .ZN(n583) );
  XOR2_X1 U399 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XOR2_X1 U400 ( .A(G99GAT), .B(G134GAT), .Z(n331) );
  XNOR2_X1 U401 ( .A(G43GAT), .B(G190GAT), .ZN(n330) );
  XNOR2_X1 U402 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U403 ( .A(n439), .B(n332), .Z(n334) );
  NAND2_X1 U404 ( .A1(G227GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U405 ( .A(n334), .B(n333), .ZN(n347) );
  XOR2_X1 U406 ( .A(KEYINPUT79), .B(KEYINPUT81), .Z(n336) );
  XNOR2_X1 U407 ( .A(KEYINPUT80), .B(KEYINPUT64), .ZN(n335) );
  XNOR2_X1 U408 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U409 ( .A(KEYINPUT20), .B(G176GAT), .Z(n338) );
  XNOR2_X1 U410 ( .A(G15GAT), .B(G183GAT), .ZN(n337) );
  XNOR2_X1 U411 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U412 ( .A(n340), .B(n339), .Z(n345) );
  XOR2_X1 U413 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n342) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n341) );
  XNOR2_X1 U415 ( .A(n342), .B(n341), .ZN(n356) );
  XNOR2_X1 U416 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n343) );
  XNOR2_X1 U417 ( .A(n343), .B(G127GAT), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n356), .B(n360), .ZN(n344) );
  XNOR2_X1 U419 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U420 ( .A(G64GAT), .B(G92GAT), .Z(n349) );
  XNOR2_X1 U421 ( .A(G176GAT), .B(G204GAT), .ZN(n348) );
  XNOR2_X1 U422 ( .A(n349), .B(n348), .ZN(n446) );
  XOR2_X1 U423 ( .A(n446), .B(n350), .Z(n352) );
  NAND2_X1 U424 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U425 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U426 ( .A(n354), .B(n353), .Z(n358) );
  XNOR2_X1 U427 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n355) );
  XNOR2_X1 U428 ( .A(n294), .B(n355), .ZN(n389) );
  XNOR2_X1 U429 ( .A(n356), .B(n389), .ZN(n357) );
  XNOR2_X1 U430 ( .A(n358), .B(n357), .ZN(n473) );
  XOR2_X1 U431 ( .A(n473), .B(KEYINPUT27), .Z(n409) );
  XOR2_X1 U432 ( .A(n359), .B(KEYINPUT3), .Z(n396) );
  XNOR2_X1 U433 ( .A(n360), .B(n396), .ZN(n385) );
  XOR2_X1 U434 ( .A(KEYINPUT90), .B(KEYINPUT84), .Z(n362) );
  XNOR2_X1 U435 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n361) );
  XNOR2_X1 U436 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U437 ( .A(KEYINPUT91), .B(n363), .Z(n367) );
  XNOR2_X1 U438 ( .A(KEYINPUT86), .B(KEYINPUT6), .ZN(n365) );
  NAND2_X1 U439 ( .A1(G225GAT), .A2(G233GAT), .ZN(n364) );
  XOR2_X1 U440 ( .A(KEYINPUT5), .B(KEYINPUT83), .Z(n369) );
  XNOR2_X1 U441 ( .A(G1GAT), .B(G57GAT), .ZN(n368) );
  XNOR2_X1 U442 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U443 ( .A(n371), .B(n370), .Z(n383) );
  XOR2_X1 U444 ( .A(G85GAT), .B(G148GAT), .Z(n373) );
  XNOR2_X1 U445 ( .A(G141GAT), .B(G120GAT), .ZN(n372) );
  XNOR2_X1 U446 ( .A(n373), .B(n372), .ZN(n375) );
  XOR2_X1 U447 ( .A(n375), .B(n374), .Z(n377) );
  XNOR2_X1 U448 ( .A(G29GAT), .B(G162GAT), .ZN(n376) );
  XNOR2_X1 U449 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U450 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n379) );
  XNOR2_X1 U451 ( .A(KEYINPUT85), .B(KEYINPUT89), .ZN(n378) );
  XNOR2_X1 U452 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U453 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U454 ( .A(n383), .B(n382), .ZN(n384) );
  NOR2_X1 U455 ( .A1(n409), .A2(n572), .ZN(n526) );
  NAND2_X1 U456 ( .A1(G228GAT), .A2(G233GAT), .ZN(n387) );
  XOR2_X1 U457 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n391) );
  XNOR2_X1 U458 ( .A(G218GAT), .B(G204GAT), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U460 ( .A(n393), .B(n392), .Z(n398) );
  XOR2_X1 U461 ( .A(G78GAT), .B(G148GAT), .Z(n395) );
  XNOR2_X1 U462 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n447) );
  XOR2_X1 U464 ( .A(G141GAT), .B(G22GAT), .Z(n426) );
  XOR2_X2 U465 ( .A(KEYINPUT28), .B(n477), .Z(n530) );
  NAND2_X1 U466 ( .A1(n526), .A2(n530), .ZN(n401) );
  XOR2_X1 U467 ( .A(KEYINPUT92), .B(n401), .Z(n402) );
  NAND2_X1 U468 ( .A1(n528), .A2(n402), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n404), .B(n403), .ZN(n415) );
  NOR2_X1 U470 ( .A1(n528), .A2(n519), .ZN(n405) );
  NOR2_X1 U471 ( .A1(n477), .A2(n405), .ZN(n406) );
  XOR2_X1 U472 ( .A(n406), .B(KEYINPUT25), .Z(n407) );
  XNOR2_X1 U473 ( .A(KEYINPUT94), .B(n407), .ZN(n411) );
  NAND2_X1 U474 ( .A1(n477), .A2(n528), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n408), .B(KEYINPUT26), .ZN(n575) );
  NOR2_X1 U476 ( .A1(n575), .A2(n409), .ZN(n410) );
  NOR2_X1 U477 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U478 ( .A(KEYINPUT95), .B(n412), .ZN(n413) );
  NAND2_X1 U479 ( .A1(n413), .A2(n572), .ZN(n414) );
  NAND2_X1 U480 ( .A1(n415), .A2(n414), .ZN(n416) );
  XOR2_X1 U481 ( .A(KEYINPUT96), .B(n416), .Z(n491) );
  NOR2_X1 U482 ( .A1(n583), .A2(n491), .ZN(n417) );
  NAND2_X1 U483 ( .A1(n585), .A2(n417), .ZN(n418) );
  XOR2_X1 U484 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n420) );
  XNOR2_X1 U485 ( .A(G113GAT), .B(G8GAT), .ZN(n419) );
  XNOR2_X1 U486 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U487 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n422) );
  XNOR2_X1 U488 ( .A(KEYINPUT70), .B(KEYINPUT67), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U490 ( .A(n424), .B(n423), .ZN(n437) );
  XOR2_X1 U491 ( .A(G50GAT), .B(G36GAT), .Z(n428) );
  XNOR2_X1 U492 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U494 ( .A(n429), .B(G197GAT), .Z(n435) );
  XOR2_X1 U495 ( .A(n430), .B(KEYINPUT69), .Z(n432) );
  NAND2_X1 U496 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U497 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n436) );
  INV_X1 U500 ( .A(n576), .ZN(n532) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n451) );
  XOR2_X1 U502 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n441) );
  XNOR2_X1 U503 ( .A(KEYINPUT32), .B(KEYINPUT73), .ZN(n440) );
  XNOR2_X1 U504 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U505 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U506 ( .A1(G230GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U508 ( .A(n447), .B(n446), .Z(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(n461) );
  INV_X1 U511 ( .A(n461), .ZN(n579) );
  NOR2_X1 U512 ( .A1(n532), .A2(n579), .ZN(n492) );
  NOR2_X1 U513 ( .A1(n503), .A2(n572), .ZN(n456) );
  XNOR2_X1 U514 ( .A(KEYINPUT99), .B(KEYINPUT39), .ZN(n454) );
  INV_X1 U515 ( .A(G29GAT), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n456), .B(n455), .ZN(G1328GAT) );
  INV_X1 U518 ( .A(KEYINPUT123), .ZN(n482) );
  NAND2_X1 U519 ( .A1(n583), .A2(n585), .ZN(n458) );
  NOR2_X1 U520 ( .A1(n579), .A2(n576), .ZN(n459) );
  AND2_X1 U521 ( .A1(n460), .A2(n459), .ZN(n470) );
  XOR2_X1 U522 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n463) );
  XOR2_X1 U523 ( .A(KEYINPUT41), .B(n461), .Z(n534) );
  INV_X1 U524 ( .A(n534), .ZN(n563) );
  NAND2_X1 U525 ( .A1(n563), .A2(n576), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n463), .B(n462), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n464), .A2(n583), .ZN(n465) );
  NAND2_X1 U528 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U529 ( .A(KEYINPUT108), .B(n467), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n468), .B(KEYINPUT47), .ZN(n469) );
  NOR2_X1 U531 ( .A1(n470), .A2(n469), .ZN(n472) );
  NAND2_X1 U532 ( .A1(n473), .A2(n527), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n474), .B(KEYINPUT121), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT54), .ZN(n573) );
  INV_X1 U535 ( .A(n572), .ZN(n476) );
  AND2_X1 U536 ( .A1(n573), .A2(n292), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U539 ( .A1(n528), .A2(n480), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(n567) );
  NAND2_X1 U541 ( .A1(n567), .A2(n583), .ZN(n485) );
  XOR2_X1 U542 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n483) );
  NOR2_X1 U543 ( .A1(n528), .A2(n503), .ZN(n488) );
  INV_X1 U544 ( .A(n583), .ZN(n538) );
  NOR2_X1 U545 ( .A1(n464), .A2(n538), .ZN(n489) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n489), .Z(n490) );
  NOR2_X1 U547 ( .A1(n491), .A2(n490), .ZN(n505) );
  NAND2_X1 U548 ( .A1(n492), .A2(n505), .ZN(n499) );
  NOR2_X1 U549 ( .A1(n572), .A2(n499), .ZN(n494) );
  XNOR2_X1 U550 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(n495), .ZN(G1324GAT) );
  NOR2_X1 U553 ( .A1(n519), .A2(n499), .ZN(n496) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  NOR2_X1 U555 ( .A1(n528), .A2(n499), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n530), .A2(n499), .ZN(n500) );
  XOR2_X1 U559 ( .A(KEYINPUT98), .B(n500), .Z(n501) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n501), .ZN(G1327GAT) );
  NOR2_X1 U561 ( .A1(n503), .A2(n519), .ZN(n502) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U563 ( .A1(n503), .A2(n530), .ZN(n504) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n291), .ZN(G1331GAT) );
  NOR2_X1 U565 ( .A1(n534), .A2(n576), .ZN(n516) );
  NAND2_X1 U566 ( .A1(n516), .A2(n505), .ZN(n512) );
  NOR2_X1 U567 ( .A1(n572), .A2(n512), .ZN(n507) );
  XNOR2_X1 U568 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n519), .A2(n512), .ZN(n509) );
  XOR2_X1 U572 ( .A(KEYINPUT104), .B(n509), .Z(n510) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n510), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n528), .A2(n512), .ZN(n511) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n511), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n530), .A2(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n515), .Z(G1335GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n516), .ZN(n522) );
  NOR2_X1 U581 ( .A1(n572), .A2(n522), .ZN(n518) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n522), .ZN(n520) );
  XOR2_X1 U584 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U585 ( .A1(n528), .A2(n522), .ZN(n521) );
  XOR2_X1 U586 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U587 ( .A1(n530), .A2(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT106), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U590 ( .A(G106GAT), .B(n525), .Z(G1339GAT) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n548) );
  NOR2_X1 U592 ( .A1(n528), .A2(n548), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(KEYINPUT110), .ZN(n531) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n543) );
  NOR2_X1 U595 ( .A1(n532), .A2(n543), .ZN(n533) );
  XOR2_X1 U596 ( .A(G113GAT), .B(n533), .Z(G1340GAT) );
  NOR2_X1 U597 ( .A1(n534), .A2(n543), .ZN(n536) );
  XNOR2_X1 U598 ( .A(KEYINPUT111), .B(KEYINPUT49), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  NOR2_X1 U601 ( .A1(n538), .A2(n543), .ZN(n540) );
  XNOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT112), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U604 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  INV_X1 U605 ( .A(n464), .ZN(n542) );
  NOR2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n547) );
  XOR2_X1 U607 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n545) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT113), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n550) );
  NOR2_X1 U612 ( .A1(n575), .A2(n548), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n559), .A2(n576), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n553) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(n554), .Z(n556) );
  NAND2_X1 U620 ( .A1(n559), .A2(n563), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT119), .Z(n558) );
  NAND2_X1 U623 ( .A1(n559), .A2(n583), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n464), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT120), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n567), .A2(n576), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n565) );
  NAND2_X1 U631 ( .A1(n567), .A2(n563), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n464), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT58), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(n569), .ZN(G1351GAT) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n570), .B(KEYINPUT126), .ZN(n571) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(n571), .Z(n578) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n586) );
  NAND2_X1 U642 ( .A1(n586), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n586), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  NAND2_X1 U648 ( .A1(n586), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(KEYINPUT62), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

