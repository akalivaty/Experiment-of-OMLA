//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n562, new_n563, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G238), .A3(G237), .A4(G235), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(G137), .A3(new_n464), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n472), .A2(new_n464), .A3(G101), .A4(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n475), .ZN(G160));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(KEYINPUT69), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n464), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n492), .B2(G114), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(KEYINPUT70), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n477), .B2(new_n478), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n477), .B2(new_n478), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n501), .B(new_n504), .C1(new_n478), .C2(new_n477), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT71), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT5), .B1(new_n508), .B2(KEYINPUT71), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g086(.A(KEYINPUT71), .B(KEYINPUT5), .C1(new_n507), .C2(new_n508), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(G88), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n508), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n511), .A2(new_n512), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n521), .B1(new_n520), .B2(new_n526), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  AOI21_X1  g106(.A(new_n523), .B1(new_n514), .B2(new_n515), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n518), .A2(G51), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n533), .A2(new_n534), .A3(new_n537), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n518), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n513), .A2(new_n516), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n513), .A2(G64), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n544), .A2(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n523), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n511), .A2(G81), .A3(new_n512), .A4(new_n516), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n518), .A2(G43), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G860), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT76), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT77), .ZN(G188));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n523), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n511), .A2(G91), .A3(new_n512), .A4(new_n516), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT78), .B(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n518), .A2(new_n572), .A3(G53), .A4(new_n573), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n518), .A2(G53), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n518), .A2(G53), .A3(new_n573), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(KEYINPUT79), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n570), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  NAND2_X1  g159(.A1(new_n532), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n518), .A2(G49), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  NAND3_X1  g163(.A1(new_n513), .A2(G86), .A3(new_n516), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n518), .A2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n523), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n518), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n542), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n513), .A2(G60), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n545), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT81), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n511), .A2(G92), .A3(new_n512), .A4(new_n516), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n608), .A2(KEYINPUT82), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n608), .A2(KEYINPUT82), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  OR3_X1    g186(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n609), .B2(new_n610), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n523), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n612), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n607), .B1(G868), .B2(new_n619), .ZN(G284));
  XOR2_X1   g195(.A(G284), .B(KEYINPUT83), .Z(G321));
  MUX2_X1   g196(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g197(.A(G280), .B(KEYINPUT84), .Z(G297));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n619), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n619), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(new_n557), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(G868), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n488), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n483), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n464), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  XOR2_X1   g211(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n636), .A2(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT14), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n663), .B2(new_n659), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(new_n684), .B(new_n683), .S(new_n676), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT89), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n688), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n690), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n691), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n691), .B2(new_n695), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n673), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n691), .A2(new_n695), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(new_n696), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n691), .A2(new_n695), .A3(new_n697), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n702), .A2(new_n672), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(new_n704), .ZN(G229));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G21), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G168), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G1966), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT97), .ZN(new_n710));
  NOR2_X1   g285(.A1(G29), .A2(G35), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G162), .B2(G29), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G2090), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n619), .A2(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G4), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G1348), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G27), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G164), .B2(new_n721), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT98), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(G33), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n728));
  NAND3_X1  g303(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n464), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G139), .B2(new_n488), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n733), .B2(new_n721), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2072), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G1966), .B2(new_n708), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n716), .A2(new_n720), .A3(new_n726), .A4(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n718), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(G1348), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G299), .A2(G16), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n706), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT23), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G1956), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n706), .A2(G19), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT91), .Z(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n628), .B2(new_n706), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT92), .Z(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n721), .A2(G26), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT28), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n483), .A2(G128), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n756));
  INV_X1    g331(.A(G116), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G2105), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n488), .B2(G140), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n752), .B1(new_n760), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  AND2_X1   g337(.A1(KEYINPUT24), .A2(G34), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n721), .B1(KEYINPUT24), .B2(G34), .ZN(new_n764));
  OAI22_X1  g339(.A1(G160), .A2(new_n721), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G28), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT30), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n768), .B2(KEYINPUT30), .ZN(new_n770));
  OR2_X1    g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  NAND2_X1  g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n767), .B(new_n773), .C1(new_n721), .C2(new_n635), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n706), .A2(G5), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G171), .B2(new_n706), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n776), .A2(G1961), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(G1961), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n774), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AND3_X1   g354(.A1(new_n750), .A2(new_n762), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n721), .A2(G32), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n488), .A2(G141), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n488), .A2(KEYINPUT95), .A3(G141), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT26), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n788), .B(new_n789), .C1(new_n483), .C2(G129), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n786), .A2(KEYINPUT96), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n781), .B1(new_n796), .B2(new_n721), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT27), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1996), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n739), .A2(new_n745), .A3(new_n780), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G6), .A2(G16), .ZN(new_n801));
  INV_X1    g376(.A(new_n596), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(new_n591), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n801), .B1(new_n803), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT32), .ZN(new_n805));
  INV_X1    g380(.A(G1981), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n706), .A2(G22), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G166), .B2(new_n706), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(G1971), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n706), .A2(G23), .ZN(new_n811));
  INV_X1    g386(.A(G288), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n706), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT33), .B(G1976), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n809), .B2(G1971), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n807), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G24), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n604), .B(KEYINPUT90), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(G16), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1986), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n488), .A2(G131), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n483), .A2(G119), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n464), .A2(G107), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  MUX2_X1   g403(.A(G25), .B(new_n828), .S(G29), .Z(new_n829));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G1991), .Z(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n829), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n818), .A2(new_n819), .A3(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n800), .B1(new_n835), .B2(new_n836), .ZN(G311));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  INV_X1    g413(.A(new_n800), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(G150));
  NOR2_X1   g415(.A1(new_n618), .A2(new_n624), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n511), .A2(G67), .A3(new_n512), .ZN(new_n844));
  NAND2_X1  g419(.A1(G80), .A2(G543), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n545), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n511), .A2(G93), .A3(new_n512), .A4(new_n516), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n518), .A2(G55), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n557), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n846), .A2(new_n849), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n851), .A2(new_n553), .A3(new_n556), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n843), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n856), .B2(new_n855), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n851), .A2(new_n558), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n828), .B(new_n639), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n483), .A2(G130), .ZN(new_n863));
  OR2_X1    g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(G142), .B2(new_n488), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n862), .B(new_n867), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT102), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n492), .A2(G114), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n494), .A2(KEYINPUT70), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(G2105), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n872), .A2(new_n491), .B1(new_n465), .B2(new_n497), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n504), .B1(new_n465), .B2(new_n501), .ZN(new_n874));
  INV_X1    g449(.A(new_n505), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n794), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT96), .B1(new_n786), .B2(new_n790), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n793), .A2(G164), .A3(new_n794), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n879), .A2(new_n760), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n760), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n733), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n760), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n877), .A2(new_n876), .A3(new_n878), .ZN(new_n886));
  AOI21_X1  g461(.A(G164), .B1(new_n793), .B2(new_n794), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n879), .A2(new_n760), .A3(new_n880), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n733), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n869), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n635), .B(G160), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G162), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n883), .B1(new_n881), .B2(new_n882), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n888), .A2(new_n733), .A3(new_n889), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n895), .A2(KEYINPUT102), .A3(new_n896), .A4(new_n868), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n868), .B1(new_n884), .B2(new_n890), .ZN(new_n899));
  INV_X1    g474(.A(new_n868), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n893), .A3(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(KEYINPUT101), .B(G37), .Z(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n898), .A2(new_n902), .A3(KEYINPUT103), .A4(new_n903), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n906), .A2(KEYINPUT40), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT40), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(G395));
  XNOR2_X1  g485(.A(new_n626), .B(new_n854), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n613), .A2(new_n617), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n612), .A4(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n618), .B1(new_n581), .B2(new_n582), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n911), .A2(KEYINPUT104), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT104), .B1(new_n911), .B2(new_n918), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT41), .B1(new_n915), .B2(new_n916), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT41), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n911), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n925));
  XNOR2_X1  g500(.A(G305), .B(new_n604), .ZN(new_n926));
  INV_X1    g501(.A(new_n526), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n517), .A2(new_n519), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT73), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n527), .A3(G288), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G288), .B1(new_n929), .B2(new_n527), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n604), .B(new_n803), .ZN(new_n934));
  INV_X1    g509(.A(new_n932), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n919), .A2(new_n939), .A3(new_n920), .A4(new_n923), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n925), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n938), .B1(new_n925), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(G868), .B2(new_n851), .ZN(G295));
  OAI21_X1  g519(.A(new_n943), .B1(G868), .B2(new_n851), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n946));
  AOI21_X1  g521(.A(G286), .B1(G171), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT106), .B1(new_n544), .B2(new_n548), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n850), .A2(new_n949), .A3(new_n852), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n850), .B2(new_n852), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n949), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n853), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n850), .A2(new_n949), .A3(new_n852), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n947), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n952), .A2(new_n956), .A3(new_n917), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n922), .A2(new_n959), .B1(new_n952), .B2(new_n956), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n917), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT41), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(KEYINPUT108), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n958), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n965), .A2(new_n938), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n952), .A2(new_n956), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n922), .B2(new_n921), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n938), .A3(new_n957), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n969), .A2(new_n903), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n966), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n903), .B(new_n969), .C1(new_n965), .C2(new_n938), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT109), .B1(new_n974), .B2(KEYINPUT43), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n962), .A2(new_n963), .B1(new_n956), .B2(new_n952), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n937), .B1(new_n976), .B2(new_n958), .ZN(new_n977));
  INV_X1    g552(.A(G37), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n969), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT43), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n979), .B2(KEYINPUT43), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n973), .B(new_n975), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n977), .A2(new_n969), .A3(new_n972), .A4(new_n978), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(KEYINPUT44), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n987), .A2(new_n991), .A3(KEYINPUT44), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n986), .A2(new_n993), .ZN(G397));
  INV_X1    g569(.A(G2067), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n885), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n760), .A2(G2067), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n996), .A2(KEYINPUT114), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT114), .B1(new_n996), .B2(new_n997), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n796), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1996), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n998), .B2(new_n999), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT111), .B(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n876), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1005), .A2(KEYINPUT112), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G40), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n468), .A2(new_n475), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1000), .A2(new_n1002), .A3(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n828), .A2(new_n831), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n828), .A2(new_n831), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1013), .A2(new_n795), .A3(G1996), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT113), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n604), .B(G1986), .Z(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n503), .A2(new_n505), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1384), .B1(new_n1024), .B2(new_n873), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1012), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT115), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(KEYINPUT115), .A3(new_n1026), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1384), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1025), .A2(KEYINPUT117), .A3(KEYINPUT45), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1003), .B1(G164), .B2(G1384), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1012), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1031), .A2(new_n766), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G8), .ZN(new_n1041));
  OR3_X1    g616(.A1(new_n1040), .A2(new_n1041), .A3(G168), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1043));
  INV_X1    g618(.A(G125), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n467), .B1(new_n479), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(G2105), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(G40), .A3(new_n469), .A4(new_n474), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n876), .A2(new_n1032), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(KEYINPUT50), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1030), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n766), .B(new_n1049), .C1(new_n1050), .C2(new_n1028), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1041), .B1(new_n1043), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G168), .A2(new_n1041), .ZN(new_n1053));
  OR3_X1    g628(.A1(new_n1052), .A2(KEYINPUT51), .A3(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1053), .B1(new_n1052), .B2(KEYINPUT123), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1055), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1054), .B1(new_n1059), .B2(KEYINPUT124), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT124), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1061), .B(new_n1055), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1042), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT62), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1065), .B(new_n1042), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1012), .B1(new_n1025), .B2(KEYINPUT45), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1005), .A2(new_n1003), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G1971), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G2090), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1031), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1041), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n929), .A2(new_n527), .A3(G8), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n592), .A2(new_n806), .A3(new_n596), .ZN(new_n1079));
  OAI21_X1  g654(.A(G1981), .B1(new_n802), .B2(new_n591), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT49), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT49), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1012), .A2(new_n1025), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G8), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n812), .A2(G1976), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n1088), .A3(G8), .A4(new_n1083), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G288), .A2(new_n1087), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT52), .B1(new_n1090), .B2(new_n1084), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1085), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1075), .B(KEYINPUT55), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1049), .B1(KEYINPUT50), .B2(new_n1048), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(G2090), .ZN(new_n1096));
  OAI21_X1  g671(.A(G8), .B1(new_n1096), .B2(new_n1070), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1078), .A2(new_n1093), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1069), .A2(new_n724), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1049), .B1(new_n1050), .B2(new_n1028), .ZN(new_n1102));
  INV_X1    g677(.A(G1961), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1100), .A2(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n1038), .A2(new_n1101), .A3(G2078), .ZN(new_n1105));
  AOI21_X1  g680(.A(G301), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1099), .A2(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1064), .A2(new_n1066), .A3(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n580), .B(KEYINPUT57), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1047), .B1(new_n1048), .B2(new_n1003), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1095), .A2(new_n744), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1110), .A2(new_n1111), .A3(KEYINPUT118), .A4(new_n1112), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1109), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(KEYINPUT120), .A3(new_n1115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  AND4_X1   g698(.A1(new_n1109), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1083), .B(KEYINPUT119), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1128), .A2(new_n995), .B1(new_n1102), .B2(new_n719), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n618), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(new_n618), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT60), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1109), .B1(new_n1121), .B2(new_n1115), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1125), .B1(new_n1134), .B2(new_n1124), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1083), .A2(KEYINPUT119), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1012), .B2(new_n1025), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT58), .B(G1341), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1067), .A2(new_n1068), .A3(G1996), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n628), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1144), .B(new_n628), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n618), .A2(KEYINPUT60), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1143), .A2(new_n1145), .B1(new_n1129), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1127), .A2(new_n1133), .A3(new_n1135), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1124), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1149), .B(new_n1150), .C1(new_n1151), .C2(new_n1132), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1132), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT121), .B1(new_n1153), .B2(new_n1124), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1148), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n469), .A2(new_n474), .A3(KEYINPUT125), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT125), .B1(new_n469), .B2(new_n474), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n724), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1159));
  NOR4_X1   g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n468), .A4(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1110), .B(new_n1160), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1104), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(G171), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1156), .B1(new_n1163), .B2(new_n1106), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1099), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1104), .A2(G301), .A3(new_n1105), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT54), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1162), .A2(G171), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT126), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1162), .A2(new_n1170), .A3(G171), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1167), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1165), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1155), .A2(new_n1173), .A3(new_n1063), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1093), .A2(new_n1077), .A3(new_n1074), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1085), .A2(G1976), .A3(G288), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1079), .B(KEYINPUT116), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1175), .B1(new_n1178), .B2(new_n1084), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1040), .A2(new_n1041), .A3(G286), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1099), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT63), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1180), .A2(KEYINPUT63), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1184), .A2(new_n1185), .A3(new_n1078), .A4(new_n1093), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1179), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1174), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1023), .B1(new_n1108), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1015), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n996), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1190), .B1(new_n1192), .B2(new_n1014), .ZN(new_n1193));
  AOI211_X1 g768(.A(KEYINPUT127), .B(new_n1013), .C1(new_n1191), .C2(new_n996), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1000), .A2(new_n1014), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1014), .A2(new_n1001), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT46), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT47), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1198), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1013), .A2(G1986), .A3(G290), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT48), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1200), .A2(new_n1201), .B1(new_n1021), .B2(new_n1203), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1193), .A2(new_n1194), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1189), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g781(.A1(new_n906), .A2(new_n907), .ZN(new_n1208));
  NOR3_X1   g782(.A1(new_n462), .A2(G401), .A3(G227), .ZN(new_n1209));
  AND3_X1   g783(.A1(new_n700), .A2(new_n704), .A3(new_n1209), .ZN(new_n1210));
  AND3_X1   g784(.A1(new_n1208), .A2(new_n1210), .A3(new_n984), .ZN(G308));
  NAND3_X1  g785(.A1(new_n1208), .A2(new_n1210), .A3(new_n984), .ZN(G225));
endmodule


