//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT79), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G104), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT79), .A3(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(KEYINPUT78), .A3(G104), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(KEYINPUT78), .A3(KEYINPUT3), .A4(G104), .ZN(new_n197));
  AOI221_X4 g011(.A(G101), .B1(new_n191), .B2(new_n193), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n192), .A2(G107), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n192), .A2(G107), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT80), .B1(new_n198), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G116), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(KEYINPUT66), .A3(G119), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT5), .ZN(new_n212));
  INV_X1    g026(.A(G113), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT5), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(new_n206), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT2), .B(G113), .Z(new_n216));
  AOI22_X1  g030(.A1(new_n212), .A2(new_n215), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n191), .A2(new_n193), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT3), .B1(new_n200), .B2(KEYINPUT78), .ZN(new_n219));
  INV_X1    g033(.A(new_n197), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n199), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT80), .ZN(new_n222));
  INV_X1    g036(.A(new_n203), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n204), .A2(new_n217), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n211), .B(new_n216), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G101), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n221), .A2(KEYINPUT4), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n196), .A2(new_n197), .B1(new_n191), .B2(new_n193), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(new_n199), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n226), .B(new_n229), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n225), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n225), .A2(new_n233), .A3(new_n235), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(KEYINPUT6), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT0), .A4(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n242), .A2(G146), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n240), .B2(G143), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(KEYINPUT64), .A3(G146), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT0), .B(G128), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G125), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n241), .A2(new_n243), .A3(new_n253), .A4(G128), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n241), .B2(KEYINPUT1), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n249), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n252), .B1(G125), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G224), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G953), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n234), .A2(new_n262), .A3(new_n236), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n239), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n239), .A2(KEYINPUT83), .A3(new_n261), .A4(new_n263), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G902), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n235), .B(KEYINPUT8), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n203), .B1(new_n231), .B2(new_n199), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n217), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n217), .A2(new_n271), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT84), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT7), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI22_X1  g091(.A1(new_n258), .A2(new_n277), .B1(new_n276), .B2(new_n260), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n258), .A2(new_n260), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(KEYINPUT7), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n274), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n238), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n269), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n188), .B1(new_n268), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n188), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n286), .B(new_n283), .C1(new_n266), .C2(new_n267), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n187), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G469), .ZN(new_n289));
  INV_X1    g103(.A(new_n257), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT81), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n290), .B(new_n291), .C1(new_n198), .C2(new_n203), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT81), .B1(new_n271), .B2(new_n257), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n241), .A2(new_n243), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n254), .B1(new_n294), .B2(new_n256), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n271), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G137), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G134), .ZN(new_n299));
  NOR2_X1   g113(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G134), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G137), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(G137), .ZN(new_n306));
  AND2_X1   g120(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G131), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n298), .A2(G134), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(new_n299), .B2(new_n302), .ZN(new_n311));
  INV_X1    g125(.A(G131), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n306), .B1(new_n307), .B2(new_n300), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n297), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT12), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n297), .A2(KEYINPUT12), .A3(new_n315), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n227), .A2(G101), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n324), .B(new_n244), .C1(new_n249), .C2(new_n250), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n322), .A2(new_n323), .A3(new_n325), .A4(new_n229), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n204), .A2(KEYINPUT10), .A3(new_n257), .A4(new_n224), .ZN(new_n327));
  INV_X1    g141(.A(new_n315), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT10), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n296), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G110), .B(G140), .ZN(new_n332));
  INV_X1    g146(.A(G953), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n333), .A2(G227), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n332), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n320), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n326), .A2(new_n327), .A3(new_n330), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n315), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n336), .B1(new_n341), .B2(new_n331), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n289), .B(new_n269), .C1(new_n339), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n337), .A2(KEYINPUT82), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n331), .A2(new_n336), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT82), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n347), .A3(new_n341), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n320), .A2(new_n331), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n335), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n350), .A3(G469), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n289), .A2(new_n269), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n343), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT9), .B(G234), .ZN(new_n355));
  OAI21_X1  g169(.A(G221), .B1(new_n355), .B2(G902), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n288), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G217), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(G234), .B2(new_n269), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT75), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G137), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G140), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G125), .ZN(new_n367));
  INV_X1    g181(.A(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G140), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT16), .ZN(new_n370));
  OR3_X1    g184(.A1(new_n368), .A2(KEYINPUT16), .A3(G140), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G146), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(G146), .B1(new_n370), .B2(new_n371), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n255), .A2(G119), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n208), .A2(G128), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT24), .B(G110), .ZN(new_n378));
  OAI22_X1  g192(.A1(new_n373), .A2(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT73), .B1(new_n208), .B2(G128), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT23), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT23), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(KEYINPUT73), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n383), .A3(new_n376), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G110), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT74), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(KEYINPUT74), .A3(G110), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n379), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n377), .A2(new_n378), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n384), .B2(G110), .ZN(new_n391));
  XNOR2_X1  g205(.A(G125), .B(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n240), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n372), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n365), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n379), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n387), .A2(new_n388), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n394), .A3(new_n364), .ZN(new_n400));
  AOI21_X1  g214(.A(G902), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT25), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  AOI211_X1 g219(.A(G902), .B(new_n403), .C1(new_n396), .C2(new_n400), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n360), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n360), .A2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n396), .A2(new_n400), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT77), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n407), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(G472), .A2(G902), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n323), .A2(new_n315), .A3(new_n325), .ZN(new_n415));
  OAI21_X1  g229(.A(G131), .B1(new_n306), .B2(new_n310), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n257), .A2(new_n314), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(KEYINPUT30), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n257), .A2(new_n314), .A3(new_n416), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n251), .B1(new_n314), .B2(new_n309), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n422), .A3(new_n226), .ZN(new_n423));
  INV_X1    g237(.A(new_n226), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n415), .A2(new_n424), .A3(new_n417), .ZN(new_n425));
  NOR2_X1   g239(.A1(G237), .A2(G953), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G210), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT27), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT26), .B(G101), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n423), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT31), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT68), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT68), .B(KEYINPUT31), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n423), .A2(new_n425), .A3(new_n430), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n421), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n424), .B1(new_n439), .B2(new_n417), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n425), .A2(KEYINPUT28), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT28), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n415), .A2(new_n442), .A3(new_n424), .A4(new_n417), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n440), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(new_n430), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n414), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT69), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n434), .B(new_n437), .C1(new_n444), .C2(new_n430), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT69), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n414), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n424), .B1(new_n415), .B2(new_n417), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n441), .B2(new_n443), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n430), .A2(KEYINPUT29), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT71), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n423), .A2(new_n425), .ZN(new_n460));
  INV_X1    g274(.A(new_n430), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI211_X1 g276(.A(KEYINPUT71), .B(new_n430), .C1(new_n423), .C2(new_n425), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT29), .B1(new_n444), .B2(new_n430), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n458), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G472), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT72), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n460), .A2(new_n461), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT71), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n460), .A2(new_n459), .A3(new_n461), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n465), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n457), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(G472), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n448), .A2(KEYINPUT32), .A3(new_n414), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n452), .A2(new_n468), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n355), .A2(new_n359), .A3(G953), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n480));
  OR2_X1    g294(.A1(KEYINPUT88), .A2(G122), .ZN(new_n481));
  NAND2_X1  g295(.A1(KEYINPUT88), .A2(G122), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n205), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n205), .A2(G122), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n483), .A2(KEYINPUT89), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n487));
  AND2_X1   g301(.A1(KEYINPUT88), .A2(G122), .ZN(new_n488));
  NOR2_X1   g302(.A1(KEYINPUT88), .A2(G122), .ZN(new_n489));
  OAI21_X1  g303(.A(G116), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n490), .B2(new_n484), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n480), .B(new_n190), .C1(new_n486), .C2(new_n491), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n484), .A2(KEYINPUT14), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n484), .A2(KEYINPUT14), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n242), .A2(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n255), .A2(G143), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n304), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G134), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n495), .A2(G107), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT89), .B1(new_n483), .B2(new_n485), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n490), .A2(new_n487), .A3(new_n484), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n480), .B1(new_n505), .B2(new_n190), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n496), .A2(KEYINPUT13), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT13), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n508), .B(G134), .C1(new_n509), .C2(new_n499), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n498), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n190), .B1(new_n486), .B2(new_n491), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n503), .A2(G107), .A3(new_n504), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n479), .B1(new_n507), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(KEYINPUT90), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n492), .A3(new_n501), .ZN(new_n517));
  INV_X1    g331(.A(new_n514), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n518), .A3(new_n478), .ZN(new_n519));
  AOI211_X1 g333(.A(KEYINPUT91), .B(G902), .C1(new_n515), .C2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G478), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(G902), .B1(new_n515), .B2(new_n519), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n523), .B1(new_n526), .B2(new_n522), .ZN(new_n527));
  INV_X1    g341(.A(G475), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n392), .B(new_n240), .ZN(new_n529));
  OR2_X1    g343(.A1(KEYINPUT85), .A2(G143), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(G214), .A3(new_n426), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT85), .B(G143), .Z(new_n532));
  AND2_X1   g346(.A1(new_n426), .A2(G214), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(new_n312), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n530), .A2(G214), .A3(new_n426), .ZN(new_n537));
  NAND2_X1  g351(.A1(KEYINPUT85), .A2(G143), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n530), .A2(new_n538), .B1(new_n426), .B2(G214), .ZN(new_n539));
  OAI21_X1  g353(.A(G131), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI221_X1 g354(.A(new_n529), .B1(new_n534), .B2(new_n536), .C1(new_n540), .C2(new_n535), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n312), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT86), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n540), .A2(new_n542), .A3(KEYINPUT86), .A4(new_n544), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n373), .A2(new_n374), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n534), .A2(KEYINPUT17), .A3(G131), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n541), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G113), .B(G122), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(new_n192), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n552), .B(new_n541), .C1(new_n545), .C2(new_n549), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n528), .B1(new_n556), .B2(new_n269), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT19), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n392), .B(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n372), .B1(new_n559), .B2(G146), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n541), .B1(new_n543), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n553), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT87), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(G475), .A2(G902), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n555), .A2(new_n562), .A3(KEYINPUT87), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT20), .ZN(new_n569));
  NOR3_X1   g383(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n557), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G952), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(G953), .ZN(new_n574));
  NAND2_X1  g388(.A1(G234), .A2(G237), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT21), .B(G898), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(G902), .A3(G953), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n527), .A2(new_n572), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n358), .A2(new_n413), .A3(new_n477), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  OAI211_X1 g397(.A(new_n580), .B(new_n187), .C1(new_n285), .C2(new_n287), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n515), .A2(new_n519), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT33), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n515), .A2(new_n519), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(G478), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n269), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n524), .B2(new_n590), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n572), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n584), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n356), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n341), .A2(new_n331), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n335), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n599), .B2(new_n338), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n352), .B1(new_n600), .B2(new_n289), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n601), .B2(new_n351), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n447), .A2(new_n450), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n448), .A2(new_n269), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G472), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT92), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n467), .B1(new_n448), .B2(new_n269), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n603), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n596), .A2(new_n413), .A3(new_n602), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G104), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  INV_X1    g428(.A(new_n584), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT20), .ZN(new_n616));
  AND4_X1   g430(.A1(new_n616), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n569), .A3(KEYINPUT94), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n555), .A2(new_n562), .A3(KEYINPUT87), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT87), .B1(new_n555), .B2(new_n562), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n616), .B1(new_n623), .B2(new_n566), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n620), .B1(new_n624), .B2(new_n617), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n626), .A2(new_n557), .A3(new_n527), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n615), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n606), .A2(new_n609), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n354), .A2(new_n413), .A3(new_n356), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n630), .A2(new_n631), .A3(new_n603), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NAND2_X1  g449(.A1(new_n399), .A2(new_n394), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n408), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n407), .A2(KEYINPUT95), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT95), .B1(new_n407), .B2(new_n639), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n358), .A2(new_n581), .A3(new_n610), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  NOR2_X1   g459(.A1(new_n524), .A2(new_n525), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n522), .B1(new_n646), .B2(new_n520), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n524), .A2(new_n525), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n521), .A3(G478), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n557), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n579), .A2(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n576), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n619), .A2(new_n650), .A3(new_n625), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n477), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n268), .A2(new_n284), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n286), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n268), .A2(new_n188), .A3(new_n284), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n658), .A2(new_n602), .A3(new_n187), .A4(new_n642), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n255), .ZN(G30));
  XOR2_X1   g475(.A(new_n658), .B(KEYINPUT38), .Z(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n652), .B(KEYINPUT39), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n602), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(KEYINPUT40), .Z(new_n666));
  AOI21_X1  g480(.A(new_n461), .B1(new_n423), .B2(new_n425), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n425), .A2(new_n461), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n269), .B1(new_n668), .B2(new_n453), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n476), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n452), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n187), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n407), .A2(new_n639), .ZN(new_n675));
  INV_X1    g489(.A(new_n572), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n647), .A2(new_n649), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR4_X1   g492(.A1(new_n673), .A2(new_n674), .A3(new_n675), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n663), .A2(new_n666), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  INV_X1    g495(.A(new_n593), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n568), .A2(KEYINPUT20), .B1(new_n563), .B2(new_n570), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n682), .B(new_n652), .C1(new_n557), .C2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT96), .B1(new_n288), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT96), .ZN(new_n686));
  INV_X1    g500(.A(new_n652), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n572), .A2(new_n593), .A3(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n658), .A2(new_n686), .A3(new_n187), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n642), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n467), .B1(new_n472), .B2(new_n457), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n476), .B1(new_n692), .B2(new_n474), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n466), .A2(KEYINPUT72), .A3(new_n467), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n691), .B1(new_n695), .B2(new_n452), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n690), .A2(new_n602), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  INV_X1    g512(.A(new_n596), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n342), .B1(new_n320), .B2(new_n337), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n701), .A2(new_n356), .A3(new_n343), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n477), .A2(new_n413), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT41), .B(G113), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NOR2_X1   g520(.A1(new_n628), .A2(new_n703), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n205), .ZN(G18));
  NAND3_X1  g522(.A1(new_n477), .A2(new_n581), .A3(new_n642), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT97), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n701), .A2(new_n356), .A3(new_n343), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n710), .B1(new_n288), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n674), .B1(new_n656), .B2(new_n657), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(KEYINPUT97), .A3(new_n702), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n709), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n208), .ZN(G21));
  INV_X1    g530(.A(KEYINPUT99), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n676), .A2(new_n717), .A3(new_n677), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT99), .B1(new_n527), .B2(new_n572), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n434), .B(new_n437), .C1(new_n430), .C2(new_n454), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n414), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT98), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n721), .A2(KEYINPUT98), .A3(new_n414), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n413), .A3(new_n605), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n720), .A2(new_n728), .A3(new_n615), .A4(new_n702), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  AND3_X1   g544(.A1(new_n721), .A2(KEYINPUT98), .A3(new_n414), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT98), .B1(new_n721), .B2(new_n414), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n605), .B(new_n675), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT100), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n726), .A2(new_n735), .A3(new_n605), .A4(new_n675), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n684), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT97), .B1(new_n713), .B2(new_n702), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n288), .A2(new_n710), .A3(new_n711), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NOR2_X1   g555(.A1(new_n658), .A2(new_n674), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n602), .A3(new_n688), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT32), .B1(new_n448), .B2(new_n414), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n744), .B(KEYINPUT101), .Z(new_n745));
  NAND3_X1  g559(.A1(new_n468), .A2(new_n475), .A3(new_n476), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n413), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT42), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n412), .B1(new_n695), .B2(new_n452), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n658), .A2(new_n357), .A3(new_n674), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n684), .A2(KEYINPUT42), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n312), .ZN(G33));
  AND3_X1   g568(.A1(new_n749), .A2(new_n653), .A3(new_n750), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n304), .ZN(G36));
  NAND2_X1  g570(.A1(new_n348), .A2(new_n350), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT102), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n289), .B1(new_n757), .B2(new_n758), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT46), .B1(new_n762), .B2(new_n353), .ZN(new_n763));
  INV_X1    g577(.A(new_n343), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n353), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n597), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n664), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n742), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n572), .A2(new_n682), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT43), .Z(new_n772));
  OAI211_X1 g586(.A(new_n772), .B(new_n675), .C1(new_n603), .C2(new_n630), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n769), .B(new_n775), .C1(new_n774), .C2(new_n773), .ZN(new_n776));
  XOR2_X1   g590(.A(KEYINPUT103), .B(G137), .Z(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(G39));
  XNOR2_X1  g592(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n767), .B1(KEYINPUT104), .B2(new_n781), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n770), .A2(new_n413), .A3(new_n477), .A4(new_n684), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NAND2_X1  g599(.A1(new_n702), .A2(new_n674), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT110), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n662), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n772), .A2(new_n575), .A3(new_n574), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n727), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n787), .A2(new_n662), .A3(KEYINPUT111), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT50), .Z(new_n795));
  NOR3_X1   g609(.A1(new_n672), .A2(new_n412), .A3(new_n576), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n702), .A3(new_n742), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n797), .A2(new_n676), .A3(new_n682), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n791), .A2(new_n711), .A3(new_n770), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n734), .A2(new_n736), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n795), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n701), .A2(new_n343), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n356), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n780), .B2(new_n782), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n742), .B(new_n792), .C1(new_n808), .C2(new_n809), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n805), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT114), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n814));
  INV_X1    g628(.A(new_n715), .ZN(new_n815));
  INV_X1    g629(.A(new_n707), .ZN(new_n816));
  INV_X1    g630(.A(new_n703), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n596), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(new_n816), .A3(new_n818), .A4(new_n729), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n814), .B1(new_n819), .B2(new_n753), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n801), .A2(new_n688), .ZN(new_n821));
  OR4_X1    g635(.A1(new_n557), .A2(new_n626), .A3(new_n677), .A4(new_n687), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n477), .A2(new_n642), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n755), .B1(new_n824), .B2(new_n750), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n611), .A2(new_n582), .A3(new_n643), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT105), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n572), .A2(new_n677), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n615), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT105), .B1(new_n584), .B2(new_n828), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n632), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n825), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n729), .B1(new_n699), .B2(new_n703), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n715), .A3(new_n707), .ZN(new_n836));
  INV_X1    g650(.A(new_n753), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT109), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n820), .A2(new_n834), .A3(new_n838), .A4(KEYINPUT53), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n357), .A2(new_n675), .A3(new_n687), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n720), .A3(new_n713), .A4(new_n672), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n654), .A2(new_n659), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n697), .A2(new_n740), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT107), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n357), .B1(new_n685), .B2(new_n689), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n660), .B1(new_n846), .B2(new_n696), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(KEYINPUT107), .A3(new_n740), .A4(new_n841), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n843), .A2(KEYINPUT52), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n839), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT108), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n845), .A2(new_n848), .A3(KEYINPUT52), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n836), .A2(new_n837), .A3(new_n825), .A4(new_n833), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n853), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n852), .B1(new_n855), .B2(KEYINPUT53), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n845), .A2(new_n848), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n854), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n845), .A2(new_n848), .A3(KEYINPUT52), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(KEYINPUT108), .A3(new_n863), .ZN(new_n864));
  AOI211_X1 g678(.A(KEYINPUT54), .B(new_n851), .C1(new_n856), .C2(new_n864), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n860), .A2(KEYINPUT106), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n860), .A2(KEYINPUT106), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n866), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n849), .A2(new_n850), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n868), .A2(new_n869), .B1(KEYINPUT53), .B2(new_n862), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n865), .B1(KEYINPUT54), .B2(new_n870), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n808), .A2(new_n727), .A3(new_n770), .A4(new_n791), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n804), .B1(new_n872), .B2(new_n803), .ZN(new_n873));
  INV_X1    g687(.A(new_n747), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n800), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT48), .Z(new_n876));
  OAI21_X1  g690(.A(new_n792), .B1(new_n738), .B2(new_n739), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n574), .C1(new_n595), .C2(new_n797), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n813), .A2(new_n871), .A3(new_n873), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n573), .A2(new_n333), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n771), .A2(new_n412), .A3(new_n674), .A4(new_n597), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n806), .B(KEYINPUT49), .Z(new_n884));
  NAND4_X1  g698(.A1(new_n662), .A2(new_n673), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n882), .A2(new_n885), .ZN(G75));
  AOI21_X1  g700(.A(new_n851), .B1(new_n856), .B2(new_n864), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n269), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(G210), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n239), .A2(new_n263), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n261), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n889), .B(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n333), .A2(G952), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT115), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n893), .A2(new_n896), .ZN(G51));
  NOR3_X1   g711(.A1(new_n887), .A2(new_n269), .A3(new_n762), .ZN(new_n898));
  XNOR2_X1  g712(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n352), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n856), .A2(new_n864), .ZN(new_n902));
  INV_X1    g716(.A(new_n851), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n900), .B1(new_n904), .B2(new_n865), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n700), .B(KEYINPUT117), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n898), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT118), .B1(new_n907), .B2(new_n894), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n909));
  INV_X1    g723(.A(new_n894), .ZN(new_n910));
  INV_X1    g724(.A(new_n906), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n855), .A2(new_n852), .A3(KEYINPUT53), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT108), .B1(new_n862), .B2(new_n863), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n887), .A2(new_n901), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n911), .B1(new_n917), .B2(new_n900), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n909), .B(new_n910), .C1(new_n918), .C2(new_n898), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n908), .A2(new_n919), .ZN(G54));
  NAND3_X1  g734(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  INV_X1    g736(.A(new_n623), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n910), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(G60));
  XNOR2_X1  g741(.A(new_n591), .B(KEYINPUT59), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(new_n916), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n586), .A2(new_n588), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n895), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n928), .B1(new_n586), .B2(new_n588), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n917), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(KEYINPUT120), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(KEYINPUT120), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n411), .B1(new_n887), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n939), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n914), .A2(new_n638), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n942), .A3(new_n895), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT121), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n896), .A2(new_n944), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n947), .A2(new_n942), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT121), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n943), .A2(new_n951), .A3(new_n944), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n946), .A2(new_n950), .A3(new_n952), .ZN(G66));
  OAI21_X1  g767(.A(G953), .B1(new_n577), .B2(new_n259), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n836), .A2(new_n833), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n956), .B2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n890), .B1(G898), .B2(new_n333), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT123), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  INV_X1    g774(.A(new_n776), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n961), .A2(new_n753), .A3(new_n755), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n713), .A2(new_n769), .A3(new_n720), .A4(new_n874), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n847), .A2(new_n740), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n962), .A2(new_n333), .A3(new_n784), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n418), .A2(new_n422), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(new_n559), .Z(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(G900), .B2(G953), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n333), .B1(G227), .B2(G900), .ZN(new_n971));
  AOI22_X1  g785(.A1(new_n967), .A2(new_n970), .B1(KEYINPUT124), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n964), .A2(new_n680), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT62), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n595), .A2(new_n828), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n749), .A2(new_n664), .A3(new_n750), .A4(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n974), .A2(new_n784), .A3(new_n776), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n333), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n969), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n971), .A2(KEYINPUT124), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(G72));
  XNOR2_X1  g796(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n467), .A2(new_n269), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n464), .A2(new_n431), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n870), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT127), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n460), .A2(new_n430), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n962), .A2(new_n784), .A3(new_n956), .A4(new_n966), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n990), .A2(KEYINPUT126), .A3(new_n985), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT126), .B1(new_n990), .B2(new_n985), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n985), .B1(new_n977), .B2(new_n955), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n894), .B1(new_n994), .B2(new_n667), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n988), .A2(new_n993), .A3(new_n995), .ZN(G57));
endmodule


