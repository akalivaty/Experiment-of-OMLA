//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT81), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211));
  INV_X1    g010(.A(G1gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT16), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT86), .B1(new_n211), .B2(G1gat), .ZN(new_n216));
  OAI21_X1  g015(.A(G8gat), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n211), .A2(G1gat), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n218), .A2(new_n214), .A3(KEYINPUT86), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G43gat), .A2(G50gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G43gat), .A2(G50gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT15), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT83), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT83), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(KEYINPUT15), .C1(new_n223), .C2(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230));
  AND2_X1   g029(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n231), .A2(new_n232), .A3(G50gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(G43gat), .A2(G50gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT15), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n230), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G29gat), .ZN(new_n238));
  INV_X1    g037(.A(G36gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT14), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT14), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G29gat), .B2(G36gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(G29gat), .A2(G36gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n236), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT84), .B(G43gat), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n246), .B(KEYINPUT85), .C1(new_n247), .C2(G50gat), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n229), .A2(new_n237), .A3(new_n245), .A4(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G43gat), .ZN(new_n250));
  INV_X1    g049(.A(G50gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n235), .B1(new_n252), .B2(new_n234), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n244), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n244), .A2(new_n253), .A3(KEYINPUT82), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n249), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n249), .B2(new_n258), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n222), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n249), .A2(new_n258), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(new_n221), .B1(G229gat), .B2(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n210), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AOI211_X1 g067(.A(KEYINPUT88), .B(new_n266), .C1(new_n262), .C2(new_n264), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT89), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n263), .A2(KEYINPUT17), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n249), .A2(new_n258), .A3(new_n259), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n221), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n263), .A2(new_n221), .ZN(new_n275));
  NAND2_X1  g074(.A1(G229gat), .A2(G233gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(KEYINPUT18), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n262), .A2(KEYINPUT89), .A3(KEYINPUT18), .A4(new_n264), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n263), .B(new_n221), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n276), .B(KEYINPUT13), .Z(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n209), .B1(new_n270), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n286));
  INV_X1    g085(.A(new_n264), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n267), .B1(new_n274), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n207), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT24), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n297), .A2(new_n298), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(KEYINPUT24), .A3(new_n296), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n295), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT27), .B(G183gat), .Z(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n307), .A2(new_n308), .A3(G190gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT27), .B1(new_n300), .B2(KEYINPUT64), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n300), .A2(KEYINPUT27), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n301), .B(new_n310), .C1(new_n311), .C2(KEYINPUT64), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n309), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n297), .B1(KEYINPUT26), .B2(new_n293), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT26), .ZN(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n314), .B1(new_n293), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n306), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT68), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n325), .A3(new_n322), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n304), .B(KEYINPUT25), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n313), .A2(new_n319), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(KEYINPUT65), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT65), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n313), .B2(new_n319), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT29), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n324), .B(new_n326), .C1(new_n332), .C2(new_n322), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT22), .ZN(new_n335));
  INV_X1    g134(.A(G211gat), .ZN(new_n336));
  INV_X1    g135(.A(G218gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G211gat), .B(G218gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT67), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n333), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n322), .A3(new_n331), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n320), .A2(new_n346), .A3(new_n321), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n341), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G8gat), .B(G36gat), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT69), .ZN(new_n352));
  XNOR2_X1  g151(.A(G64gat), .B(G92gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  NAND2_X1  g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n348), .B1(new_n333), .B2(new_n343), .ZN(new_n356));
  INV_X1    g155(.A(new_n354), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(new_n358), .A3(KEYINPUT30), .ZN(new_n359));
  INV_X1    g158(.A(new_n358), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT30), .B1(new_n356), .B2(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G141gat), .B(G148gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(G155gat), .B2(G162gat), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT70), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G155gat), .B(G162gat), .Z(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G113gat), .B(G120gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(KEYINPUT1), .ZN(new_n371));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n371), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n369), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT5), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n369), .A2(new_n374), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT4), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n367), .B(new_n368), .Z(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n369), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n384), .A3(new_n375), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n377), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n378), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n380), .A2(KEYINPUT5), .A3(new_n377), .A4(new_n385), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G1gat), .B(G29gat), .Z(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT71), .B(KEYINPUT0), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT6), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n395), .B2(new_n390), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n390), .A2(new_n395), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT6), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n363), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n346), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n342), .B1(KEYINPUT74), .B2(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n402), .A2(KEYINPUT74), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n340), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n339), .B(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT3), .B1(new_n407), .B2(new_n346), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(new_n369), .ZN(new_n409));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(KEYINPUT72), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n402), .A2(new_n341), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT72), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n408), .B2(new_n369), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT73), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(new_n410), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n417), .B2(new_n410), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n412), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT31), .B(G50gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(G22gat), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(KEYINPUT76), .ZN(new_n428));
  XOR2_X1   g227(.A(KEYINPUT75), .B(G22gat), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n422), .B2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n412), .B(new_n429), .C1(new_n420), .C2(new_n421), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n422), .A2(new_n430), .A3(new_n428), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n427), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G71gat), .B(G99gat), .Z(new_n437));
  XNOR2_X1  g236(.A(G15gat), .B(G43gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT66), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n440), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(KEYINPUT33), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n328), .A2(KEYINPUT65), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n331), .A3(new_n306), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n375), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n329), .A2(new_n374), .A3(new_n331), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G227gat), .A2(G233gat), .ZN(new_n449));
  OAI211_X1 g248(.A(KEYINPUT32), .B(new_n443), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n446), .B2(new_n447), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT32), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n439), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n451), .A2(KEYINPUT33), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n446), .A2(new_n449), .A3(new_n447), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT34), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n455), .B(new_n457), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n401), .A2(new_n436), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT35), .ZN(new_n460));
  INV_X1    g259(.A(new_n427), .ZN(new_n461));
  INV_X1    g260(.A(new_n428), .ZN(new_n462));
  INV_X1    g261(.A(new_n421), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n463), .A2(new_n419), .B1(new_n405), .B2(new_n411), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n464), .B2(new_n429), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n432), .ZN(new_n466));
  INV_X1    g265(.A(new_n435), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n456), .B(KEYINPUT34), .Z(new_n469));
  XNOR2_X1  g268(.A(new_n455), .B(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n363), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT79), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n388), .A2(KEYINPUT78), .A3(new_n389), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT78), .B1(new_n388), .B2(new_n389), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n473), .A2(new_n474), .A3(new_n395), .ZN(new_n475));
  INV_X1    g274(.A(new_n396), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT78), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n395), .B1(new_n390), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n388), .A2(KEYINPUT78), .A3(new_n389), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(KEYINPUT79), .A3(new_n396), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n399), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n460), .ZN(new_n484));
  OAI22_X1  g283(.A1(new_n459), .A2(new_n460), .B1(new_n471), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n386), .A2(new_n387), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n376), .B2(new_n377), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n386), .A2(new_n487), .A3(new_n387), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT77), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n490), .A2(new_n491), .A3(new_n395), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n490), .B2(new_n395), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT40), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n494), .A2(new_n495), .B1(new_n479), .B2(new_n480), .ZN(new_n496));
  OAI211_X1 g295(.A(KEYINPUT40), .B(new_n489), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n496), .A2(new_n362), .A3(new_n359), .A4(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n357), .B1(new_n356), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n345), .A2(new_n341), .A3(new_n347), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n333), .B2(new_n343), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT38), .B1(new_n502), .B2(KEYINPUT37), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n360), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n354), .B1(new_n350), .B2(KEYINPUT37), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n356), .A2(new_n499), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT38), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n468), .B(new_n498), .C1(new_n483), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n401), .A2(new_n436), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n470), .A2(KEYINPUT36), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n458), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n292), .B1(new_n485), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n263), .ZN(new_n518));
  NAND2_X1  g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT92), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(G99gat), .A3(G106gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT8), .ZN(new_n523));
  OAI21_X1  g322(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n524));
  AND2_X1   g323(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527));
  INV_X1    g326(.A(G85gat), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n527), .A2(new_n528), .A3(G92gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n523), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G99gat), .B(G106gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n523), .B(new_n531), .C1(new_n529), .C2(new_n526), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n517), .B1(new_n518), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n272), .A2(new_n273), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n535), .ZN(new_n538));
  XOR2_X1   g337(.A(G190gat), .B(G218gat), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT93), .ZN(new_n541));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n538), .A2(new_n539), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n540), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n541), .A2(new_n546), .A3(new_n540), .A4(new_n544), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(G57gat), .A2(G64gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(G57gat), .A2(G64gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT90), .ZN(new_n557));
  NAND2_X1  g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n553), .A2(new_n556), .A3(new_n557), .A4(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(G57gat), .A2(G64gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(G57gat), .A2(G64gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(new_n557), .A3(new_n558), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT90), .B1(new_n551), .B2(new_n552), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n535), .A2(new_n561), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n561), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n533), .A2(new_n570), .A3(new_n534), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(KEYINPUT94), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n571), .A2(KEYINPUT94), .A3(KEYINPUT10), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n569), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n575), .B1(new_n580), .B2(new_n574), .ZN(new_n581));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT96), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n579), .A2(new_n569), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT10), .B1(new_n571), .B2(KEYINPUT94), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n578), .A2(KEYINPUT95), .A3(new_n569), .A4(new_n579), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n573), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n575), .A3(new_n584), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n570), .A2(KEYINPUT21), .ZN(new_n597));
  XOR2_X1   g396(.A(G127gat), .B(G155gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n221), .B1(KEYINPUT21), .B2(new_n570), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT91), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n601), .B(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n550), .A2(new_n596), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT97), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n516), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n400), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n212), .ZN(G1324gat));
  INV_X1    g412(.A(new_n611), .ZN(new_n614));
  INV_X1    g413(.A(new_n363), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n219), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT16), .B(G8gat), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n611), .A2(new_n363), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT42), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(KEYINPUT42), .B2(new_n618), .ZN(G1325gat));
  OAI21_X1  g419(.A(G15gat), .B1(new_n611), .B2(new_n514), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n458), .A2(G15gat), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n621), .B1(new_n611), .B2(new_n622), .ZN(G1326gat));
  NOR2_X1   g422(.A1(new_n611), .A2(new_n468), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT43), .B(G22gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(G1327gat));
  INV_X1    g425(.A(new_n608), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n596), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n550), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n516), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n400), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n238), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT45), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n485), .A2(new_n515), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n548), .A2(new_n549), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT44), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n286), .A2(new_n289), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT98), .B1(new_n284), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n286), .A2(new_n268), .A3(new_n269), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n290), .B(new_n641), .C1(new_n642), .C2(new_n209), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n550), .B1(new_n485), .B2(new_n515), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT99), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n359), .A2(new_n362), .B1(new_n397), .B2(new_n399), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT100), .B1(new_n468), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n401), .A2(new_n436), .A3(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n509), .A2(new_n650), .A3(new_n514), .A4(new_n652), .ZN(new_n653));
  AOI211_X1 g452(.A(KEYINPUT44), .B(new_n550), .C1(new_n485), .C2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n638), .B(new_n645), .C1(new_n648), .C2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(G29gat), .B1(new_n655), .B2(new_n400), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n633), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1328gat));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660));
  AOI21_X1  g459(.A(G36gat), .B1(new_n660), .B2(KEYINPUT46), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n630), .A2(new_n615), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n660), .A2(KEYINPUT46), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G36gat), .B1(new_n655), .B2(new_n363), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT103), .ZN(G1329gat));
  OAI21_X1  g466(.A(new_n247), .B1(new_n655), .B2(new_n514), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT47), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n458), .A2(new_n247), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n630), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n670), .B(new_n673), .ZN(G1330gat));
  OAI21_X1  g473(.A(G50gat), .B1(new_n655), .B2(new_n468), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n630), .A2(new_n251), .A3(new_n436), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT48), .Z(G1331gat));
  NAND4_X1  g477(.A1(new_n644), .A2(new_n550), .A3(new_n608), .A4(new_n595), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n485), .B2(new_n653), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n631), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G57gat), .ZN(G1332gat));
  INV_X1    g481(.A(KEYINPUT49), .ZN(new_n683));
  INV_X1    g482(.A(G64gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n615), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT105), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1333gat));
  INV_X1    g488(.A(new_n514), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n680), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n458), .A2(G71gat), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n691), .A2(G71gat), .B1(new_n680), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1334gat));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n436), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g496(.A1(new_n644), .A2(new_n627), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n596), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT107), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n638), .B(new_n700), .C1(new_n648), .C2(new_n654), .ZN(new_n701));
  OAI21_X1  g500(.A(G85gat), .B1(new_n701), .B2(new_n400), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n485), .A2(new_n653), .ZN(new_n703));
  INV_X1    g502(.A(new_n698), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n635), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n707), .A2(new_n528), .A3(new_n631), .A4(new_n595), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT108), .ZN(G1336gat));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n550), .B(new_n698), .C1(new_n485), .C2(new_n653), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(KEYINPUT51), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n706), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n703), .A2(new_n714), .A3(new_n635), .A4(new_n704), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n713), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n363), .A2(G92gat), .A3(new_n596), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT51), .B1(new_n705), .B2(KEYINPUT109), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n711), .A3(new_n716), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G92gat), .B1(new_n701), .B2(new_n363), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT52), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT52), .B1(new_n707), .B2(new_n719), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(KEYINPUT111), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n722), .B2(new_n723), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n723), .A2(new_n726), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n733), .ZN(G1337gat));
  XNOR2_X1  g533(.A(KEYINPUT112), .B(G99gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n707), .A2(new_n470), .A3(new_n595), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n701), .A2(new_n514), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n735), .ZN(G1338gat));
  NOR3_X1   g537(.A1(new_n468), .A2(G106gat), .A3(new_n596), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n718), .A2(new_n721), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G106gat), .B1(new_n701), .B2(new_n468), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT53), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT53), .B1(new_n707), .B2(new_n739), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1339gat));
  INV_X1    g545(.A(KEYINPUT54), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n580), .B2(new_n574), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n593), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n589), .A2(new_n590), .A3(new_n574), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n584), .B1(new_n750), .B2(new_n747), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(KEYINPUT55), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n594), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT55), .B1(new_n749), .B2(new_n751), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n640), .A2(new_n755), .A3(new_n643), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n280), .A2(KEYINPUT113), .A3(new_n281), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT113), .B1(new_n280), .B2(new_n281), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n262), .A2(new_n275), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n757), .B(new_n758), .C1(new_n276), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n206), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n595), .A2(new_n290), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n635), .B1(new_n756), .B2(new_n762), .ZN(new_n763));
  AND4_X1   g562(.A1(new_n290), .A2(new_n635), .A3(new_n755), .A4(new_n761), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n627), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n644), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n609), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n765), .A2(new_n771), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n436), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n615), .A2(new_n458), .A3(new_n400), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(G113gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n776), .A2(new_n777), .A3(new_n292), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n773), .A2(new_n400), .ZN(new_n779));
  INV_X1    g578(.A(new_n471), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n780), .A3(new_n766), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n778), .B1(new_n777), .B2(new_n781), .ZN(G1340gat));
  OAI21_X1  g581(.A(G120gat), .B1(new_n776), .B2(new_n596), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT115), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n780), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n596), .A2(G120gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(G1341gat));
  OAI21_X1  g586(.A(G127gat), .B1(new_n776), .B2(new_n627), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n627), .A2(G127gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n785), .B2(new_n789), .ZN(G1342gat));
  NOR3_X1   g589(.A1(new_n785), .A2(G134gat), .A3(new_n550), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT116), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n774), .A2(new_n635), .A3(new_n775), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n791), .A2(new_n792), .B1(G134gat), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1343gat));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n514), .A2(new_n363), .A3(new_n436), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n773), .A2(new_n400), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(G141gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n801), .A3(new_n291), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n436), .A2(KEYINPUT57), .ZN(new_n803));
  INV_X1    g602(.A(new_n753), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n749), .A2(new_n751), .ZN(new_n805));
  XNOR2_X1  g604(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n804), .B(new_n807), .C1(new_n639), .C2(new_n284), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n635), .B1(new_n808), .B2(new_n762), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n627), .B1(new_n809), .B2(new_n764), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n767), .B1(new_n810), .B2(KEYINPUT118), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n627), .C1(new_n809), .C2(new_n764), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n803), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n770), .A2(new_n436), .A3(new_n772), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n615), .A2(new_n400), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n514), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n817), .A2(new_n292), .A3(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n798), .B(new_n802), .C1(new_n820), .C2(new_n801), .ZN(new_n821));
  INV_X1    g620(.A(new_n802), .ZN(new_n822));
  INV_X1    g621(.A(new_n814), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n765), .A2(new_n768), .A3(new_n771), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n771), .B1(new_n765), .B2(new_n768), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n824), .A2(new_n825), .A3(new_n468), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n826), .B2(KEYINPUT57), .ZN(new_n827));
  INV_X1    g626(.A(new_n819), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(KEYINPUT119), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n817), .B2(new_n819), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n831), .A3(new_n766), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n822), .B1(new_n832), .B2(G141gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n821), .B1(new_n833), .B2(new_n798), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n821), .B(KEYINPUT120), .C1(new_n833), .C2(new_n798), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1344gat));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n839), .B(G148gat), .C1(new_n800), .C2(new_n595), .ZN(new_n840));
  INV_X1    g639(.A(G148gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n610), .A2(new_n292), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(new_n810), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n816), .B1(new_n843), .B2(new_n468), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n773), .B2(new_n803), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n595), .A3(new_n828), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n841), .B1(new_n846), .B2(KEYINPUT59), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n829), .A2(new_n831), .A3(new_n839), .A4(new_n595), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n840), .B1(new_n847), .B2(new_n848), .ZN(G1345gat));
  NAND2_X1  g648(.A1(new_n829), .A2(new_n831), .ZN(new_n850));
  OAI21_X1  g649(.A(G155gat), .B1(new_n850), .B2(new_n627), .ZN(new_n851));
  INV_X1    g650(.A(new_n800), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n627), .A2(G155gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(G1346gat));
  NOR3_X1   g653(.A1(new_n852), .A2(G162gat), .A3(new_n550), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT121), .Z(new_n856));
  OAI21_X1  g655(.A(G162gat), .B1(new_n850), .B2(new_n550), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1347gat));
  NAND2_X1  g657(.A1(new_n615), .A2(new_n400), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n458), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n774), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(new_n316), .A3(new_n292), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n773), .A2(new_n631), .ZN(new_n863));
  AND4_X1   g662(.A1(new_n615), .A2(new_n863), .A3(new_n468), .A4(new_n470), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n766), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n862), .B1(new_n316), .B2(new_n865), .ZN(G1348gat));
  AOI21_X1  g665(.A(G176gat), .B1(new_n864), .B2(new_n595), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n774), .A2(G176gat), .A3(new_n595), .A4(new_n860), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(KEYINPUT122), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(KEYINPUT122), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(G1349gat));
  NOR2_X1   g670(.A1(new_n627), .A2(new_n307), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G183gat), .B1(new_n861), .B2(new_n627), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(KEYINPUT123), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n875), .B2(KEYINPUT60), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n881), .B1(new_n876), .B2(new_n877), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n875), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n883));
  OAI22_X1  g682(.A1(new_n878), .A2(new_n880), .B1(new_n882), .B2(new_n883), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n861), .B2(new_n550), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT61), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n864), .A2(new_n301), .A3(new_n635), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1351gat));
  NAND4_X1  g687(.A1(new_n863), .A2(new_n615), .A3(new_n436), .A4(new_n514), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(G197gat), .A3(new_n644), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n690), .A2(new_n859), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n845), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n291), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n890), .B1(new_n894), .B2(G197gat), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n895), .B(new_n896), .ZN(G1352gat));
  INV_X1    g696(.A(G204gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n595), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n900), .B2(new_n899), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n889), .A2(G204gat), .A3(new_n596), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT62), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1353gat));
  OAI21_X1  g704(.A(G211gat), .B1(new_n892), .B2(new_n627), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT63), .B(G211gat), .C1(new_n892), .C2(new_n627), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(KEYINPUT127), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n608), .A2(new_n336), .ZN(new_n911));
  OAI221_X1 g710(.A(new_n910), .B1(KEYINPUT127), .B2(new_n908), .C1(new_n889), .C2(new_n911), .ZN(G1354gat));
  OAI21_X1  g711(.A(G218gat), .B1(new_n892), .B2(new_n550), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n635), .A2(new_n337), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n889), .B2(new_n914), .ZN(G1355gat));
endmodule


