//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n215), .A2(KEYINPUT65), .A3(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI22_X1  g0021(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G116), .ZN(new_n225));
  INV_X1    g0025(.A(G270), .ZN(new_n226));
  OAI22_X1  g0026(.A1(new_n223), .A2(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n217), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(KEYINPUT65), .B1(new_n215), .B2(new_n216), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n205), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n208), .B1(new_n212), .B2(new_n213), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n223), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n218), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT80), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n254), .B(G45), .C1(new_n255), .C2(KEYINPUT5), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT5), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G41), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n253), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n251), .B1(new_n259), .B2(new_n226), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n265), .A2(KEYINPUT80), .A3(G270), .A4(new_n253), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  INV_X1    g0068(.A(new_n209), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(new_n252), .ZN(new_n270));
  INV_X1    g0070(.A(new_n256), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT73), .B1(new_n257), .B2(G41), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT73), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(new_n255), .A3(KEYINPUT5), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n270), .A2(new_n271), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  OAI211_X1 g0077(.A(G264), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  OAI211_X1 g0079(.A(G257), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n280));
  INV_X1    g0080(.A(G303), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n278), .B(new_n280), .C1(new_n281), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n253), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n267), .A2(new_n275), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n225), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n291), .B(new_n209), .C1(new_n283), .C2(new_n205), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT72), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n283), .B2(G1), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n254), .A2(KEYINPUT72), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n292), .B1(new_n298), .B2(new_n225), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G283), .ZN(new_n300));
  INV_X1    g0100(.A(G97), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n300), .B(new_n210), .C1(G33), .C2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n209), .B1(new_n205), .B2(new_n283), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n225), .A2(G20), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT20), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT20), .A4(new_n304), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(KEYINPUT81), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT81), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(new_n310), .A3(new_n306), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n299), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n290), .A2(new_n312), .A3(G169), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT21), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n290), .A2(G200), .ZN(new_n316));
  INV_X1    g0116(.A(new_n312), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n272), .A2(new_n274), .A3(new_n263), .A4(new_n262), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n253), .A2(G274), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n288), .B2(new_n287), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n322), .A2(KEYINPUT70), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(KEYINPUT70), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n321), .B(new_n267), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n316), .A2(new_n317), .A3(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n312), .A2(G179), .A3(new_n267), .A4(new_n321), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n290), .A2(new_n312), .A3(KEYINPUT21), .A4(G169), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n315), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT82), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n328), .A2(new_n327), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT82), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n331), .A2(new_n332), .A3(new_n315), .A4(new_n326), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n286), .A2(G222), .A3(new_n279), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n286), .A2(G1698), .ZN(new_n336));
  INV_X1    g0136(.A(G223), .ZN(new_n337));
  OAI221_X1 g0137(.A(new_n335), .B1(new_n220), .B2(new_n286), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n288), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n253), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT66), .B(G226), .Z(new_n343));
  INV_X1    g0143(.A(new_n340), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n342), .A2(new_n343), .B1(new_n270), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT67), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT67), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n339), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G190), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(G200), .A3(new_n349), .ZN(new_n352));
  INV_X1    g0152(.A(new_n291), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(new_n303), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n254), .A2(G20), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G50), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(G50), .B2(new_n291), .ZN(new_n357));
  INV_X1    g0157(.A(new_n303), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n210), .A2(new_n283), .ZN(new_n359));
  INV_X1    g0159(.A(G150), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT8), .B(G58), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n283), .A2(G20), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n358), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT9), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n351), .A2(new_n352), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT10), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n351), .A2(new_n372), .A3(new_n369), .A4(new_n352), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G179), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n350), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G169), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n347), .A2(new_n377), .A3(new_n349), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n376), .A2(new_n378), .A3(new_n368), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n359), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n383));
  INV_X1    g0183(.A(new_n364), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n220), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(KEYINPUT11), .A3(new_n303), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n353), .A2(new_n218), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT12), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n354), .A2(G68), .A3(new_n355), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT11), .B1(new_n385), .B2(new_n303), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(G226), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT68), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT68), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n286), .A2(new_n395), .A3(G226), .A4(new_n279), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(G232), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n253), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n344), .A2(new_n253), .A3(G274), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n219), .B2(new_n341), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT13), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  INV_X1    g0206(.A(new_n404), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n400), .B1(new_n396), .B2(new_n394), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n406), .B(new_n407), .C1(new_n408), .C2(new_n253), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(G169), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n405), .A2(new_n409), .A3(G179), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n410), .B2(G169), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n392), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n405), .A2(new_n409), .A3(G190), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT69), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT69), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n405), .A2(new_n409), .A3(new_n419), .A4(G190), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G200), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n405), .B2(new_n409), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n392), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n284), .A2(new_n210), .A3(new_n285), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT7), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n284), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n285), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n218), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G58), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(new_n218), .ZN(new_n434));
  OAI21_X1  g0234(.A(G20), .B1(new_n434), .B2(new_n201), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n382), .A2(G159), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n427), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n276), .A2(new_n277), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT7), .B1(new_n439), .B2(new_n210), .ZN(new_n440));
  INV_X1    g0240(.A(new_n431), .ZN(new_n441));
  OAI21_X1  g0241(.A(G68), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n437), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(KEYINPUT16), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n438), .A2(new_n444), .A3(new_n303), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n362), .B1(new_n254), .B2(G20), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(new_n354), .B1(new_n353), .B2(new_n362), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n253), .A2(G232), .A3(new_n340), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n403), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n337), .A2(new_n279), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n224), .A2(G1698), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n451), .B(new_n452), .C1(new_n276), .C2(new_n277), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G87), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n253), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G179), .ZN(new_n457));
  OAI21_X1  g0257(.A(G169), .B1(new_n450), .B2(new_n455), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n448), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT18), .ZN(new_n461));
  INV_X1    g0261(.A(new_n447), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n432), .A2(new_n437), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n358), .B1(new_n463), .B2(KEYINPUT16), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(new_n438), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n323), .A2(new_n324), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n456), .A2(KEYINPUT71), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n453), .A2(new_n454), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n288), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(new_n466), .A3(new_n403), .A4(new_n449), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT71), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n422), .B1(new_n450), .B2(new_n455), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n465), .A2(KEYINPUT17), .A3(new_n467), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT18), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n448), .A2(new_n459), .A3(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n445), .A2(new_n473), .A3(new_n447), .A4(new_n467), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT17), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n461), .A2(new_n474), .A3(new_n476), .A4(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n363), .A2(new_n382), .B1(G20), .B2(G77), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT15), .B(G87), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n364), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n358), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n354), .A2(G77), .A3(new_n355), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G77), .B2(new_n291), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n403), .B1(new_n221), .B2(new_n341), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n286), .A2(G232), .A3(new_n279), .ZN(new_n491));
  INV_X1    g0291(.A(G107), .ZN(new_n492));
  OAI221_X1 g0292(.A(new_n491), .B1(new_n492), .B2(new_n286), .C1(new_n336), .C2(new_n219), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n493), .B2(new_n288), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n375), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n489), .B(new_n495), .C1(G169), .C2(new_n494), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(G190), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(new_n488), .C1(new_n422), .C2(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR4_X1   g0299(.A1(new_n381), .A2(new_n426), .A3(new_n480), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT74), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n265), .A2(G257), .A3(new_n253), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n503), .B2(new_n320), .ZN(new_n504));
  OAI211_X1 g0304(.A(G250), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n300), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n288), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n275), .A2(KEYINPUT74), .A3(new_n502), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n504), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G200), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n291), .A2(G97), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n298), .B2(G97), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(G107), .B1(new_n440), .B2(new_n441), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n301), .A2(new_n492), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n492), .A2(KEYINPUT6), .A3(G97), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n382), .A2(G77), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n517), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n516), .B1(new_n526), .B2(new_n303), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n513), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n275), .A2(KEYINPUT74), .A3(new_n502), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT74), .B1(new_n275), .B2(new_n502), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT75), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(G190), .A4(new_n510), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT75), .B1(new_n512), .B2(new_n322), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n528), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(new_n375), .A3(new_n510), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n512), .A2(new_n377), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n526), .A2(new_n303), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n515), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G238), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n541));
  OAI211_X1 g0341(.A(G244), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G116), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT76), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT76), .A4(new_n543), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n288), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n262), .A2(G250), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n288), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n262), .A2(new_n268), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n377), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n253), .B1(new_n544), .B2(new_n545), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n547), .B1(new_n551), .B2(new_n550), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n375), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n483), .A2(new_n291), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n286), .A2(new_n210), .A3(G68), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n384), .B2(new_n301), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n210), .B1(new_n399), .B2(new_n560), .ZN(new_n562));
  INV_X1    g0362(.A(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n520), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT77), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT77), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n559), .B(new_n561), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n558), .B1(new_n567), .B2(new_n303), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT79), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n482), .B(KEYINPUT78), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n354), .A2(new_n296), .A3(new_n295), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT78), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n482), .B(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(KEYINPUT79), .A3(new_n298), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n568), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n554), .A2(new_n557), .A3(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n293), .A2(new_n297), .A3(new_n563), .ZN(new_n578));
  AOI211_X1 g0378(.A(new_n558), .B(new_n578), .C1(new_n567), .C2(new_n303), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n548), .A2(G190), .A3(new_n552), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n579), .B(new_n580), .C1(new_n422), .C2(new_n556), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n535), .A2(new_n540), .A3(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(G257), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n584));
  OAI211_X1 g0384(.A(G250), .B(new_n279), .C1(new_n276), .C2(new_n277), .ZN(new_n585));
  INV_X1    g0385(.A(G294), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n584), .B(new_n585), .C1(new_n283), .C2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n259), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n288), .B1(new_n588), .B2(G264), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT85), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n589), .A2(new_n590), .A3(G179), .A4(new_n275), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n210), .B(G87), .C1(new_n276), .C2(new_n277), .ZN(new_n592));
  XNOR2_X1  g0392(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT22), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n595), .A2(KEYINPUT83), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n286), .A2(new_n210), .A3(G87), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT84), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n598), .B(KEYINPUT23), .C1(new_n210), .C2(G107), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT23), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(new_n492), .A3(G20), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT84), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n594), .A2(new_n597), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT24), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n605), .A2(new_n599), .A3(new_n600), .A4(new_n602), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT24), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n597), .A4(new_n594), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n358), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n291), .A2(G107), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(KEYINPUT25), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n492), .B2(new_n571), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n591), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n587), .A2(new_n288), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n588), .A2(G264), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n616), .A2(G179), .A3(new_n617), .A4(new_n275), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT85), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n377), .B1(new_n589), .B2(new_n275), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n616), .A2(new_n275), .A3(new_n617), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n589), .A2(G190), .A3(new_n275), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n626), .A2(new_n611), .A3(new_n614), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT86), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  OAI221_X1 g0428(.A(new_n591), .B1(new_n611), .B2(new_n614), .C1(new_n620), .C2(new_n619), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT86), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n611), .A2(new_n614), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n625), .A3(new_n624), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n334), .A2(new_n500), .A3(new_n583), .A4(new_n634), .ZN(G372));
  NAND3_X1  g0435(.A1(new_n629), .A2(new_n315), .A3(new_n331), .ZN(new_n636));
  INV_X1    g0436(.A(new_n528), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n534), .A2(new_n533), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n377), .A2(new_n512), .B1(new_n538), .B2(new_n515), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n637), .A2(new_n638), .B1(new_n536), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n582), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n636), .A2(new_n640), .A3(new_n641), .A4(new_n632), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n639), .A2(new_n536), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n582), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n540), .A2(KEYINPUT26), .A3(new_n577), .A4(new_n581), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(KEYINPUT87), .B(new_n643), .C1(new_n582), .C2(new_n644), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n642), .A2(new_n648), .A3(new_n577), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n500), .A2(new_n650), .ZN(new_n651));
  AOI211_X1 g0451(.A(new_n392), .B(new_n423), .C1(new_n418), .C2(new_n420), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n416), .B1(new_n652), .B2(new_n496), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(new_n479), .A3(new_n474), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(new_n461), .A3(new_n476), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n379), .B1(new_n655), .B2(new_n374), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n656), .ZN(G369));
  NAND3_X1  g0457(.A1(new_n254), .A2(new_n210), .A3(G13), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n658), .A2(KEYINPUT88), .A3(KEYINPUT27), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT88), .B1(new_n658), .B2(KEYINPUT27), .ZN(new_n660));
  OAI221_X1 g0460(.A(G213), .B1(KEYINPUT27), .B2(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n312), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n334), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n331), .A2(new_n315), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n664), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(KEYINPUT89), .A3(G330), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT89), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n665), .A2(new_n667), .ZN(new_n671));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n663), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n634), .B1(new_n631), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n622), .A2(new_n663), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n666), .A2(new_n663), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n633), .B2(new_n628), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n622), .B2(new_n676), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n206), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n254), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n564), .A2(G116), .ZN(new_n689));
  INV_X1    g0489(.A(new_n213), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n688), .A2(new_n689), .B1(new_n690), .B2(new_n687), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT28), .Z(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n531), .A2(new_n556), .A3(new_n510), .A4(new_n589), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n321), .A2(G179), .A3(new_n267), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AND4_X1   g0496(.A1(new_n510), .A2(new_n504), .A3(new_n589), .A4(new_n511), .ZN(new_n697));
  INV_X1    g0497(.A(new_n695), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(KEYINPUT30), .A4(new_n556), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n290), .A2(new_n623), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n375), .A3(new_n512), .A4(new_n553), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n663), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT31), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(new_n703), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n634), .A2(new_n334), .A3(new_n583), .A4(new_n676), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n672), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n650), .A2(new_n676), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n645), .A2(new_n647), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n642), .A2(new_n577), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n709), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n692), .B1(new_n716), .B2(G1), .ZN(G364));
  NAND2_X1  g0517(.A1(new_n210), .A2(G13), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT91), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G45), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n688), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n668), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n686), .A2(new_n439), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n728), .A2(G355), .B1(new_n225), .B2(new_n686), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n249), .A2(new_n261), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n686), .A2(new_n286), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G45), .B2(new_n213), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT92), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(KEYINPUT92), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n209), .B1(G20), .B2(new_n377), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n725), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n210), .A2(new_n375), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G190), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n422), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G190), .ZN(new_n743));
  AOI22_X1  g0543(.A1(G68), .A2(new_n741), .B1(new_n743), .B2(G77), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n466), .A2(new_n742), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n744), .B1(new_n433), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n210), .A2(G190), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n375), .A3(G200), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT94), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT94), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G107), .ZN(new_n754));
  NOR4_X1   g0554(.A1(new_n210), .A2(new_n322), .A3(new_n422), .A4(G179), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n439), .B1(new_n755), .B2(G87), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n466), .A2(new_n740), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n754), .B(new_n756), .C1(new_n223), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n375), .A2(new_n422), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT93), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n210), .B1(new_n762), .B2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n747), .B(new_n759), .C1(G97), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n748), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n757), .A2(G326), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n286), .B1(new_n755), .B2(G303), .ZN(new_n771));
  INV_X1    g0571(.A(G329), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n770), .B(new_n771), .C1(new_n766), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(G283), .B2(new_n753), .ZN(new_n774));
  INV_X1    g0574(.A(G317), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT33), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(KEYINPUT33), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n741), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n743), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n778), .B1(new_n779), .B2(new_n780), .C1(new_n746), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G294), .B2(new_n764), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n765), .A2(new_n769), .B1(new_n774), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n736), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n738), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n722), .B1(new_n727), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n674), .B1(new_n672), .B2(new_n671), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n722), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT95), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  INV_X1    g0591(.A(KEYINPUT99), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n489), .A2(new_n663), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n496), .A2(new_n498), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT97), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT97), .A4(new_n793), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT98), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n496), .B2(new_n676), .ZN(new_n799));
  INV_X1    g0599(.A(new_n494), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n488), .B1(new_n800), .B2(new_n377), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n801), .A2(KEYINPUT98), .A3(new_n495), .A4(new_n663), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n796), .A2(new_n797), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n710), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n709), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n792), .B1(new_n806), .B2(new_n721), .ZN(new_n807));
  AOI211_X1 g0607(.A(KEYINPUT99), .B(new_n722), .C1(new_n805), .C2(new_n709), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(new_n709), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n785), .A2(new_n724), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n722), .B1(G77), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT96), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n757), .A2(G303), .B1(new_n743), .B2(G116), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n814), .B1(new_n586), .B2(new_n746), .C1(new_n763), .C2(new_n301), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n752), .A2(new_n563), .ZN(new_n816));
  INV_X1    g0616(.A(new_n741), .ZN(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n755), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n439), .B1(new_n820), .B2(new_n492), .ZN(new_n821));
  OR3_X1    g0621(.A1(new_n816), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n766), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n815), .B(new_n822), .C1(G311), .C2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n745), .A2(G143), .B1(new_n741), .B2(G150), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n825), .B1(new_n826), .B2(new_n758), .C1(new_n767), .C2(new_n779), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT34), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(G132), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n753), .A2(G68), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n439), .B1(new_n755), .B2(G50), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G58), .B2(new_n764), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n824), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n813), .B1(new_n785), .B2(new_n834), .C1(new_n804), .C2(new_n724), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT100), .B1(new_n810), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n806), .A2(new_n721), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n809), .B1(new_n838), .B2(KEYINPUT99), .ZN(new_n839));
  INV_X1    g0639(.A(new_n808), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT100), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(new_n835), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n837), .A2(new_n843), .ZN(G384));
  NOR2_X1   g0644(.A1(new_n719), .A2(new_n254), .ZN(new_n845));
  INV_X1    g0645(.A(new_n661), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT103), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n432), .B2(new_n437), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n442), .A2(KEYINPUT103), .A3(new_n443), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n849), .A3(new_n427), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n464), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n447), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n480), .A2(new_n846), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT104), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n846), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n852), .A2(new_n459), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n477), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n854), .B1(new_n857), .B2(KEYINPUT37), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n462), .B1(new_n850), .B2(new_n464), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n477), .B1(new_n859), .B2(new_n661), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n851), .A2(new_n447), .B1(new_n458), .B2(new_n457), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n854), .B(KEYINPUT37), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n448), .A2(new_n846), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n460), .A2(new_n863), .A3(new_n864), .A4(new_n477), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(KEYINPUT38), .B(new_n853), .C1(new_n858), .C2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n460), .A2(new_n863), .A3(new_n477), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n865), .ZN(new_n870));
  INV_X1    g0670(.A(new_n480), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(new_n863), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n706), .B1(KEYINPUT90), .B2(KEYINPUT106), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n702), .A2(new_n663), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n704), .A2(KEYINPUT106), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n702), .B2(new_n663), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n708), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n410), .A2(G169), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT14), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n413), .A3(new_n412), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n392), .B(new_n663), .C1(new_n652), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n392), .A2(new_n663), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n416), .A2(new_n425), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n803), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT40), .B1(new_n875), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n881), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n853), .B1(new_n858), .B2(new_n866), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n873), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n867), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n500), .A2(new_n881), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n672), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT107), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n894), .B2(new_n867), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n867), .A2(new_n874), .A3(new_n903), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT105), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n867), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT104), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n865), .A3(new_n862), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n910), .B2(new_n853), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT39), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n867), .A2(new_n874), .A3(new_n903), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n884), .A2(new_n392), .A3(new_n676), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n906), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n846), .B1(new_n461), .B2(new_n476), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n885), .A2(new_n887), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n650), .A2(new_n676), .A3(new_n804), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n801), .A2(new_n495), .A3(new_n676), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n919), .B1(new_n924), .B2(new_n895), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n918), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n712), .A2(new_n500), .A3(new_n715), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n656), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n845), .B1(new_n902), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n902), .B2(new_n929), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n523), .B(KEYINPUT101), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(KEYINPUT35), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n933), .A2(new_n225), .A3(new_n212), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n935), .A2(KEYINPUT102), .B1(KEYINPUT35), .B2(new_n932), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(KEYINPUT102), .B2(new_n935), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n213), .A2(new_n220), .A3(new_n434), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n223), .B2(G68), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n940), .A2(new_n254), .A3(G13), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n931), .A2(new_n938), .A3(new_n941), .ZN(G367));
  AOI211_X1 g0742(.A(new_n540), .B(new_n535), .C1(new_n539), .C2(new_n663), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n644), .A2(new_n676), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n683), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n622), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n663), .B1(new_n948), .B2(new_n644), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n946), .B2(KEYINPUT42), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n579), .A2(new_n676), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n641), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n577), .B2(new_n952), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n947), .A2(new_n950), .B1(KEYINPUT43), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n680), .A2(new_n945), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n687), .B(KEYINPUT41), .Z(new_n960));
  MUX2_X1   g0760(.A(new_n634), .B(new_n679), .S(new_n682), .Z(new_n961));
  XNOR2_X1  g0761(.A(new_n674), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n716), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT109), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n684), .A2(new_n945), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n684), .A2(new_n945), .ZN(new_n967));
  XOR2_X1   g0767(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n680), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT109), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n962), .A2(new_n972), .A3(new_n716), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n681), .A2(new_n966), .A3(new_n969), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n964), .A2(new_n971), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n960), .B1(new_n975), .B2(new_n716), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n720), .A2(G1), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n959), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n731), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n737), .B1(new_n206), .B2(new_n482), .C1(new_n240), .C2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(new_n722), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n746), .A2(new_n281), .B1(new_n817), .B2(new_n586), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n286), .B(new_n982), .C1(G283), .C2(new_n743), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n753), .A2(G97), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(new_n775), .C2(new_n766), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n755), .A2(G116), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT46), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G311), .A2(new_n757), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n987), .B2(new_n986), .C1(new_n763), .C2(new_n492), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n766), .A2(new_n826), .B1(new_n433), .B2(new_n820), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT110), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n817), .A2(new_n767), .B1(new_n779), .B2(new_n223), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G143), .B2(new_n757), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n763), .A2(new_n218), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n753), .A2(G77), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n439), .B1(new_n745), .B2(G150), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n985), .A2(new_n989), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n981), .B1(new_n726), .B2(new_n954), .C1(new_n1000), .C2(new_n785), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n978), .A2(new_n1001), .ZN(G387));
  NAND2_X1  g0802(.A1(new_n964), .A2(new_n973), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1003), .B(new_n687), .C1(new_n716), .C2(new_n962), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n728), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n1005), .A2(new_n689), .B1(G107), .B2(new_n206), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n237), .A2(new_n261), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n689), .ZN(new_n1008));
  AOI211_X1 g0808(.A(G45), .B(new_n1008), .C1(G68), .C2(G77), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n362), .A2(G50), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT50), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n979), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1006), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n737), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n722), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n757), .A2(G322), .B1(new_n741), .B2(G311), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n281), .B2(new_n779), .C1(new_n775), .C2(new_n746), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n764), .A2(G283), .B1(G294), .B2(new_n755), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT49), .Z(new_n1023));
  AOI21_X1  g0823(.A(new_n286), .B1(new_n823), .B2(G326), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n225), .B2(new_n752), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n823), .A2(G150), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n745), .A2(G50), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n439), .B1(new_n755), .B2(G77), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1026), .A2(new_n984), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n764), .A2(new_n574), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n757), .A2(G159), .B1(new_n741), .B2(new_n363), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n218), .C2(new_n779), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1023), .A2(new_n1025), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1015), .B1(new_n1033), .B2(new_n736), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n679), .A2(new_n725), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n962), .A2(new_n977), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT111), .Z(new_n1038));
  NAND3_X1  g0838(.A1(new_n1004), .A2(new_n1036), .A3(new_n1038), .ZN(G393));
  INV_X1    g0839(.A(KEYINPUT112), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n971), .A2(new_n1040), .A3(new_n974), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n681), .A2(KEYINPUT112), .A3(new_n966), .A4(new_n969), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1003), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(new_n687), .A3(new_n975), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n737), .B1(new_n301), .B2(new_n206), .C1(new_n244), .C2(new_n979), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n722), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT113), .Z(new_n1047));
  OAI22_X1  g0847(.A1(new_n817), .A2(new_n281), .B1(new_n779), .B2(new_n586), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G311), .A2(new_n745), .B1(new_n757), .B2(G317), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(G116), .C2(new_n764), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n286), .B1(new_n755), .B2(G283), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n754), .B(new_n1052), .C1(new_n781), .C2(new_n766), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT114), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n439), .B1(new_n755), .B2(G68), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n779), .B2(new_n362), .C1(new_n223), .C2(new_n817), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n816), .B(new_n1056), .C1(G143), .C2(new_n823), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G150), .A2(new_n757), .B1(new_n745), .B2(G159), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1058), .A2(KEYINPUT51), .B1(new_n763), .B2(new_n220), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(KEYINPUT51), .B2(new_n1058), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1051), .A2(new_n1054), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1047), .B1(new_n1061), .B2(new_n785), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n945), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1062), .B1(new_n1063), .B2(new_n725), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n977), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1044), .A2(new_n1066), .ZN(G390));
  NOR3_X1   g0867(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT105), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1068), .A2(new_n1069), .B1(new_n917), .B2(new_n924), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n867), .A2(new_n874), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n714), .A2(new_n804), .A3(new_n676), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1072), .A2(new_n923), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1071), .B(new_n916), .C1(new_n1073), .C2(new_n921), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n709), .A2(new_n804), .A3(new_n920), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1070), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n672), .B1(new_n880), .B2(new_n708), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1077), .A2(new_n888), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n922), .A2(new_n923), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n917), .B1(new_n1079), .B2(new_n920), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n906), .B2(new_n915), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1074), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1076), .A2(new_n1083), .A3(new_n977), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT115), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1076), .A2(new_n1083), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n500), .A2(new_n1077), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n927), .A2(new_n656), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n920), .B1(new_n709), .B2(new_n804), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1079), .B1(new_n1089), .B2(new_n1078), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1077), .A2(new_n804), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1075), .B(new_n1073), .C1(new_n920), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1088), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1076), .A2(new_n1083), .A3(new_n1093), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n687), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n723), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n722), .B1(new_n363), .B2(new_n811), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n830), .B1(new_n586), .B2(new_n766), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT116), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n439), .B1(new_n820), .B2(new_n563), .C1(new_n817), .C2(new_n492), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n758), .A2(new_n818), .B1(new_n779), .B2(new_n301), .ZN(new_n1103));
  OR3_X1    g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n763), .A2(new_n220), .B1(new_n225), .B2(new_n746), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT117), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT53), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n820), .B2(new_n360), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n755), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n823), .A2(G125), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n439), .B1(new_n741), .B2(G137), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n223), .C2(new_n752), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n745), .A2(G132), .B1(new_n743), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n757), .A2(G128), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(new_n763), .C2(new_n767), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1104), .A2(new_n1106), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1099), .B1(new_n1118), .B2(new_n736), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT118), .Z(new_n1120));
  NAND2_X1  g0920(.A1(new_n1098), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1085), .A2(new_n1097), .A3(new_n1121), .ZN(G378));
  NOR2_X1   g0922(.A1(new_n752), .A2(new_n433), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n574), .B2(new_n743), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n818), .B2(new_n766), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n286), .A2(G41), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n820), .B2(new_n220), .C1(new_n817), .C2(new_n301), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n492), .A2(new_n746), .B1(new_n758), .B2(new_n225), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n1125), .A2(new_n994), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1129), .A2(KEYINPUT58), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(KEYINPUT58), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n764), .A2(G150), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n743), .A2(G137), .B1(new_n755), .B2(new_n1114), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n745), .A2(G128), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n757), .A2(G125), .B1(new_n741), .B2(G132), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n1136), .A2(KEYINPUT59), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(KEYINPUT59), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n283), .B(new_n255), .C1(new_n752), .C2(new_n767), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G124), .B2(new_n823), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(G50), .B(new_n1126), .C1(new_n283), .C2(new_n255), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n1130), .A2(new_n1131), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n722), .B1(G50), .B2(new_n811), .C1(new_n1143), .C2(new_n785), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n368), .A2(new_n846), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT55), .Z(new_n1146));
  NAND2_X1  g0946(.A1(new_n381), .A2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1148));
  AOI21_X1  g0948(.A(new_n379), .B1(new_n371), .B2(new_n373), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1146), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1148), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1146), .B(new_n379), .C1(new_n371), .C2(new_n373), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1144), .B1(new_n1157), .B2(new_n723), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT120), .Z(new_n1159));
  NAND2_X1  g0959(.A1(new_n926), .A2(KEYINPUT121), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1157), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n897), .A2(new_n1161), .A3(G330), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1071), .A2(new_n881), .A3(new_n888), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(KEYINPUT40), .B1(new_n892), .B2(new_n895), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1157), .B1(new_n1164), .B2(new_n672), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1160), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1161), .B1(new_n897), .B2(G330), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n672), .B(new_n1157), .C1(new_n890), .C2(new_n896), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n926), .B(KEYINPUT121), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1159), .B1(new_n1170), .B2(new_n977), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1088), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1096), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n918), .B(new_n925), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n926), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(KEYINPUT57), .A3(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(KEYINPUT122), .B(new_n687), .C1(new_n1173), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1096), .A2(new_n1172), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1170), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n687), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1174), .A2(KEYINPUT57), .A3(new_n1175), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1184), .B2(new_n1178), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(KEYINPUT122), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1171), .B1(new_n1182), .B2(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(new_n1172), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1189), .A2(new_n960), .A3(new_n1093), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT123), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n921), .A2(new_n723), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n722), .B1(G68), .B2(new_n811), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G132), .A2(new_n757), .B1(new_n745), .B2(G137), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n439), .B1(new_n755), .B2(G159), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n817), .C2(new_n1113), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1123), .B(new_n1196), .C1(G128), .C2(new_n823), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n763), .A2(new_n223), .B1(new_n360), .B2(new_n779), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT124), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n439), .B1(new_n820), .B2(new_n301), .C1(new_n817), .C2(new_n225), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G77), .B2(new_n753), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n758), .A2(new_n586), .B1(new_n779), .B2(new_n492), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G283), .B2(new_n745), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n823), .A2(G303), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1030), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1200), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1193), .B1(new_n1207), .B2(new_n736), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1188), .A2(new_n977), .B1(new_n1192), .B2(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1191), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(G381));
  NOR3_X1   g1011(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1212));
  INV_X1    g1012(.A(G390), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1210), .ZN(new_n1214));
  OR4_X1    g1014(.A1(G387), .A2(new_n1214), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1015(.A(new_n1171), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1185), .A2(KEYINPUT122), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1185), .A2(KEYINPUT122), .B1(new_n1180), .B2(new_n1179), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(G378), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n662), .A2(G213), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(G407), .A2(G213), .A3(new_n1223), .ZN(G409));
  NAND2_X1  g1024(.A1(G387), .A2(new_n1213), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(G390), .A2(new_n978), .A3(new_n1001), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(G393), .B(new_n790), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1225), .A2(new_n1228), .A3(new_n1226), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G378), .B(new_n1171), .C1(new_n1182), .C2(new_n1186), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1159), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1174), .A2(new_n977), .A3(new_n1175), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n1179), .C2(new_n960), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1220), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1221), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1222), .A2(G2897), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1090), .A2(new_n1092), .A3(new_n1088), .A4(KEYINPUT60), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1242), .A2(new_n687), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT60), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1093), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1245), .B2(new_n1189), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1209), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(G384), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n837), .A3(new_n843), .A4(new_n1209), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1249), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1241), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT126), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1248), .A2(new_n1250), .A3(new_n1249), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1240), .A3(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT61), .B1(new_n1239), .B2(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1254), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n1239), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1222), .B1(new_n1233), .B2(new_n1237), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(KEYINPUT63), .A3(new_n1254), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1232), .A2(new_n1259), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1263), .A2(new_n1266), .A3(new_n1254), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1268), .B1(new_n1263), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1266), .B1(new_n1263), .B2(new_n1254), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1267), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1265), .B1(new_n1272), .B2(new_n1232), .ZN(G405));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1233), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1254), .B1(new_n1219), .B2(G378), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G375), .A2(new_n1261), .A3(new_n1220), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1232), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1276), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1282), .A2(new_n1278), .A3(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1281), .A2(new_n1284), .ZN(G402));
endmodule


