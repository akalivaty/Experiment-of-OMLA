//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n460), .B1(new_n449), .B2(new_n453), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n467), .A3(G137), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n466), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n478), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .A3(G138), .ZN(new_n486));
  NOR3_X1   g061(.A1(new_n486), .A2(new_n464), .A3(new_n465), .ZN(new_n487));
  AND2_X1   g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n467), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n472), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n492), .B(new_n493), .C1(new_n476), .C2(new_n477), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n489), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT71), .A3(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT5), .B2(new_n504), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n504), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n511), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G89), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n517), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n521), .B(new_n522), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(G168));
  AOI22_X1  g105(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n510), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n508), .A2(G90), .A3(new_n516), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n514), .A2(G52), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n533), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n532), .B(new_n540), .C1(new_n536), .C2(new_n537), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n510), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n514), .A2(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n517), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  AND2_X1   g130(.A1(new_n508), .A2(new_n516), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n516), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n514), .A2(new_n560), .A3(G53), .ZN(new_n561));
  AOI22_X1  g136(.A1(G91), .A2(new_n556), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(new_n510), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  INV_X1    g143(.A(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT77), .B1(new_n517), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n508), .A2(new_n571), .A3(G87), .A4(new_n516), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n508), .A2(G74), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G49), .B2(new_n514), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n514), .A2(G48), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n505), .A2(new_n507), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n578), .B1(new_n584), .B2(G651), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n508), .A2(G86), .A3(new_n516), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n556), .A2(KEYINPUT78), .A3(G86), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n556), .A2(G85), .B1(G47), .B2(new_n514), .ZN(new_n591));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n582), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(new_n556), .A2(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT79), .B(G66), .Z(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n582), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g181(.A(new_n605), .B1(G868), .B2(G171), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G280));
  INV_X1    g186(.A(G860), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n604), .B1(G559), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT80), .ZN(G148));
  OR2_X1    g189(.A1(new_n604), .A2(G559), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n472), .A2(G2104), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n478), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(G2100), .ZN(new_n626));
  AOI22_X1  g201(.A1(G123), .A2(new_n479), .B1(new_n482), .B2(G135), .ZN(new_n627));
  OAI221_X1 g202(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT83), .B(G2096), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n625), .A2(G2100), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n626), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT84), .ZN(G156));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n638), .B(new_n644), .Z(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT86), .Z(new_n656));
  INV_X1    g231(.A(new_n654), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n651), .A2(new_n652), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2096), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g248(.A(new_n673), .B(new_n672), .S(new_n665), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT87), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT96), .B(KEYINPUT24), .Z(new_n685));
  INV_X1    g260(.A(G34), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n686), .B2(new_n685), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT97), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G160), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n684), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G2084), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(G162), .A2(G29), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G29), .B2(G35), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT29), .B(G2090), .Z(new_n697));
  OAI21_X1  g272(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT30), .B(G28), .ZN(new_n700));
  OR2_X1    g275(.A1(KEYINPUT31), .A2(G11), .ZN(new_n701));
  NAND2_X1  g276(.A1(KEYINPUT31), .A2(G11), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n700), .A2(new_n684), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n699), .B(new_n703), .C1(new_n684), .C2(new_n629), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n684), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n479), .A2(G129), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n482), .A2(G141), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n705), .B1(new_n713), .B2(new_n684), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n714), .B(new_n715), .Z(new_n716));
  NOR3_X1   g291(.A1(new_n698), .A2(new_n704), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n684), .A2(G33), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n482), .A2(G139), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT25), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n719), .B1(new_n466), .B2(new_n720), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI211_X1 g305(.A(G2072), .B(new_n718), .C1(new_n730), .C2(new_n684), .ZN(new_n731));
  INV_X1    g306(.A(G2072), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n684), .B1(new_n727), .B2(new_n728), .ZN(new_n733));
  INV_X1    g308(.A(new_n718), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n690), .B(G2084), .C1(new_n684), .C2(new_n691), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT98), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n684), .A2(G27), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT100), .Z(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n501), .B2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G2078), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n717), .A2(new_n736), .A3(new_n738), .A4(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G168), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G1966), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(G1966), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n604), .A2(G16), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n746), .A2(G4), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(G1348), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G1348), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n755), .B(new_n752), .C1(new_n604), .C2(G16), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n749), .B(new_n750), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n684), .A2(G26), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  AOI22_X1  g334(.A1(G128), .A2(new_n479), .B1(new_n482), .B2(G140), .ZN(new_n760));
  OAI221_X1 g335(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(KEYINPUT94), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(KEYINPUT94), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n759), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n746), .A2(G19), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT93), .Z(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n548), .B2(new_n746), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1341), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n746), .A2(G20), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT23), .Z(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G299), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1956), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n768), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n745), .A2(new_n757), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n746), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n746), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G1961), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT99), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n780), .A2(G1961), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n778), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(G303), .A2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G22), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(G16), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G1971), .ZN(new_n788));
  INV_X1    g363(.A(G1971), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n785), .B(new_n789), .C1(G16), .C2(new_n786), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT32), .B(G1981), .Z(new_n791));
  AND2_X1   g366(.A1(new_n746), .A2(G6), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G305), .B2(G16), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n788), .B(new_n790), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n746), .A2(G23), .ZN(new_n795));
  INV_X1    g370(.A(G288), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n746), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT33), .B(G1976), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n798), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n795), .B(new_n800), .C1(new_n796), .C2(new_n746), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n793), .A2(new_n791), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n794), .A2(KEYINPUT34), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT89), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n482), .A2(G131), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n466), .A2(G107), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n810), .A2(new_n812), .B1(new_n479), .B2(G119), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n806), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n809), .A2(new_n806), .A3(new_n813), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G29), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n684), .A2(G25), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT90), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n823), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n818), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  MUX2_X1   g402(.A(G24), .B(G290), .S(G16), .Z(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(G1986), .Z(new_n829));
  NAND4_X1  g404(.A1(new_n804), .A2(new_n805), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n829), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n794), .A2(KEYINPUT34), .A3(new_n803), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT91), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(KEYINPUT34), .B1(new_n794), .B2(new_n803), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n830), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n836));
  NOR2_X1   g411(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n784), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n830), .A2(new_n833), .A3(new_n836), .A4(new_n834), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT101), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n835), .A2(new_n838), .ZN(new_n842));
  INV_X1    g417(.A(new_n784), .ZN(new_n843));
  AND4_X1   g418(.A1(KEYINPUT101), .A2(new_n842), .A3(new_n843), .A4(new_n840), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(G311));
  AOI21_X1  g420(.A(KEYINPUT102), .B1(new_n839), .B2(new_n840), .ZN(new_n846));
  AND4_X1   g421(.A1(KEYINPUT102), .A2(new_n842), .A3(new_n843), .A4(new_n840), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(G150));
  INV_X1    g423(.A(new_n604), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  INV_X1    g426(.A(new_n548), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n514), .A2(G55), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT103), .B(G93), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n517), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n508), .A2(G67), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n510), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n548), .A2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n851), .B(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n612), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n859), .A2(new_n612), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n872));
  INV_X1    g447(.A(new_n816), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(new_n814), .ZN(new_n874));
  AOI22_X1  g449(.A1(G130), .A2(new_n479), .B1(new_n482), .B2(G142), .ZN(new_n875));
  OAI221_X1 g450(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n622), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(new_n878), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n882), .A3(new_n880), .ZN(new_n885));
  XNOR2_X1  g460(.A(G164), .B(new_n762), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n729), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n729), .A2(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n713), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n713), .B1(new_n887), .B2(new_n888), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n884), .B(new_n885), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n691), .B(new_n629), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(G162), .Z(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT106), .B1(new_n890), .B2(new_n891), .ZN(new_n897));
  INV_X1    g472(.A(new_n891), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n889), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n884), .A2(new_n885), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n897), .A2(new_n900), .A3(KEYINPUT107), .A4(new_n901), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n896), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n901), .A2(new_n889), .A3(new_n898), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n892), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n909), .B2(new_n894), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n872), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n910), .ZN(new_n912));
  INV_X1    g487(.A(new_n872), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n912), .A2(new_n906), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n911), .A2(new_n914), .ZN(G395));
  NAND2_X1  g490(.A1(new_n860), .A2(new_n608), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n917));
  XNOR2_X1  g492(.A(G290), .B(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n796), .ZN(new_n919));
  XNOR2_X1  g494(.A(G303), .B(G305), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n918), .B(G288), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n921), .A3(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT42), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n615), .B(new_n863), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n604), .B(G299), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g506(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(KEYINPUT41), .B2(new_n930), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n931), .B1(new_n935), .B2(new_n929), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n928), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n916), .B1(new_n937), .B2(new_n608), .ZN(G295));
  OAI21_X1  g513(.A(new_n916), .B1(new_n937), .B2(new_n608), .ZN(G331));
  XNOR2_X1  g514(.A(G171), .B(G286), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n864), .ZN(new_n941));
  XNOR2_X1  g516(.A(G171), .B(G168), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n863), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n935), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n924), .A2(new_n926), .ZN(new_n946));
  INV_X1    g521(.A(new_n930), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G37), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n946), .B1(new_n945), .B2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT41), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n930), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n930), .B2(new_n932), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n941), .B2(new_n943), .ZN(new_n957));
  INV_X1    g532(.A(new_n948), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n927), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n950), .A4(new_n949), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n953), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n951), .B2(new_n952), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n959), .A2(KEYINPUT43), .A3(new_n950), .A4(new_n949), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  MUX2_X1   g540(.A(new_n962), .B(new_n965), .S(KEYINPUT44), .Z(G397));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n501), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT50), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n466), .A2(new_n467), .A3(G138), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n499), .B1(new_n970), .B2(new_n490), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n971), .B2(new_n489), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n470), .A2(new_n474), .A3(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n969), .A2(new_n974), .A3(new_n693), .A4(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT118), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1966), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n976), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n982), .B(G1384), .C1(new_n971), .C2(new_n489), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n468), .A2(new_n469), .ZN(new_n985));
  INV_X1    g560(.A(new_n466), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n471), .A2(new_n473), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(G40), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n990), .A2(KEYINPUT118), .A3(new_n693), .A4(new_n974), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n979), .A2(new_n984), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT115), .B(G8), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(G168), .A2(new_n993), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(KEYINPUT51), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n992), .A2(G286), .A3(new_n994), .ZN(new_n999));
  XOR2_X1   g574(.A(KEYINPUT121), .B(KEYINPUT51), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n992), .B2(G8), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT62), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n998), .B(KEYINPUT62), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n989), .B1(new_n968), .B2(new_n982), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n972), .A2(KEYINPUT45), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1971), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n976), .B1(new_n972), .B2(new_n973), .ZN(new_n1011));
  AOI211_X1 g586(.A(KEYINPUT50), .B(G1384), .C1(new_n971), .C2(new_n489), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1011), .A2(G2090), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1007), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n789), .B1(new_n981), .B2(new_n983), .ZN(new_n1015));
  INV_X1    g590(.A(G2090), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n969), .A2(new_n974), .A3(new_n1016), .A4(new_n976), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(KEYINPUT117), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n994), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1020), .B1(G166), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT55), .B(G8), .C1(new_n511), .C2(new_n519), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  AOI221_X4 g601(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n993), .B1(new_n976), .B2(new_n972), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n573), .A2(new_n575), .A3(G1976), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT52), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G288), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n585), .A2(new_n1036), .A3(new_n588), .A4(new_n589), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n577), .B(new_n586), .C1(new_n1038), .C2(new_n510), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G1981), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT116), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n1028), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1042), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1031), .B(new_n1035), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1027), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1008), .A2(new_n742), .A3(new_n1009), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n969), .A2(new_n976), .A3(new_n974), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1048), .A2(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1049), .A2(G2078), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1008), .A2(new_n1009), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  AND4_X1   g630(.A1(G171), .A2(new_n1026), .A3(new_n1047), .A4(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1005), .A2(new_n1006), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1037), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G288), .A2(G1976), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1028), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(G8), .A3(new_n1024), .ZN(new_n1064));
  OAI22_X1  g639(.A1(new_n1061), .A2(new_n1062), .B1(new_n1064), .B2(new_n1046), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n992), .A2(G168), .A3(new_n994), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1026), .A2(new_n1047), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT63), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1063), .A2(G8), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1068), .B1(new_n1070), .B2(new_n1025), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1047), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1065), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n562), .A2(new_n564), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n561), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n560), .B1(new_n514), .B2(G53), .ZN(new_n1077));
  INV_X1    g652(.A(G91), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1076), .A2(new_n1077), .B1(new_n1078), .B2(new_n517), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n563), .A2(new_n510), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1956), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1008), .A2(new_n1009), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1082), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1050), .A2(new_n755), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n976), .A2(new_n972), .A3(new_n767), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n604), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1082), .A2(new_n1086), .A3(new_n1084), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1087), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1082), .A2(new_n1086), .A3(new_n1084), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1087), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1086), .A2(new_n1084), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1082), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(KEYINPUT61), .A3(new_n1091), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n968), .A2(new_n982), .ZN(new_n1100));
  INV_X1    g675(.A(G1996), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1100), .A2(new_n1009), .A3(new_n1101), .A4(new_n976), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n968), .B2(new_n989), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n852), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT120), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1095), .A2(new_n1099), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n1089), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n849), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n604), .A4(new_n1089), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1092), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1000), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n991), .A2(new_n984), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n993), .B1(new_n1118), .B2(new_n979), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1119), .B2(G286), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1002), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1120), .A2(new_n1121), .B1(new_n995), .B2(new_n997), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  NAND2_X1  g698(.A1(G171), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n539), .A2(KEYINPUT54), .A3(new_n541), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1055), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n474), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n471), .A2(KEYINPUT122), .A3(new_n473), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1129), .A2(G40), .A3(new_n987), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT112), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT45), .B1(new_n968), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n972), .A2(KEYINPUT112), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1133), .A2(new_n1137), .A3(new_n1009), .A4(new_n1053), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1052), .A2(new_n1138), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1127), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n993), .B1(new_n1063), .B2(new_n1007), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1024), .B1(new_n1141), .B2(new_n1018), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1059), .A2(new_n1064), .A3(new_n1031), .A4(new_n1035), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1116), .A2(new_n1122), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1057), .A2(new_n1073), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT113), .B1(new_n1137), .B2(new_n989), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT113), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1135), .A2(new_n1148), .A3(new_n976), .A4(new_n1136), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n762), .B(new_n767), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT114), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n713), .B(G1996), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n874), .A2(new_n822), .ZN(new_n1157));
  INV_X1    g732(.A(new_n822), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n817), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(G290), .B(G1986), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1151), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1146), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n762), .A2(G2067), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1157), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1156), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n1150), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n1168));
  NOR2_X1   g743(.A1(G290), .A2(G1986), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1151), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1169), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT125), .B1(new_n1150), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT48), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1173), .A2(new_n1174), .B1(new_n1160), .B2(new_n1151), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1170), .A2(KEYINPUT48), .A3(new_n1172), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1167), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT47), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT46), .B1(new_n1150), .B2(G1996), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT46), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1147), .A2(new_n1149), .A3(new_n1180), .A4(new_n1101), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n713), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1151), .B1(new_n1183), .B2(new_n1153), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1182), .A2(KEYINPUT124), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT124), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1178), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1191), .A2(KEYINPUT47), .A3(new_n1185), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1177), .A2(new_n1188), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1163), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1163), .A2(new_n1193), .A3(KEYINPUT126), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g773(.A1(G227), .A2(new_n462), .ZN(new_n1200));
  XOR2_X1   g774(.A(new_n1200), .B(KEYINPUT127), .Z(new_n1201));
  INV_X1    g775(.A(G401), .ZN(new_n1202));
  AND3_X1   g776(.A1(new_n1201), .A2(new_n682), .A3(new_n1202), .ZN(new_n1203));
  OAI211_X1 g777(.A(new_n962), .B(new_n1203), .C1(new_n906), .C2(new_n912), .ZN(G225));
  INV_X1    g778(.A(G225), .ZN(G308));
endmodule


