//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n530, new_n532, new_n533, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n553, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1154,
    new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n468), .B(KEYINPUT64), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n467), .ZN(new_n473));
  OAI22_X1  g048(.A1(new_n469), .A2(new_n470), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n463), .A2(new_n467), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT65), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT66), .Z(new_n481));
  NOR2_X1   g056(.A1(new_n463), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n478), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT67), .Z(G162));
  OR2_X1    g060(.A1(new_n467), .A2(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n476), .A2(G126), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n467), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n472), .A2(new_n492), .A3(G138), .A4(new_n467), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G543), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT6), .B(G651), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(G543), .ZN(new_n500));
  AOI22_X1  g075(.A1(G88), .A2(new_n499), .B1(new_n500), .B2(G50), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n501), .B1(new_n504), .B2(KEYINPUT68), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n504), .A2(KEYINPUT68), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(G166));
  NAND2_X1  g082(.A1(new_n497), .A2(new_n498), .ZN(new_n508));
  INV_X1    g083(.A(G89), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n498), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G51), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n497), .A2(G63), .A3(G651), .ZN(new_n513));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT7), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n512), .A2(new_n518), .ZN(G168));
  AOI22_X1  g094(.A1(G90), .A2(new_n499), .B1(new_n500), .B2(G52), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n497), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(new_n503), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(G171));
  NAND2_X1  g098(.A1(new_n499), .A2(G81), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n500), .A2(G43), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n497), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n524), .B(new_n525), .C1(new_n503), .C2(new_n526), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT69), .Z(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G860), .ZN(G153));
  AND3_X1   g104(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G36), .ZN(G176));
  NAND2_X1  g106(.A1(G1), .A2(G3), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT8), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(G188));
  NAND2_X1  g109(.A1(G78), .A2(G543), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT71), .ZN(new_n536));
  INV_X1    g111(.A(G65), .ZN(new_n537));
  INV_X1    g112(.A(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT5), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n536), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n503), .B1(new_n543), .B2(KEYINPUT72), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n544), .B1(KEYINPUT72), .B2(new_n543), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT70), .B(KEYINPUT9), .Z(new_n546));
  NAND3_X1  g121(.A1(new_n500), .A2(G53), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n499), .A2(G91), .ZN(new_n548));
  NOR2_X1   g123(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n549));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n510), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n545), .A2(new_n547), .A3(new_n548), .A4(new_n551), .ZN(G299));
  XNOR2_X1  g127(.A(G171), .B(KEYINPUT73), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(G301));
  INV_X1    g129(.A(G168), .ZN(G286));
  INV_X1    g130(.A(G166), .ZN(G303));
  OAI21_X1  g131(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT74), .ZN(new_n558));
  AOI22_X1  g133(.A1(G87), .A2(new_n499), .B1(new_n500), .B2(G49), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(G288));
  NAND3_X1  g135(.A1(new_n539), .A2(new_n541), .A3(G61), .ZN(new_n561));
  NAND2_X1  g136(.A1(G73), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n565), .A2(new_n567), .A3(G48), .A4(G543), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n563), .A2(G651), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n498), .A2(KEYINPUT76), .A3(G48), .A4(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n497), .A2(new_n498), .A3(G86), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT75), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n497), .A2(new_n498), .A3(new_n573), .A4(G86), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n569), .A2(new_n570), .A3(new_n572), .A4(new_n574), .ZN(G305));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  INV_X1    g151(.A(G47), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n508), .A2(new_n576), .B1(new_n510), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n503), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n499), .A2(KEYINPUT10), .A3(G92), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  INV_X1    g160(.A(G92), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n508), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n584), .A2(new_n587), .B1(G54), .B2(new_n500), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n542), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n503), .B1(new_n591), .B2(KEYINPUT77), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(KEYINPUT77), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT78), .Z(new_n595));
  OAI21_X1  g170(.A(new_n583), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n583), .B1(new_n595), .B2(G868), .ZN(G321));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  XOR2_X1   g173(.A(G299), .B(KEYINPUT79), .Z(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  INV_X1    g178(.A(new_n595), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G559), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n528), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g184(.A(KEYINPUT64), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n468), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(new_n472), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n476), .A2(G123), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n482), .A2(G135), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(G156));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT80), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2430), .Z(new_n628));
  AOI21_X1  g203(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n627), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT16), .B(G1341), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(G14), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n630), .B2(new_n636), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(KEYINPUT17), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n640), .A2(new_n641), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n642), .A2(KEYINPUT17), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n647), .C1(new_n648), .C2(new_n644), .ZN(new_n649));
  OR3_X1    g224(.A1(new_n647), .A2(KEYINPUT18), .A3(new_n643), .ZN(new_n650));
  OAI21_X1  g225(.A(KEYINPUT18), .B1(new_n647), .B2(new_n643), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2096), .B(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n657), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(KEYINPUT81), .B1(new_n658), .B2(new_n659), .ZN(new_n666));
  OR3_X1    g241(.A1(new_n665), .A2(new_n657), .A3(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n661), .B(new_n663), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n668), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1991), .ZN(new_n671));
  INV_X1    g246(.A(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  AOI22_X1  g252(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n678), .A2(new_n467), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT25), .ZN(new_n681));
  INV_X1    g256(.A(G103), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n468), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g258(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n684));
  AOI22_X1  g259(.A1(new_n482), .A2(G139), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G29), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G29), .B2(G33), .ZN(new_n688));
  INV_X1    g263(.A(G2072), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT90), .Z(new_n691));
  AOI22_X1  g266(.A1(G105), .A2(new_n611), .B1(new_n476), .B2(G129), .ZN(new_n692));
  NAND3_X1  g267(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT26), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G141), .B2(new_n482), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G29), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G29), .B2(G32), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT27), .B(G1996), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  AND2_X1   g276(.A1(KEYINPUT24), .A2(G34), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(KEYINPUT24), .B2(G34), .ZN(new_n703));
  OAI22_X1  g278(.A1(G160), .A2(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n699), .A2(new_n700), .B1(G2084), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n688), .B2(new_n689), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n691), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT91), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n701), .A2(G35), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT95), .Z(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G162), .B2(new_n701), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT29), .ZN(new_n712));
  INV_X1    g287(.A(G2090), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n701), .A2(G26), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n476), .A2(G128), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n482), .A2(G140), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n467), .A2(G116), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n715), .B1(new_n720), .B2(G29), .ZN(new_n721));
  MUX2_X1   g296(.A(new_n715), .B(new_n721), .S(KEYINPUT28), .Z(new_n722));
  INV_X1    g297(.A(G2067), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G21), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G168), .B2(new_n725), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1966), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT31), .B(G11), .Z(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT92), .B(KEYINPUT30), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(G28), .ZN(new_n731));
  AOI21_X1  g306(.A(G29), .B1(new_n730), .B2(G28), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G164), .A2(new_n701), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G27), .B2(new_n701), .ZN(new_n735));
  INV_X1    g310(.A(G2078), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n733), .B1(new_n701), .B2(new_n621), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n728), .B(new_n737), .C1(new_n736), .C2(new_n735), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n725), .A2(G5), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G171), .B2(new_n725), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT93), .ZN(new_n741));
  INV_X1    g316(.A(new_n722), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n741), .A2(G1961), .B1(G2067), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G16), .A2(G19), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n528), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT88), .B(G1341), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  AND4_X1   g322(.A1(new_n724), .A2(new_n738), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT23), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G299), .B2(G16), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n725), .A2(G20), .ZN(new_n751));
  MUX2_X1   g326(.A(new_n749), .B(new_n750), .S(new_n751), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1956), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n714), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n704), .A2(G2084), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n755), .B1(new_n699), .B2(new_n700), .C1(new_n741), .C2(G1961), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT94), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n725), .A2(G4), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n595), .B2(new_n725), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1348), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n708), .A2(new_n754), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G6), .B(G305), .S(G16), .Z(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT84), .Z(new_n763));
  XOR2_X1   g338(.A(KEYINPUT32), .B(G1981), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT85), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G166), .A2(new_n725), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n725), .B2(G22), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(G1971), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G23), .ZN(new_n771));
  INV_X1    g346(.A(G288), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G16), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT33), .B(G1976), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n769), .B2(G1971), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n763), .A2(new_n765), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n766), .A2(new_n770), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT83), .B(KEYINPUT34), .Z(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n701), .A2(G25), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n476), .A2(G119), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n482), .A2(G131), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n467), .A2(G107), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT82), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n782), .B1(new_n789), .B2(new_n701), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT35), .B(G1991), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n725), .A2(G24), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n581), .B2(new_n725), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1986), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n780), .A2(new_n781), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n799));
  MUX2_X1   g374(.A(new_n799), .B(KEYINPUT36), .S(KEYINPUT87), .Z(new_n800));
  OR2_X1    g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n799), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n761), .A2(new_n801), .A3(new_n802), .ZN(G150));
  INV_X1    g378(.A(G150), .ZN(G311));
  NAND2_X1  g379(.A1(G80), .A2(G543), .ZN(new_n805));
  INV_X1    g380(.A(G67), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n542), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G651), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT96), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT98), .B(G93), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT97), .B(G55), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n499), .A2(new_n810), .B1(new_n500), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT37), .Z(new_n815));
  INV_X1    g390(.A(G860), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n595), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n817), .B(new_n818), .Z(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n528), .A2(new_n813), .ZN(new_n821));
  INV_X1    g396(.A(new_n813), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(new_n527), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(KEYINPUT99), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n528), .A2(new_n813), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n826), .A2(new_n827), .A3(new_n823), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n816), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n819), .B1(new_n825), .B2(new_n828), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n815), .B1(new_n830), .B2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(G162), .B(KEYINPUT100), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G160), .ZN(new_n834));
  INV_X1    g409(.A(new_n621), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G160), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n833), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n621), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n696), .B(new_n720), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n489), .A2(new_n842), .A3(new_n494), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n489), .B2(new_n494), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n841), .B(new_n845), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n686), .ZN(new_n847));
  INV_X1    g422(.A(G142), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n467), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n473), .A2(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n476), .A2(G130), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(KEYINPUT102), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(KEYINPUT102), .B2(new_n852), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n613), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n788), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n847), .B(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n840), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n847), .B(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n836), .A2(new_n839), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n858), .A2(KEYINPUT104), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT104), .B1(new_n858), .B2(new_n862), .ZN(new_n864));
  OR3_X1    g439(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT40), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT40), .B1(new_n863), .B2(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(G395));
  XOR2_X1   g442(.A(G299), .B(new_n594), .Z(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n829), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n605), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n829), .B(KEYINPUT105), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n606), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n869), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(KEYINPUT41), .B2(new_n869), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n872), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G288), .B(G305), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G166), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n581), .B(KEYINPUT107), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT42), .Z(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n876), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT108), .ZN(new_n888));
  INV_X1    g463(.A(new_n880), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n889), .B2(new_n875), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT109), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n876), .A2(new_n893), .A3(new_n880), .A4(new_n886), .ZN(new_n894));
  OAI211_X1 g469(.A(KEYINPUT109), .B(new_n885), .C1(new_n889), .C2(new_n875), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n888), .A2(new_n892), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(G868), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n822), .A2(G868), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(G295));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n898), .ZN(G331));
  NAND2_X1  g475(.A1(G171), .A2(G286), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n553), .B2(G286), .ZN(new_n902));
  INV_X1    g477(.A(new_n828), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n827), .B1(new_n826), .B2(new_n823), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n902), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n825), .A2(new_n828), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT110), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n829), .A2(KEYINPUT110), .A3(new_n902), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n869), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n905), .A2(new_n907), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n879), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n911), .B2(new_n912), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n917), .B2(new_n884), .ZN(new_n918));
  INV_X1    g493(.A(new_n884), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n913), .B2(new_n916), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT43), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n911), .A2(new_n912), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n911), .A2(new_n912), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n922), .A2(new_n884), .A3(new_n923), .A4(new_n915), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n868), .A2(KEYINPUT41), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n868), .B2(new_n877), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n909), .A2(new_n910), .A3(new_n927), .ZN(new_n928));
  OAI22_X1  g503(.A1(new_n928), .A2(KEYINPUT112), .B1(new_n869), .B2(new_n914), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n928), .A2(KEYINPUT112), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n919), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND4_X1   g506(.A1(KEYINPUT43), .A2(new_n924), .A3(new_n925), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT44), .B1(new_n921), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n918), .B2(new_n920), .ZN(new_n936));
  AND4_X1   g511(.A1(new_n935), .A2(new_n924), .A3(new_n925), .A4(new_n931), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(new_n938), .ZN(G397));
  INV_X1    g514(.A(G1384), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n845), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI22_X1  g518(.A1(G101), .A2(new_n611), .B1(new_n482), .B2(G137), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n465), .A2(G2105), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(G40), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n696), .B(new_n672), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n720), .B(new_n723), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT113), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n788), .A2(new_n791), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n788), .A2(new_n791), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n581), .B(G1986), .Z(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n947), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G40), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n466), .A2(new_n474), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n489), .B2(new_n494), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1976), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n962), .B(G8), .C1(new_n963), .C2(G288), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n772), .B2(G1976), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(KEYINPUT52), .B2(new_n964), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(G8), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT115), .B1(G305), .B2(G1981), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n568), .A2(new_n564), .ZN(new_n972));
  INV_X1    g547(.A(new_n562), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n497), .B2(G61), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n972), .B(new_n570), .C1(new_n974), .C2(new_n503), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n572), .A2(new_n574), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n978));
  INV_X1    g553(.A(G1981), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n976), .A2(new_n977), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n971), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n571), .ZN(new_n982));
  OAI21_X1  g557(.A(G1981), .B1(new_n975), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT116), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n985), .B(G1981), .C1(new_n975), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n970), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n971), .A2(new_n980), .B1(new_n984), .B2(new_n986), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT117), .B1(new_n991), .B2(KEYINPUT49), .ZN(new_n992));
  AND4_X1   g567(.A1(KEYINPUT117), .A2(new_n981), .A3(KEYINPUT49), .A4(new_n987), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT118), .B(new_n990), .C1(new_n992), .C2(new_n993), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n969), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(G166), .B2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT55), .B(G8), .C1(new_n505), .C2(new_n506), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT45), .B(new_n940), .C1(new_n843), .C2(new_n844), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n495), .A2(new_n940), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n946), .B1(new_n1006), .B2(new_n942), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1971), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(KEYINPUT50), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n961), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1009), .A2(new_n713), .A3(new_n1011), .A4(new_n960), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1004), .B(G8), .C1(new_n1008), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1012), .B1(new_n1017), .B2(G1971), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(KEYINPUT114), .A3(G8), .A4(new_n1004), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT119), .B(new_n1012), .C1(new_n1017), .C2(G1971), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n1013), .B2(new_n1008), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1023), .A3(G8), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1004), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1020), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n999), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT56), .B(G2072), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1017), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1009), .A2(new_n960), .A3(new_n1011), .ZN(new_n1031));
  INV_X1    g606(.A(G1956), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G299), .B(KEYINPUT57), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1035), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1038));
  INV_X1    g613(.A(G1348), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(G2067), .B2(new_n962), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(new_n595), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1036), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1038), .A2(new_n1036), .A3(KEYINPUT61), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1041), .A2(new_n595), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT60), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1051));
  INV_X1    g626(.A(new_n962), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT124), .B(KEYINPUT58), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(G1341), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1051), .A2(G1996), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1055), .A2(new_n528), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1056), .A2(KEYINPUT59), .ZN(new_n1057));
  OR3_X1    g632(.A1(new_n1041), .A2(new_n604), .A3(KEYINPUT60), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(KEYINPUT59), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1050), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1036), .B(new_n1043), .C1(new_n1048), .C2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(new_n1051), .B2(G2078), .ZN(new_n1063));
  INV_X1    g638(.A(G1961), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1031), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1007), .B1(new_n942), .B2(new_n1006), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n736), .A2(KEYINPUT53), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1063), .B(new_n1065), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n553), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n467), .B1(new_n465), .B2(KEYINPUT125), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(KEYINPUT125), .B2(new_n465), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n474), .A2(new_n959), .A3(new_n1067), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n943), .A2(new_n1005), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1069), .B1(new_n553), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1074), .B2(G171), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1068), .A2(new_n553), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1075), .A2(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n1080));
  INV_X1    g655(.A(G1966), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n960), .B1(KEYINPUT45), .B2(new_n961), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1006), .A2(new_n942), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT120), .B(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1009), .A2(new_n1085), .A3(new_n1011), .A4(new_n960), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT120), .B1(new_n1066), .B2(new_n1081), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1080), .B(G8), .C1(new_n1089), .C2(G286), .ZN(new_n1090));
  OAI21_X1  g665(.A(G8), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(KEYINPUT51), .C1(new_n1001), .C2(G168), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(G8), .A3(G286), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1061), .A2(new_n1079), .A3(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1094), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1096), .A2(new_n1101), .A3(new_n1069), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1028), .B1(new_n1095), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n996), .A2(new_n997), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G288), .A2(G1976), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1104), .A2(new_n1105), .B1(new_n971), .B2(new_n980), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1106), .A2(new_n970), .B1(new_n999), .B2(new_n1020), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1018), .A2(G8), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1020), .B(KEYINPUT63), .C1(new_n1004), .C2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(G8), .B(G168), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n997), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n981), .A2(new_n987), .A3(KEYINPUT49), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n991), .A2(KEYINPUT117), .A3(KEYINPUT49), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT118), .B1(new_n1117), .B2(new_n990), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n968), .B(new_n1111), .C1(new_n1112), .C2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1109), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1119), .B2(new_n1027), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1016), .A2(new_n1019), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n998), .A2(new_n1124), .A3(KEYINPUT121), .A4(new_n1111), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1122), .A2(new_n1125), .A3(KEYINPUT122), .A4(new_n1123), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1107), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1103), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g707(.A(KEYINPUT123), .B(new_n1107), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n958), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n947), .A2(new_n672), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT46), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n949), .A2(new_n697), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1135), .A2(new_n1136), .B1(new_n947), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1136), .B2(new_n1135), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT47), .ZN(new_n1140));
  NOR4_X1   g715(.A1(new_n943), .A2(G1986), .A3(G290), .A4(new_n946), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT48), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n956), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n952), .A2(new_n954), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(G2067), .B2(new_n720), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(KEYINPUT127), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1146), .A2(new_n946), .A3(new_n943), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(KEYINPUT127), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1143), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1134), .A2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g725(.A1(new_n654), .A2(G319), .ZN(new_n1152));
  NOR3_X1   g726(.A1(G229), .A2(G401), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g727(.A(new_n1153), .B1(new_n863), .B2(new_n864), .ZN(new_n1154));
  NOR2_X1   g728(.A1(new_n936), .A2(new_n937), .ZN(new_n1155));
  NOR2_X1   g729(.A1(new_n1154), .A2(new_n1155), .ZN(G308));
  OAI221_X1 g730(.A(new_n1153), .B1(new_n863), .B2(new_n864), .C1(new_n936), .C2(new_n937), .ZN(G225));
endmodule


