

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720;

  NOR2_X1 U365 ( .A1(n677), .A2(n696), .ZN(n678) );
  AND2_X1 U366 ( .A1(n371), .A2(n369), .ZN(n571) );
  AND2_X1 U367 ( .A1(n403), .A2(n344), .ZN(n401) );
  OR2_X1 U368 ( .A1(n653), .A2(n404), .ZN(n403) );
  XNOR2_X1 U369 ( .A(n418), .B(n467), .ZN(n691) );
  INV_X1 U370 ( .A(G137), .ZN(n426) );
  XNOR2_X1 U371 ( .A(n419), .B(n706), .ZN(n418) );
  NOR2_X1 U372 ( .A1(n596), .A2(n696), .ZN(n598) );
  XNOR2_X2 U373 ( .A(n450), .B(n449), .ZN(n705) );
  XNOR2_X2 U374 ( .A(n513), .B(n442), .ZN(n450) );
  INV_X1 U375 ( .A(n376), .ZN(n573) );
  INV_X1 U376 ( .A(n479), .ZN(n586) );
  NOR2_X1 U377 ( .A1(n688), .A2(n696), .ZN(n690) );
  NOR2_X1 U378 ( .A1(n590), .A2(n696), .ZN(n592) );
  XNOR2_X1 U379 ( .A(n395), .B(n430), .ZN(n349) );
  OR2_X2 U380 ( .A1(n626), .A2(n627), .ZN(n634) );
  NOR2_X1 U381 ( .A1(n691), .A2(G902), .ZN(n472) );
  XNOR2_X1 U382 ( .A(n365), .B(KEYINPUT78), .ZN(n364) );
  XNOR2_X1 U383 ( .A(n413), .B(KEYINPUT65), .ZN(n537) );
  XNOR2_X1 U384 ( .A(n423), .B(KEYINPUT104), .ZN(n719) );
  NAND2_X1 U385 ( .A1(n414), .A2(n630), .ZN(n413) );
  NAND2_X1 U386 ( .A1(n401), .A2(n400), .ZN(n528) );
  NAND2_X1 U387 ( .A1(n349), .A2(n389), .ZN(n529) );
  AND2_X1 U388 ( .A1(n549), .A2(n548), .ZN(n568) );
  NOR2_X1 U389 ( .A1(n523), .A2(n376), .ZN(n524) );
  XNOR2_X1 U390 ( .A(n433), .B(n411), .ZN(n633) );
  XNOR2_X1 U391 ( .A(n472), .B(n471), .ZN(n626) );
  XNOR2_X1 U392 ( .A(n426), .B(G140), .ZN(n459) );
  INV_X2 U393 ( .A(G143), .ZN(n392) );
  XNOR2_X1 U394 ( .A(n466), .B(KEYINPUT10), .ZN(n706) );
  INV_X1 U395 ( .A(G134), .ZN(n441) );
  NAND2_X1 U396 ( .A1(n366), .A2(n362), .ZN(n580) );
  NOR2_X1 U397 ( .A1(n364), .A2(n363), .ZN(n362) );
  XNOR2_X1 U398 ( .A(n368), .B(n367), .ZN(n366) );
  NAND2_X1 U399 ( .A1(n621), .A2(n563), .ZN(n363) );
  XOR2_X1 U400 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n500) );
  XNOR2_X1 U401 ( .A(KEYINPUT12), .B(KEYINPUT97), .ZN(n499) );
  XOR2_X1 U402 ( .A(G140), .B(G104), .Z(n498) );
  NOR2_X1 U403 ( .A1(G237), .A2(G953), .ZN(n443) );
  OR2_X2 U404 ( .A1(n715), .A2(n720), .ZN(n368) );
  NAND2_X1 U405 ( .A1(n559), .A2(n558), .ZN(n365) );
  INV_X1 U406 ( .A(KEYINPUT83), .ZN(n407) );
  XOR2_X1 U407 ( .A(KEYINPUT5), .B(G146), .Z(n444) );
  XNOR2_X1 U408 ( .A(n512), .B(KEYINPUT7), .ZN(n417) );
  XNOR2_X1 U409 ( .A(KEYINPUT4), .B(G131), .ZN(n442) );
  XNOR2_X1 U410 ( .A(G146), .B(G125), .ZN(n466) );
  OR2_X1 U411 ( .A1(n717), .A2(n535), .ZN(n410) );
  NOR2_X1 U412 ( .A1(n716), .A2(KEYINPUT44), .ZN(n538) );
  XNOR2_X1 U413 ( .A(n480), .B(KEYINPUT85), .ZN(n481) );
  INV_X1 U414 ( .A(G469), .ZN(n412) );
  NOR2_X1 U415 ( .A1(n680), .A2(G902), .ZN(n454) );
  INV_X1 U416 ( .A(KEYINPUT22), .ZN(n430) );
  XNOR2_X1 U417 ( .A(n388), .B(n440), .ZN(n474) );
  XOR2_X1 U418 ( .A(KEYINPUT3), .B(G116), .Z(n440) );
  XNOR2_X1 U419 ( .A(n439), .B(n438), .ZN(n388) );
  INV_X1 U420 ( .A(G119), .ZN(n438) );
  XNOR2_X1 U421 ( .A(n360), .B(n358), .ZN(n510) );
  XNOR2_X1 U422 ( .A(n359), .B(KEYINPUT67), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n361), .B(n465), .ZN(n360) );
  INV_X1 U424 ( .A(KEYINPUT8), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n353), .B(n466), .ZN(n352) );
  NAND2_X1 U426 ( .A1(n708), .A2(G224), .ZN(n353) );
  NAND2_X1 U427 ( .A1(n355), .A2(n390), .ZN(n707) );
  XNOR2_X1 U428 ( .A(n580), .B(n348), .ZN(n355) );
  INV_X1 U429 ( .A(n624), .ZN(n391) );
  BUF_X1 U430 ( .A(n633), .Z(n389) );
  BUF_X1 U431 ( .A(n584), .Z(n393) );
  XOR2_X1 U432 ( .A(n509), .B(n508), .Z(n527) );
  NOR2_X1 U433 ( .A1(G902), .A2(n685), .ZN(n508) );
  XNOR2_X1 U434 ( .A(n474), .B(n384), .ZN(n702) );
  XNOR2_X1 U435 ( .A(n473), .B(n385), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n386), .B(G122), .ZN(n385) );
  INV_X1 U437 ( .A(KEYINPUT16), .ZN(n386) );
  INV_X1 U438 ( .A(KEYINPUT46), .ZN(n367) );
  OR2_X1 U439 ( .A1(G237), .A2(G902), .ZN(n483) );
  INV_X1 U440 ( .A(KEYINPUT99), .ZN(n518) );
  XNOR2_X1 U441 ( .A(G113), .B(G101), .ZN(n439) );
  NAND2_X1 U442 ( .A1(n476), .A2(G234), .ZN(n361) );
  INV_X1 U443 ( .A(KEYINPUT68), .ZN(n465) );
  INV_X1 U444 ( .A(KEYINPUT11), .ZN(n399) );
  XNOR2_X1 U445 ( .A(G131), .B(G143), .ZN(n497) );
  XOR2_X1 U446 ( .A(KEYINPUT15), .B(G902), .Z(n479) );
  XNOR2_X1 U447 ( .A(n408), .B(n407), .ZN(n406) );
  INV_X1 U448 ( .A(KEYINPUT69), .ZN(n382) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n487) );
  INV_X1 U450 ( .A(KEYINPUT1), .ZN(n411) );
  XNOR2_X1 U451 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U452 ( .A(n630), .B(n375), .ZN(n376) );
  INV_X1 U453 ( .A(KEYINPUT6), .ZN(n375) );
  XNOR2_X1 U454 ( .A(n427), .B(n425), .ZN(n587) );
  XNOR2_X1 U455 ( .A(n474), .B(n426), .ZN(n425) );
  XNOR2_X1 U456 ( .A(n450), .B(n446), .ZN(n427) );
  XNOR2_X1 U457 ( .A(G119), .B(G110), .ZN(n460) );
  XNOR2_X1 U458 ( .A(n416), .B(n415), .ZN(n593) );
  XNOR2_X1 U459 ( .A(n513), .B(n343), .ZN(n415) );
  XNOR2_X1 U460 ( .A(n511), .B(n417), .ZN(n416) );
  XNOR2_X1 U461 ( .A(n507), .B(n506), .ZN(n685) );
  XNOR2_X1 U462 ( .A(n706), .B(n398), .ZN(n507) );
  XNOR2_X1 U463 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U464 ( .A(n496), .B(n399), .ZN(n398) );
  XNOR2_X1 U465 ( .A(KEYINPUT75), .B(KEYINPUT90), .ZN(n437) );
  XNOR2_X1 U466 ( .A(n387), .B(G107), .ZN(n473) );
  XNOR2_X1 U467 ( .A(G104), .B(G110), .ZN(n387) );
  NAND2_X1 U468 ( .A1(n556), .A2(n433), .ZN(n565) );
  INV_X1 U469 ( .A(KEYINPUT100), .ZN(n429) );
  XNOR2_X1 U470 ( .A(n705), .B(n434), .ZN(n680) );
  XNOR2_X1 U471 ( .A(n436), .B(n435), .ZN(n434) );
  INV_X1 U472 ( .A(n473), .ZN(n435) );
  XNOR2_X1 U473 ( .A(n453), .B(n437), .ZN(n436) );
  XNOR2_X1 U474 ( .A(n351), .B(n432), .ZN(n478) );
  XNOR2_X1 U475 ( .A(n352), .B(n477), .ZN(n351) );
  NOR2_X1 U476 ( .A1(G952), .A2(n708), .ZN(n696) );
  INV_X1 U477 ( .A(KEYINPUT2), .ZN(n372) );
  INV_X1 U478 ( .A(n707), .ZN(n354) );
  INV_X1 U479 ( .A(n572), .ZN(n369) );
  NOR2_X1 U480 ( .A1(n532), .A2(n396), .ZN(n534) );
  OR2_X1 U481 ( .A1(n531), .A2(n397), .ZN(n396) );
  AND2_X1 U482 ( .A1(n550), .A2(n551), .ZN(n424) );
  XNOR2_X1 U483 ( .A(G107), .B(KEYINPUT9), .ZN(n343) );
  AND2_X1 U484 ( .A1(n402), .A2(n550), .ZN(n344) );
  AND2_X1 U485 ( .A1(n522), .A2(n599), .ZN(n345) );
  XNOR2_X1 U486 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n346) );
  XNOR2_X1 U487 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n347) );
  BUF_X1 U488 ( .A(n626), .Z(n394) );
  XNOR2_X1 U489 ( .A(KEYINPUT48), .B(KEYINPUT81), .ZN(n348) );
  INV_X1 U490 ( .A(n618), .ZN(n370) );
  NAND2_X1 U491 ( .A1(n349), .A2(n578), .ZN(n532) );
  NOR2_X2 U492 ( .A1(n350), .A2(n493), .ZN(n431) );
  NOR2_X1 U493 ( .A1(n565), .A2(n350), .ZN(n612) );
  XNOR2_X1 U494 ( .A(n486), .B(n485), .ZN(n350) );
  NAND2_X1 U495 ( .A1(n428), .A2(n354), .ZN(n373) );
  XNOR2_X2 U496 ( .A(n356), .B(KEYINPUT45), .ZN(n428) );
  NAND2_X1 U497 ( .A1(n357), .A2(n379), .ZN(n356) );
  NOR2_X1 U498 ( .A1(n381), .A2(n380), .ZN(n357) );
  NAND2_X1 U499 ( .A1(n510), .A2(G221), .ZN(n419) );
  AND2_X1 U500 ( .A1(n371), .A2(n370), .ZN(n622) );
  XNOR2_X1 U501 ( .A(n569), .B(n346), .ZN(n371) );
  XNOR2_X2 U502 ( .A(n373), .B(n372), .ZN(n666) );
  XNOR2_X2 U503 ( .A(n374), .B(n441), .ZN(n513) );
  XNOR2_X1 U504 ( .A(n374), .B(n475), .ZN(n432) );
  XNOR2_X2 U505 ( .A(n392), .B(G128), .ZN(n374) );
  XNOR2_X2 U506 ( .A(n447), .B(n448), .ZN(n630) );
  XNOR2_X2 U507 ( .A(n377), .B(KEYINPUT71), .ZN(n523) );
  NOR2_X2 U508 ( .A1(n633), .A2(n634), .ZN(n377) );
  INV_X1 U509 ( .A(n378), .ZN(n525) );
  NAND2_X1 U510 ( .A1(n378), .A2(n520), .ZN(n395) );
  XNOR2_X2 U511 ( .A(n431), .B(n347), .ZN(n378) );
  NAND2_X1 U512 ( .A1(n378), .A2(n405), .ZN(n404) );
  XNOR2_X1 U513 ( .A(n383), .B(n382), .ZN(n379) );
  NAND2_X1 U514 ( .A1(n406), .A2(n345), .ZN(n380) );
  XNOR2_X1 U515 ( .A(n409), .B(KEYINPUT64), .ZN(n381) );
  NAND2_X1 U516 ( .A1(n539), .A2(n607), .ZN(n383) );
  XNOR2_X1 U517 ( .A(n529), .B(n429), .ZN(n414) );
  XNOR2_X1 U518 ( .A(n540), .B(KEYINPUT103), .ZN(n421) );
  XNOR2_X1 U519 ( .A(n482), .B(n481), .ZN(n584) );
  NOR2_X1 U520 ( .A1(n391), .A2(n622), .ZN(n390) );
  NAND2_X1 U521 ( .A1(n433), .A2(n422), .ZN(n540) );
  NAND2_X1 U522 ( .A1(n536), .A2(n410), .ZN(n409) );
  BUF_X2 U523 ( .A(n653), .Z(n663) );
  INV_X1 U524 ( .A(n394), .ZN(n397) );
  NAND2_X1 U525 ( .A1(n663), .A2(KEYINPUT34), .ZN(n400) );
  NAND2_X1 U526 ( .A1(n525), .A2(KEYINPUT34), .ZN(n402) );
  INV_X1 U527 ( .A(KEYINPUT34), .ZN(n405) );
  XNOR2_X1 U528 ( .A(n524), .B(KEYINPUT33), .ZN(n653) );
  NAND2_X1 U529 ( .A1(n716), .A2(KEYINPUT44), .ZN(n408) );
  XNOR2_X2 U530 ( .A(n454), .B(n412), .ZN(n433) );
  XNOR2_X1 U531 ( .A(n420), .B(KEYINPUT73), .ZN(n549) );
  NAND2_X1 U532 ( .A1(n421), .A2(n545), .ZN(n420) );
  INV_X1 U533 ( .A(n634), .ZN(n422) );
  XNOR2_X1 U534 ( .A(n719), .B(KEYINPUT80), .ZN(n559) );
  NAND2_X1 U535 ( .A1(n568), .A2(n424), .ZN(n423) );
  AND2_X1 U536 ( .A1(n428), .A2(n476), .ZN(n699) );
  NAND2_X1 U537 ( .A1(n537), .A2(n530), .ZN(n536) );
  XNOR2_X1 U538 ( .A(KEYINPUT4), .B(KEYINPUT84), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U540 ( .A(n587), .B(KEYINPUT62), .ZN(n588) );
  XNOR2_X1 U541 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U542 ( .A(n687), .B(n686), .ZN(n688) );
  INV_X1 U543 ( .A(KEYINPUT125), .ZN(n597) );
  XNOR2_X1 U544 ( .A(G472), .B(KEYINPUT70), .ZN(n448) );
  XNOR2_X1 U545 ( .A(n443), .B(KEYINPUT72), .ZN(n503) );
  NAND2_X1 U546 ( .A1(n503), .A2(G210), .ZN(n445) );
  NOR2_X1 U547 ( .A1(n587), .A2(G902), .ZN(n447) );
  INV_X1 U548 ( .A(n459), .ZN(n449) );
  XOR2_X1 U549 ( .A(G101), .B(G146), .Z(n452) );
  INV_X2 U550 ( .A(G953), .ZN(n476) );
  NAND2_X1 U551 ( .A1(G227), .A2(n476), .ZN(n451) );
  XNOR2_X1 U552 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U553 ( .A1(n586), .A2(G234), .ZN(n456) );
  XNOR2_X1 U554 ( .A(KEYINPUT92), .B(KEYINPUT20), .ZN(n455) );
  XNOR2_X1 U555 ( .A(n456), .B(n455), .ZN(n468) );
  NAND2_X1 U556 ( .A1(n468), .A2(G221), .ZN(n457) );
  XNOR2_X1 U557 ( .A(n457), .B(KEYINPUT94), .ZN(n458) );
  XNOR2_X1 U558 ( .A(KEYINPUT21), .B(n458), .ZN(n627) );
  XNOR2_X1 U559 ( .A(n460), .B(n459), .ZN(n464) );
  XOR2_X1 U560 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n462) );
  XNOR2_X1 U561 ( .A(G128), .B(KEYINPUT91), .ZN(n461) );
  XNOR2_X1 U562 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U563 ( .A(n464), .B(n463), .Z(n467) );
  NAND2_X1 U564 ( .A1(n468), .A2(G217), .ZN(n470) );
  XNOR2_X1 U565 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n469) );
  BUF_X2 U566 ( .A(n476), .Z(n708) );
  XNOR2_X1 U567 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n477) );
  XNOR2_X1 U568 ( .A(n702), .B(n478), .ZN(n671) );
  NOR2_X1 U569 ( .A1(n671), .A2(n479), .ZN(n482) );
  NAND2_X1 U570 ( .A1(G210), .A2(n483), .ZN(n480) );
  NAND2_X1 U571 ( .A1(G214), .A2(n483), .ZN(n484) );
  XNOR2_X1 U572 ( .A(KEYINPUT86), .B(n484), .ZN(n643) );
  INV_X1 U573 ( .A(n643), .ZN(n546) );
  NOR2_X1 U574 ( .A1(n584), .A2(n546), .ZN(n486) );
  XNOR2_X1 U575 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n485) );
  XOR2_X1 U576 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n488) );
  XNOR2_X1 U577 ( .A(n488), .B(n487), .ZN(n490) );
  NAND2_X1 U578 ( .A1(G952), .A2(n490), .ZN(n660) );
  NOR2_X1 U579 ( .A1(G953), .A2(n660), .ZN(n544) );
  NOR2_X1 U580 ( .A1(G898), .A2(n708), .ZN(n489) );
  XOR2_X1 U581 ( .A(KEYINPUT88), .B(n489), .Z(n701) );
  NAND2_X1 U582 ( .A1(G902), .A2(n490), .ZN(n541) );
  NOR2_X1 U583 ( .A1(n701), .A2(n541), .ZN(n491) );
  NOR2_X1 U584 ( .A1(n544), .A2(n491), .ZN(n492) );
  XOR2_X1 U585 ( .A(KEYINPUT89), .B(n492), .Z(n493) );
  NOR2_X1 U586 ( .A1(n540), .A2(n525), .ZN(n494) );
  NAND2_X1 U587 ( .A1(n630), .A2(n494), .ZN(n602) );
  NOR2_X1 U588 ( .A1(n630), .A2(n523), .ZN(n640) );
  NAND2_X1 U589 ( .A1(n640), .A2(n378), .ZN(n495) );
  XOR2_X1 U590 ( .A(KEYINPUT31), .B(n495), .Z(n617) );
  NAND2_X1 U591 ( .A1(n602), .A2(n617), .ZN(n517) );
  XNOR2_X1 U592 ( .A(KEYINPUT13), .B(G475), .ZN(n509) );
  XNOR2_X1 U593 ( .A(G113), .B(G122), .ZN(n496) );
  XNOR2_X1 U594 ( .A(n498), .B(n497), .ZN(n502) );
  XNOR2_X1 U595 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U596 ( .A(n502), .B(n501), .ZN(n505) );
  NAND2_X1 U597 ( .A1(n503), .A2(G214), .ZN(n504) );
  NAND2_X1 U598 ( .A1(n510), .A2(G217), .ZN(n511) );
  XNOR2_X1 U599 ( .A(G116), .B(G122), .ZN(n512) );
  NOR2_X1 U600 ( .A1(G902), .A2(n593), .ZN(n515) );
  XNOR2_X1 U601 ( .A(KEYINPUT98), .B(G478), .ZN(n514) );
  XNOR2_X1 U602 ( .A(n515), .B(n514), .ZN(n526) );
  INV_X1 U603 ( .A(n526), .ZN(n516) );
  OR2_X1 U604 ( .A1(n527), .A2(n516), .ZN(n572) );
  NAND2_X1 U605 ( .A1(n527), .A2(n516), .ZN(n618) );
  NAND2_X1 U606 ( .A1(n572), .A2(n618), .ZN(n648) );
  XOR2_X1 U607 ( .A(KEYINPUT79), .B(n648), .Z(n560) );
  NAND2_X1 U608 ( .A1(n517), .A2(n560), .ZN(n522) );
  NAND2_X1 U609 ( .A1(n526), .A2(n527), .ZN(n646) );
  NOR2_X1 U610 ( .A1(n646), .A2(n627), .ZN(n519) );
  XNOR2_X1 U611 ( .A(n519), .B(n518), .ZN(n520) );
  NOR2_X1 U612 ( .A1(n573), .A2(n529), .ZN(n521) );
  NAND2_X1 U613 ( .A1(n521), .A2(n397), .ZN(n599) );
  NOR2_X1 U614 ( .A1(n527), .A2(n526), .ZN(n550) );
  XNOR2_X2 U615 ( .A(n528), .B(KEYINPUT35), .ZN(n716) );
  AND2_X1 U616 ( .A1(n394), .A2(KEYINPUT44), .ZN(n530) );
  INV_X1 U617 ( .A(KEYINPUT44), .ZN(n535) );
  INV_X1 U618 ( .A(n389), .ZN(n578) );
  XNOR2_X1 U619 ( .A(KEYINPUT76), .B(n573), .ZN(n531) );
  INV_X1 U620 ( .A(KEYINPUT32), .ZN(n533) );
  XNOR2_X1 U621 ( .A(n534), .B(n533), .ZN(n717) );
  NAND2_X1 U622 ( .A1(n537), .A2(n394), .ZN(n607) );
  AND2_X1 U623 ( .A1(n538), .A2(n717), .ZN(n539) );
  INV_X1 U624 ( .A(n393), .ZN(n551) );
  OR2_X1 U625 ( .A1(n708), .A2(n541), .ZN(n542) );
  NOR2_X1 U626 ( .A1(G900), .A2(n542), .ZN(n543) );
  NOR2_X1 U627 ( .A1(n544), .A2(n543), .ZN(n552) );
  INV_X1 U628 ( .A(n552), .ZN(n545) );
  NOR2_X1 U629 ( .A1(n630), .A2(n546), .ZN(n547) );
  XNOR2_X1 U630 ( .A(KEYINPUT30), .B(n547), .ZN(n548) );
  NOR2_X1 U631 ( .A1(n552), .A2(n627), .ZN(n553) );
  NAND2_X1 U632 ( .A1(n394), .A2(n553), .ZN(n575) );
  NOR2_X1 U633 ( .A1(n630), .A2(n575), .ZN(n555) );
  XOR2_X1 U634 ( .A(KEYINPUT28), .B(KEYINPUT105), .Z(n554) );
  XNOR2_X1 U635 ( .A(n555), .B(n554), .ZN(n556) );
  NAND2_X1 U636 ( .A1(n612), .A2(n648), .ZN(n557) );
  NAND2_X1 U637 ( .A1(KEYINPUT47), .A2(n557), .ZN(n558) );
  INV_X1 U638 ( .A(n560), .ZN(n561) );
  NOR2_X1 U639 ( .A1(n561), .A2(KEYINPUT47), .ZN(n562) );
  NAND2_X1 U640 ( .A1(n612), .A2(n562), .ZN(n563) );
  XNOR2_X1 U641 ( .A(KEYINPUT38), .B(n393), .ZN(n644) );
  NAND2_X1 U642 ( .A1(n644), .A2(n643), .ZN(n650) );
  NOR2_X1 U643 ( .A1(n646), .A2(n650), .ZN(n564) );
  XNOR2_X1 U644 ( .A(n564), .B(KEYINPUT41), .ZN(n662) );
  NOR2_X1 U645 ( .A1(n565), .A2(n662), .ZN(n567) );
  XOR2_X1 U646 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n566) );
  XNOR2_X1 U647 ( .A(n567), .B(n566), .ZN(n720) );
  NAND2_X1 U648 ( .A1(n568), .A2(n644), .ZN(n569) );
  XNOR2_X1 U649 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n570) );
  XNOR2_X1 U650 ( .A(n571), .B(n570), .ZN(n715) );
  XNOR2_X1 U651 ( .A(KEYINPUT101), .B(n572), .ZN(n611) );
  NAND2_X1 U652 ( .A1(n611), .A2(n573), .ZN(n574) );
  NOR2_X1 U653 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U654 ( .A1(n643), .A2(n576), .ZN(n581) );
  NOR2_X1 U655 ( .A1(n393), .A2(n581), .ZN(n577) );
  XNOR2_X1 U656 ( .A(n577), .B(KEYINPUT36), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n579), .A2(n578), .ZN(n621) );
  XOR2_X1 U658 ( .A(n581), .B(KEYINPUT102), .Z(n582) );
  NAND2_X1 U659 ( .A1(n582), .A2(n389), .ZN(n583) );
  XNOR2_X1 U660 ( .A(n583), .B(KEYINPUT43), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n585), .A2(n393), .ZN(n624) );
  NOR2_X4 U662 ( .A1(n666), .A2(n586), .ZN(n692) );
  NAND2_X1 U663 ( .A1(n692), .A2(G472), .ZN(n589) );
  INV_X1 U664 ( .A(KEYINPUT63), .ZN(n591) );
  XNOR2_X1 U665 ( .A(n592), .B(n591), .ZN(G57) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT124), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G478), .A2(n692), .ZN(n594) );
  XNOR2_X1 U668 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n598), .B(n597), .ZN(G63) );
  XNOR2_X1 U670 ( .A(G101), .B(KEYINPUT108), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(n599), .ZN(G3) );
  INV_X1 U672 ( .A(n611), .ZN(n615) );
  NOR2_X1 U673 ( .A1(n615), .A2(n602), .ZN(n601) );
  XOR2_X1 U674 ( .A(G104), .B(n601), .Z(G6) );
  NOR2_X1 U675 ( .A1(n602), .A2(n618), .ZN(n606) );
  XOR2_X1 U676 ( .A(KEYINPUT26), .B(KEYINPUT109), .Z(n604) );
  XNOR2_X1 U677 ( .A(G107), .B(KEYINPUT27), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U679 ( .A(n606), .B(n605), .ZN(G9) );
  XNOR2_X1 U680 ( .A(G110), .B(n607), .ZN(G12) );
  XOR2_X1 U681 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n609) );
  NAND2_X1 U682 ( .A1(n370), .A2(n612), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U684 ( .A(G128), .B(n610), .ZN(G30) );
  XOR2_X1 U685 ( .A(G146), .B(KEYINPUT111), .Z(n614) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(G48) );
  NOR2_X1 U688 ( .A1(n615), .A2(n617), .ZN(n616) );
  XOR2_X1 U689 ( .A(G113), .B(n616), .Z(G15) );
  NOR2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U691 ( .A(G116), .B(n619), .Z(G18) );
  XOR2_X1 U692 ( .A(G125), .B(KEYINPUT37), .Z(n620) );
  XNOR2_X1 U693 ( .A(n621), .B(n620), .ZN(G27) );
  XOR2_X1 U694 ( .A(G134), .B(n622), .Z(n623) );
  XNOR2_X1 U695 ( .A(KEYINPUT112), .B(n623), .ZN(G36) );
  XNOR2_X1 U696 ( .A(G140), .B(n624), .ZN(G42) );
  XNOR2_X1 U697 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n625), .B(KEYINPUT119), .ZN(n659) );
  NAND2_X1 U699 ( .A1(n627), .A2(n394), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(KEYINPUT113), .ZN(n629) );
  XNOR2_X1 U701 ( .A(KEYINPUT49), .B(n629), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U703 ( .A(KEYINPUT114), .B(n632), .ZN(n638) );
  NAND2_X1 U704 ( .A1(n634), .A2(n389), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n635), .B(KEYINPUT115), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n636), .B(KEYINPUT50), .ZN(n637) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U709 ( .A(KEYINPUT51), .B(n641), .Z(n642) );
  NOR2_X1 U710 ( .A1(n662), .A2(n642), .ZN(n657) );
  NOR2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n647), .B(KEYINPUT116), .ZN(n652) );
  INV_X1 U714 ( .A(n648), .ZN(n649) );
  NOR2_X1 U715 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U716 ( .A1(n652), .A2(n651), .ZN(n654) );
  NOR2_X1 U717 ( .A1(n654), .A2(n663), .ZN(n655) );
  XOR2_X1 U718 ( .A(KEYINPUT117), .B(n655), .Z(n656) );
  NOR2_X1 U719 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U720 ( .A(n659), .B(n658), .Z(n661) );
  NOR2_X1 U721 ( .A1(n661), .A2(n660), .ZN(n665) );
  NOR2_X1 U722 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U723 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U724 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U725 ( .A(KEYINPUT120), .B(n668), .ZN(n669) );
  NOR2_X1 U726 ( .A1(n669), .A2(G953), .ZN(n670) );
  XNOR2_X1 U727 ( .A(n670), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U728 ( .A(KEYINPUT55), .B(KEYINPUT77), .Z(n673) );
  XNOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n672) );
  XNOR2_X1 U730 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U731 ( .A(n671), .B(n674), .ZN(n676) );
  NAND2_X1 U732 ( .A1(G210), .A2(n692), .ZN(n675) );
  XNOR2_X1 U733 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U734 ( .A(n678), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U735 ( .A1(n692), .A2(G469), .ZN(n682) );
  XOR2_X1 U736 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n679) );
  XNOR2_X1 U737 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U738 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U739 ( .A1(n696), .A2(n683), .ZN(G54) );
  NAND2_X1 U740 ( .A1(n692), .A2(G475), .ZN(n687) );
  XOR2_X1 U741 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n684) );
  XNOR2_X1 U742 ( .A(n685), .B(n684), .ZN(n686) );
  XOR2_X1 U743 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n689) );
  XNOR2_X1 U744 ( .A(n690), .B(n689), .ZN(G60) );
  XNOR2_X1 U745 ( .A(n691), .B(KEYINPUT126), .ZN(n694) );
  NAND2_X1 U746 ( .A1(G217), .A2(n692), .ZN(n693) );
  XNOR2_X1 U747 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U748 ( .A1(n696), .A2(n695), .ZN(G66) );
  NAND2_X1 U749 ( .A1(G953), .A2(G224), .ZN(n697) );
  XNOR2_X1 U750 ( .A(KEYINPUT61), .B(n697), .ZN(n698) );
  AND2_X1 U751 ( .A1(n698), .A2(G898), .ZN(n700) );
  NOR2_X1 U752 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U753 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U754 ( .A(n704), .B(n703), .ZN(G69) );
  XOR2_X1 U755 ( .A(n706), .B(n705), .Z(n710) );
  XNOR2_X1 U756 ( .A(n707), .B(n710), .ZN(n709) );
  NAND2_X1 U757 ( .A1(n709), .A2(n708), .ZN(n714) );
  XNOR2_X1 U758 ( .A(G227), .B(n710), .ZN(n711) );
  NAND2_X1 U759 ( .A1(n711), .A2(G900), .ZN(n712) );
  NAND2_X1 U760 ( .A1(n712), .A2(G953), .ZN(n713) );
  NAND2_X1 U761 ( .A1(n714), .A2(n713), .ZN(G72) );
  XOR2_X1 U762 ( .A(n715), .B(G131), .Z(G33) );
  XOR2_X1 U763 ( .A(n716), .B(G122), .Z(G24) );
  XOR2_X1 U764 ( .A(G119), .B(n717), .Z(n718) );
  XNOR2_X1 U765 ( .A(KEYINPUT127), .B(n718), .ZN(G21) );
  XNOR2_X1 U766 ( .A(G143), .B(n719), .ZN(G45) );
  XOR2_X1 U767 ( .A(G137), .B(n720), .Z(G39) );
endmodule

