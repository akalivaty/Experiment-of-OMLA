

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  NOR2_X1 U324 ( .A1(n426), .A2(n520), .ZN(n574) );
  XNOR2_X1 U325 ( .A(n443), .B(n332), .ZN(n333) );
  XNOR2_X1 U326 ( .A(n343), .B(n298), .ZN(n301) );
  AND2_X1 U327 ( .A1(n445), .A2(n532), .ZN(n569) );
  XNOR2_X1 U328 ( .A(n427), .B(KEYINPUT55), .ZN(n445) );
  XOR2_X1 U329 ( .A(n358), .B(n357), .Z(n561) );
  XNOR2_X1 U330 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U331 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n292) );
  XOR2_X1 U332 ( .A(n320), .B(n319), .Z(n293) );
  XOR2_X1 U333 ( .A(KEYINPUT64), .B(n350), .Z(n294) );
  XOR2_X1 U334 ( .A(n352), .B(KEYINPUT78), .Z(n295) );
  XNOR2_X1 U335 ( .A(n455), .B(KEYINPUT25), .ZN(n456) );
  XNOR2_X1 U336 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U337 ( .A(G155GAT), .B(G22GAT), .Z(n362) );
  XNOR2_X1 U338 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n298) );
  XNOR2_X1 U339 ( .A(n345), .B(n292), .ZN(n332) );
  INV_X1 U340 ( .A(n431), .ZN(n305) );
  XNOR2_X1 U341 ( .A(n470), .B(KEYINPUT37), .ZN(n471) );
  NOR2_X1 U342 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U343 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U344 ( .A(n472), .B(n471), .ZN(n518) );
  XNOR2_X1 U345 ( .A(n308), .B(n307), .ZN(n310) );
  XNOR2_X1 U346 ( .A(n327), .B(n326), .ZN(n462) );
  INV_X1 U347 ( .A(KEYINPUT124), .ZN(n449) );
  NOR2_X1 U348 ( .A1(n538), .A2(n446), .ZN(n448) );
  XNOR2_X1 U349 ( .A(n339), .B(n338), .ZN(n508) );
  XNOR2_X1 U350 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U351 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U352 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  XOR2_X1 U353 ( .A(G99GAT), .B(G106GAT), .Z(n297) );
  XNOR2_X1 U354 ( .A(G85GAT), .B(KEYINPUT75), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n343) );
  XOR2_X1 U356 ( .A(G148GAT), .B(G78GAT), .Z(n316) );
  XNOR2_X1 U357 ( .A(n316), .B(KEYINPUT31), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n299), .B(KEYINPUT32), .ZN(n300) );
  XOR2_X1 U359 ( .A(n301), .B(n300), .Z(n308) );
  XNOR2_X1 U360 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n302), .B(KEYINPUT13), .ZN(n368) );
  XOR2_X1 U362 ( .A(G204GAT), .B(G176GAT), .Z(n304) );
  XNOR2_X1 U363 ( .A(G92GAT), .B(G64GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n336) );
  XNOR2_X1 U365 ( .A(n368), .B(n336), .ZN(n306) );
  XOR2_X1 U366 ( .A(G120GAT), .B(G71GAT), .Z(n431) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n580) );
  XOR2_X1 U369 ( .A(n580), .B(KEYINPUT41), .Z(n553) );
  XNOR2_X1 U370 ( .A(n553), .B(KEYINPUT109), .ZN(n538) );
  XOR2_X1 U371 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n312) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n416) );
  XOR2_X1 U374 ( .A(G211GAT), .B(G197GAT), .Z(n313) );
  XOR2_X1 U375 ( .A(KEYINPUT21), .B(n313), .Z(n337) );
  XNOR2_X1 U376 ( .A(n416), .B(n337), .ZN(n327) );
  XOR2_X1 U377 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n315) );
  XNOR2_X1 U378 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n314) );
  XNOR2_X1 U379 ( .A(n315), .B(n314), .ZN(n320) );
  XOR2_X1 U380 ( .A(n316), .B(n362), .Z(n318) );
  XNOR2_X1 U381 ( .A(G218GAT), .B(G106GAT), .ZN(n317) );
  XNOR2_X1 U382 ( .A(n318), .B(n317), .ZN(n319) );
  NAND2_X1 U383 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n293), .B(n321), .ZN(n322) );
  XOR2_X1 U385 ( .A(n322), .B(KEYINPUT88), .Z(n325) );
  XNOR2_X1 U386 ( .A(G162GAT), .B(G50GAT), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n323), .B(KEYINPUT76), .ZN(n340) );
  XNOR2_X1 U388 ( .A(n340), .B(KEYINPUT23), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U390 ( .A(G169GAT), .B(KEYINPUT86), .Z(n329) );
  XNOR2_X1 U391 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n330), .B(KEYINPUT19), .ZN(n443) );
  XNOR2_X1 U394 ( .A(G218GAT), .B(G36GAT), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n331), .B(G190GAT), .ZN(n345) );
  XOR2_X1 U396 ( .A(G8GAT), .B(G183GAT), .Z(n361) );
  XNOR2_X1 U397 ( .A(n333), .B(n361), .ZN(n335) );
  AND2_X1 U398 ( .A1(G226GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n339) );
  INV_X1 U400 ( .A(n508), .ZN(n522) );
  XNOR2_X1 U401 ( .A(n522), .B(KEYINPUT122), .ZN(n405) );
  XOR2_X1 U402 ( .A(KEYINPUT79), .B(G92GAT), .Z(n342) );
  XNOR2_X1 U403 ( .A(KEYINPUT77), .B(n340), .ZN(n341) );
  XNOR2_X1 U404 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U405 ( .A(n344), .B(n343), .Z(n347) );
  XNOR2_X1 U406 ( .A(G134GAT), .B(n345), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n358) );
  XOR2_X1 U408 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n349) );
  XNOR2_X1 U409 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n350) );
  NAND2_X1 U411 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n294), .B(n351), .ZN(n352) );
  XOR2_X1 U413 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n354) );
  XNOR2_X1 U414 ( .A(KEYINPUT70), .B(G43GAT), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U416 ( .A(G29GAT), .B(n355), .Z(n396) );
  XNOR2_X1 U417 ( .A(n396), .B(KEYINPUT80), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n295), .B(n356), .ZN(n357) );
  XNOR2_X1 U419 ( .A(KEYINPUT81), .B(n561), .ZN(n570) );
  XNOR2_X1 U420 ( .A(KEYINPUT36), .B(n570), .ZN(n585) );
  XOR2_X1 U421 ( .A(G78GAT), .B(G71GAT), .Z(n360) );
  XNOR2_X1 U422 ( .A(G1GAT), .B(G64GAT), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n375) );
  XOR2_X1 U424 ( .A(n362), .B(n361), .Z(n364) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U427 ( .A(G127GAT), .B(G15GAT), .Z(n430) );
  XOR2_X1 U428 ( .A(n365), .B(n430), .Z(n373) );
  XOR2_X1 U429 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n367) );
  XNOR2_X1 U430 ( .A(KEYINPUT83), .B(G211GAT), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n368), .B(KEYINPUT82), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n369), .B(KEYINPUT14), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n583) );
  NAND2_X1 U437 ( .A1(n585), .A2(n583), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n376), .B(KEYINPUT45), .ZN(n377) );
  NOR2_X1 U439 ( .A1(n580), .A2(n377), .ZN(n397) );
  XOR2_X1 U440 ( .A(KEYINPUT66), .B(KEYINPUT72), .Z(n379) );
  XNOR2_X1 U441 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U443 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n381) );
  XNOR2_X1 U444 ( .A(G22GAT), .B(G169GAT), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U446 ( .A(n383), .B(n382), .Z(n394) );
  XOR2_X1 U447 ( .A(KEYINPUT69), .B(KEYINPUT71), .Z(n385) );
  XNOR2_X1 U448 ( .A(G141GAT), .B(G15GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n392) );
  XOR2_X1 U450 ( .A(G113GAT), .B(G1GAT), .Z(n417) );
  XOR2_X1 U451 ( .A(G197GAT), .B(G8GAT), .Z(n387) );
  XNOR2_X1 U452 ( .A(G36GAT), .B(G50GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U454 ( .A(n417), .B(n388), .Z(n390) );
  NAND2_X1 U455 ( .A1(G229GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n575) );
  NAND2_X1 U460 ( .A1(n397), .A2(n575), .ZN(n403) );
  INV_X1 U461 ( .A(n575), .ZN(n563) );
  NAND2_X1 U462 ( .A1(n563), .A2(n553), .ZN(n398) );
  XNOR2_X1 U463 ( .A(KEYINPUT46), .B(n398), .ZN(n399) );
  NAND2_X1 U464 ( .A1(n399), .A2(n561), .ZN(n400) );
  NOR2_X1 U465 ( .A1(n583), .A2(n400), .ZN(n401) );
  XNOR2_X1 U466 ( .A(KEYINPUT47), .B(n401), .ZN(n402) );
  NAND2_X1 U467 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n404), .B(KEYINPUT48), .ZN(n530) );
  NAND2_X1 U469 ( .A1(n405), .A2(n530), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n406), .B(KEYINPUT54), .ZN(n426) );
  XOR2_X1 U471 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n408) );
  XNOR2_X1 U472 ( .A(G127GAT), .B(G155GAT), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n425) );
  XOR2_X1 U474 ( .A(G134GAT), .B(KEYINPUT0), .Z(n438) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(n438), .ZN(n409) );
  XNOR2_X1 U476 ( .A(n409), .B(G85GAT), .ZN(n413) );
  XOR2_X1 U477 ( .A(G148GAT), .B(G120GAT), .Z(n411) );
  XNOR2_X1 U478 ( .A(G162GAT), .B(G57GAT), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U480 ( .A(n413), .B(n412), .Z(n423) );
  XOR2_X1 U481 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n415) );
  XNOR2_X1 U482 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n421) );
  XOR2_X1 U484 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U485 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n520) );
  NAND2_X1 U490 ( .A1(n462), .A2(n574), .ZN(n427) );
  XOR2_X1 U491 ( .A(G176GAT), .B(G183GAT), .Z(n429) );
  XNOR2_X1 U492 ( .A(G113GAT), .B(G43GAT), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n442) );
  XOR2_X1 U494 ( .A(n431), .B(n430), .Z(n433) );
  XNOR2_X1 U495 ( .A(G190GAT), .B(G99GAT), .ZN(n432) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U497 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n435) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U500 ( .A(n437), .B(n436), .Z(n440) );
  XNOR2_X1 U501 ( .A(n438), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n532) );
  INV_X1 U505 ( .A(n532), .ZN(n511) );
  INV_X1 U506 ( .A(n569), .ZN(n446) );
  XNOR2_X1 U507 ( .A(KEYINPUT125), .B(KEYINPUT57), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n452) );
  XNOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n452), .B(n451), .ZN(G1349GAT) );
  NOR2_X1 U511 ( .A1(n532), .A2(n462), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n453), .B(KEYINPUT26), .ZN(n573) );
  XNOR2_X1 U513 ( .A(KEYINPUT27), .B(n522), .ZN(n463) );
  NAND2_X1 U514 ( .A1(n573), .A2(n463), .ZN(n459) );
  NAND2_X1 U515 ( .A1(n532), .A2(n522), .ZN(n454) );
  NAND2_X1 U516 ( .A1(n454), .A2(n462), .ZN(n457) );
  INV_X1 U517 ( .A(KEYINPUT94), .ZN(n455) );
  NAND2_X1 U518 ( .A1(n459), .A2(n458), .ZN(n460) );
  INV_X1 U519 ( .A(n520), .ZN(n503) );
  NAND2_X1 U520 ( .A1(n460), .A2(n503), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n461), .B(KEYINPUT95), .ZN(n466) );
  XNOR2_X1 U522 ( .A(KEYINPUT28), .B(n462), .ZN(n514) );
  INV_X1 U523 ( .A(n514), .ZN(n534) );
  AND2_X1 U524 ( .A1(n520), .A2(n463), .ZN(n529) );
  NAND2_X1 U525 ( .A1(n529), .A2(n511), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n534), .A2(n464), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT96), .ZN(n482) );
  NOR2_X1 U528 ( .A1(n482), .A2(n583), .ZN(n468) );
  XNOR2_X1 U529 ( .A(KEYINPUT102), .B(n468), .ZN(n469) );
  NAND2_X1 U530 ( .A1(n469), .A2(n585), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n470) );
  NOR2_X1 U532 ( .A1(n580), .A2(n575), .ZN(n483) );
  NAND2_X1 U533 ( .A1(n518), .A2(n483), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(KEYINPUT38), .ZN(n474) );
  XNOR2_X1 U535 ( .A(KEYINPUT105), .B(n474), .ZN(n499) );
  AND2_X1 U536 ( .A1(n499), .A2(n532), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n476) );
  INV_X1 U538 ( .A(G43GAT), .ZN(n475) );
  XOR2_X1 U539 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n486) );
  INV_X1 U540 ( .A(n583), .ZN(n479) );
  NOR2_X1 U541 ( .A1(n479), .A2(n570), .ZN(n480) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n480), .Z(n481) );
  NOR2_X1 U543 ( .A1(n482), .A2(n481), .ZN(n502) );
  NAND2_X1 U544 ( .A1(n483), .A2(n502), .ZN(n484) );
  XNOR2_X1 U545 ( .A(KEYINPUT97), .B(n484), .ZN(n492) );
  NAND2_X1 U546 ( .A1(n492), .A2(n520), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U548 ( .A(G1GAT), .B(n487), .Z(G1324GAT) );
  XOR2_X1 U549 ( .A(G8GAT), .B(KEYINPUT99), .Z(n489) );
  NAND2_X1 U550 ( .A1(n492), .A2(n522), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U553 ( .A1(n492), .A2(n532), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n494) );
  NAND2_X1 U556 ( .A1(n492), .A2(n534), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n495), .ZN(G1327GAT) );
  XOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .Z(n497) );
  NAND2_X1 U560 ( .A1(n499), .A2(n520), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NAND2_X1 U562 ( .A1(n499), .A2(n522), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT107), .Z(n501) );
  NAND2_X1 U565 ( .A1(n534), .A2(n499), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  NOR2_X1 U567 ( .A1(n563), .A2(n538), .ZN(n517) );
  NAND2_X1 U568 ( .A1(n517), .A2(n502), .ZN(n513) );
  NOR2_X1 U569 ( .A1(n513), .A2(n503), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT108), .B(KEYINPUT110), .Z(n505) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n508), .A2(n513), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NOR2_X1 U577 ( .A1(n511), .A2(n513), .ZN(n512) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U583 ( .A(KEYINPUT112), .B(n519), .Z(n525) );
  NAND2_X1 U584 ( .A1(n520), .A2(n525), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n525), .A2(n522), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n532), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n527) );
  NAND2_X1 U591 ( .A1(n534), .A2(n525), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT115), .Z(n536) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(n531), .Z(n550) );
  NAND2_X1 U597 ( .A1(n532), .A2(n550), .ZN(n533) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n546), .A2(n563), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  INV_X1 U601 ( .A(n546), .ZN(n537) );
  NOR2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n543) );
  NAND2_X1 U608 ( .A1(n546), .A2(n583), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n548) );
  NAND2_X1 U612 ( .A1(n546), .A2(n570), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U614 ( .A(G134GAT), .B(n549), .Z(G1343GAT) );
  NAND2_X1 U615 ( .A1(n550), .A2(n573), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT120), .B(n551), .Z(n559) );
  NAND2_X1 U617 ( .A1(n559), .A2(n563), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n559), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n583), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U626 ( .A(n559), .ZN(n560) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT123), .Z(n565) );
  NAND2_X1 U630 ( .A1(n569), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n567) );
  NAND2_X1 U633 ( .A1(n569), .A2(n583), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G183GAT), .B(n568), .ZN(G1350GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(n572), .ZN(G1351GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n579) );
  NOR2_X1 U640 ( .A1(n575), .A2(n579), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U645 ( .A(n579), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n586), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n586), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(KEYINPUT62), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

