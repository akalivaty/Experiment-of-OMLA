//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT69), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n191), .B1(new_n188), .B2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n193), .A2(KEYINPUT69), .A3(G116), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT70), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT69), .B1(new_n193), .B2(G116), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n191), .A2(new_n188), .A3(G119), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n189), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n187), .B1(new_n196), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n187), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n195), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n202), .A2(KEYINPUT72), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT72), .ZN(new_n206));
  AOI211_X1 g020(.A(KEYINPUT70), .B(new_n189), .C1(new_n198), .C2(new_n197), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n197), .A2(new_n198), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n200), .B1(new_n208), .B2(new_n190), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n203), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n204), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n206), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n205), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G134), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(G137), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT11), .A3(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(G137), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n216), .A2(new_n218), .A3(new_n222), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(KEYINPUT71), .A3(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G143), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n231), .B1(new_n236), .B2(G146), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT0), .A3(G128), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n235), .A3(new_n229), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT64), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n239), .A2(new_n240), .B1(new_n248), .B2(G128), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT66), .B(G143), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n230), .B(new_n251), .C1(new_n252), .C2(new_n229), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n236), .A2(G146), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(new_n230), .A4(new_n251), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n249), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n217), .A2(G134), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n219), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(KEYINPUT67), .A3(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI22_X1  g079(.A1(new_n228), .A2(new_n247), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n213), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n238), .A2(new_n246), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n221), .A2(KEYINPUT71), .A3(new_n223), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT71), .B1(new_n221), .B2(new_n223), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n249), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n256), .B1(new_n237), .B2(new_n251), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n229), .B1(new_n233), .B2(new_n235), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n275));
  NOR4_X1   g089(.A1(new_n274), .A2(new_n231), .A3(new_n275), .A4(KEYINPUT68), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n272), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n264), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n262), .B2(new_n259), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n268), .A2(new_n271), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT72), .B1(new_n202), .B2(new_n204), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n210), .A2(new_n206), .A3(new_n211), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n267), .A2(new_n284), .A3(KEYINPUT76), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n213), .A2(new_n286), .A3(new_n266), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(KEYINPUT28), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(G237), .A2(G953), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G210), .ZN(new_n290));
  INV_X1    g104(.A(G101), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n292), .B(new_n293), .Z(new_n294));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n213), .B2(new_n266), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n288), .A2(KEYINPUT29), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n224), .ZN(new_n300));
  OAI22_X1  g114(.A1(new_n258), .A2(new_n265), .B1(new_n247), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n210), .A2(new_n211), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n213), .B2(new_n266), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(KEYINPUT73), .A3(KEYINPUT28), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n295), .B1(new_n284), .B2(new_n303), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(new_n294), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n313), .B(new_n302), .C1(new_n312), .C2(new_n266), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n284), .ZN(new_n315));
  INV_X1    g129(.A(new_n294), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n280), .A2(new_n283), .B1(new_n302), .B2(new_n301), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n306), .B(new_n296), .C1(new_n320), .C2(new_n295), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n316), .B1(new_n321), .B2(new_n305), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n319), .B1(new_n322), .B2(new_n310), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n299), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G472), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n305), .B(new_n316), .C1(new_n307), .C2(new_n308), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n316), .A4(new_n305), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n314), .A2(new_n294), .A3(new_n284), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT31), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n314), .A2(KEYINPUT31), .A3(new_n294), .A4(new_n284), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n328), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(G472), .A2(G902), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(KEYINPUT32), .A3(new_n336), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n325), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n342), .A2(KEYINPUT16), .A3(G140), .ZN(new_n343));
  XNOR2_X1  g157(.A(G125), .B(G140), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(KEYINPUT16), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G146), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n229), .B(new_n343), .C1(KEYINPUT16), .C2(new_n344), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n250), .A2(G119), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT23), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n193), .A2(G128), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n351), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n250), .A2(KEYINPUT79), .A3(KEYINPUT23), .A4(G119), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n348), .B1(G110), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n250), .B2(G119), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n193), .A2(KEYINPUT77), .A3(G128), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n361), .A2(KEYINPUT78), .A3(new_n350), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT78), .B1(new_n361), .B2(new_n350), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT24), .B(G110), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n357), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n365), .B1(new_n362), .B2(new_n363), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n356), .A2(G110), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT80), .ZN(new_n369));
  INV_X1    g183(.A(new_n347), .ZN(new_n370));
  INV_X1    g184(.A(G140), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n342), .A2(G140), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT81), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT81), .B1(new_n372), .B2(new_n373), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n229), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n369), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT80), .B1(new_n367), .B2(new_n368), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n366), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT22), .B(G137), .ZN(new_n380));
  INV_X1    g194(.A(G953), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n381), .A2(G221), .A3(G234), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n380), .B(new_n382), .Z(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n366), .B(new_n383), .C1(new_n377), .C2(new_n378), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n298), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(KEYINPUT25), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(G234), .B2(new_n298), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n388), .A2(KEYINPUT25), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n385), .A2(new_n386), .A3(new_n298), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n385), .A2(new_n386), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n391), .A2(G902), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT83), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n399), .A3(new_n396), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n394), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n341), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n341), .A2(KEYINPUT84), .A3(new_n402), .ZN(new_n406));
  INV_X1    g220(.A(G475), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n233), .A2(new_n235), .B1(new_n289), .B2(G214), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n289), .A2(G143), .A3(G214), .ZN(new_n409));
  OAI21_X1  g223(.A(G131), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n289), .A2(G143), .A3(G214), .ZN(new_n412));
  INV_X1    g226(.A(G214), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n413), .A2(G237), .A3(G953), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n222), .B(new_n412), .C1(new_n252), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT17), .B(G131), .C1(new_n408), .C2(new_n409), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n348), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n344), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G146), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n376), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT18), .B(G131), .C1(new_n408), .C2(new_n409), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n408), .A2(new_n409), .ZN(new_n423));
  NAND2_X1  g237(.A1(KEYINPUT18), .A2(G131), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n418), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G113), .B(G122), .ZN(new_n428));
  INV_X1    g242(.A(G104), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n418), .A2(new_n430), .A3(new_n426), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n407), .B1(new_n434), .B2(new_n298), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n418), .A2(new_n430), .A3(new_n426), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n410), .A2(new_n415), .B1(G146), .B2(new_n345), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n374), .B2(new_n375), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n419), .A2(KEYINPUT19), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n229), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n426), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT91), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n430), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n376), .A2(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n422), .A2(new_n447), .B1(new_n438), .B2(new_n442), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT91), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n437), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(G475), .A2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n450), .A2(KEYINPUT20), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n431), .B1(new_n448), .B2(KEYINPUT91), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n444), .A2(new_n445), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n433), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n457), .B2(new_n451), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n436), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT92), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT20), .B1(new_n450), .B2(new_n452), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n454), .A3(new_n451), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n436), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n188), .A2(G122), .ZN(new_n468));
  INV_X1    g282(.A(G122), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G116), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n468), .A2(new_n470), .A3(G107), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(G116), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n472), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT95), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n470), .A2(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n475), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n471), .B1(new_n479), .B2(G107), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n236), .A2(G128), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n250), .A2(G143), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G134), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n215), .A3(new_n482), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT94), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n468), .A2(new_n470), .ZN(new_n491));
  INV_X1    g305(.A(G107), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(new_n471), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(KEYINPUT93), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(KEYINPUT93), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n481), .A2(KEYINPUT13), .A3(new_n482), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n497), .B(G134), .C1(KEYINPUT13), .C2(new_n481), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n495), .A2(new_n496), .A3(new_n498), .A4(new_n485), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT9), .B(G234), .Z(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(G217), .A3(new_n381), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n490), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n490), .B2(new_n499), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n298), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n506), .B(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(G234), .A2(G237), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(G952), .A3(new_n381), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT21), .B(G898), .Z(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(G902), .A3(G953), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n467), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G210), .B1(G237), .B2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n258), .A2(new_n342), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n247), .A2(G125), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n381), .A2(G224), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT89), .Z(new_n523));
  XNOR2_X1  g337(.A(new_n521), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G110), .B(G122), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n429), .A2(G107), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n429), .A2(G107), .ZN(new_n529));
  OAI21_X1  g343(.A(G101), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT3), .B1(new_n429), .B2(G107), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT3), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n492), .A3(G104), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n531), .A2(new_n533), .A3(new_n291), .A4(new_n527), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n196), .A2(new_n201), .A3(KEYINPUT5), .ZN(new_n536));
  OAI21_X1  g350(.A(G113), .B1(new_n190), .B2(KEYINPUT5), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI211_X1 g352(.A(new_n204), .B(new_n535), .C1(new_n536), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n533), .A3(new_n527), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G101), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT4), .A3(new_n534), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT4), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n543), .A3(G101), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n210), .B2(new_n211), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n526), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n535), .ZN(new_n548));
  INV_X1    g362(.A(new_n536), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n211), .B(new_n548), .C1(new_n549), .C2(new_n537), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n542), .A2(new_n544), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n302), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n552), .A3(new_n525), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n553), .A3(KEYINPUT6), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT6), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(new_n526), .C1(new_n539), .C2(new_n546), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n524), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n537), .B1(new_n199), .B2(KEYINPUT5), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n548), .B1(new_n558), .B2(new_n204), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n525), .B(KEYINPUT8), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n211), .B1(new_n549), .B2(new_n537), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n548), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n521), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT7), .A4(new_n522), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n562), .A2(new_n553), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n298), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n518), .B1(new_n557), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n567), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n524), .A2(new_n554), .A3(new_n556), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n517), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n571), .A3(KEYINPUT90), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT90), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n569), .A2(new_n573), .A3(new_n517), .A4(new_n570), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(G214), .B1(G237), .B2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G221), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n500), .B2(new_n298), .ZN(new_n580));
  INV_X1    g394(.A(G469), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n298), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G128), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n255), .A2(new_n230), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n254), .A2(new_n257), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n587), .B2(new_n535), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n277), .A2(KEYINPUT10), .A3(new_n548), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n551), .A2(new_n268), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n588), .A2(new_n589), .A3(new_n228), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n381), .A2(G227), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT85), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G140), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n591), .A2(KEYINPUT86), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT86), .B1(new_n591), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n271), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT87), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT87), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n603), .A3(new_n271), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI221_X4 g419(.A(new_n249), .B1(new_n534), .B2(new_n530), .C1(new_n254), .C2(new_n257), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n254), .A2(new_n257), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n585), .A2(new_n586), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n535), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n271), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT12), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(KEYINPUT12), .B(new_n224), .C1(new_n606), .C2(new_n609), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n591), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n599), .A2(new_n605), .B1(new_n615), .B2(new_n595), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n582), .B1(new_n616), .B2(G469), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n596), .B1(new_n605), .B2(new_n591), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT88), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n608), .B1(new_n273), .B2(new_n276), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n548), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n258), .A2(new_n535), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n228), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n613), .B(new_n619), .C1(new_n623), .C2(KEYINPUT12), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n619), .B1(new_n612), .B2(new_n613), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n591), .A2(new_n596), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n581), .B(new_n298), .C1(new_n618), .C2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n580), .B1(new_n617), .B2(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n516), .A2(new_n578), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n405), .A2(new_n406), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT96), .B(G101), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G3));
  INV_X1    g448(.A(G472), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n335), .B2(new_n298), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n336), .B2(new_n335), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n617), .A2(new_n629), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n401), .A2(new_n580), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n641), .B1(new_n504), .B2(new_n505), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n490), .A2(new_n499), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n501), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(KEYINPUT33), .A3(new_n503), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n507), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n507), .B(new_n298), .C1(new_n504), .C2(new_n505), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n507), .A2(new_n298), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n466), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT97), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n466), .A2(KEYINPUT97), .A3(new_n650), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n568), .A2(new_n571), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n515), .A2(new_n576), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n653), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n640), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT98), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  INV_X1    g477(.A(new_n658), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n664), .A2(new_n459), .A3(new_n510), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n640), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  OR3_X1    g482(.A1(new_n379), .A2(KEYINPUT36), .A3(new_n384), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n379), .B1(KEYINPUT36), .B2(new_n384), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n396), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n394), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n631), .A2(new_n637), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT99), .B(KEYINPUT100), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT37), .B(G110), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  OR2_X1    g491(.A1(new_n514), .A2(G900), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n512), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n459), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n509), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n630), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n655), .A2(new_n576), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n341), .A2(new_n684), .A3(new_n672), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  XNOR2_X1  g502(.A(new_n575), .B(KEYINPUT38), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n679), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n630), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n689), .B1(KEYINPUT40), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n466), .A2(new_n509), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n335), .A2(KEYINPUT32), .A3(new_n336), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT32), .B1(new_n335), .B2(new_n336), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n285), .A2(new_n316), .A3(new_n287), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(G472), .A3(new_n330), .ZN(new_n701));
  NAND2_X1  g515(.A1(G472), .A2(G902), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n703), .B(KEYINPUT101), .Z(new_n704));
  NAND2_X1  g518(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n672), .A2(new_n577), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n693), .A2(new_n696), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n252), .ZN(G45));
  INV_X1    g522(.A(new_n672), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n699), .B2(new_n325), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n464), .B1(new_n463), .B2(new_n436), .ZN(new_n711));
  AOI211_X1 g525(.A(KEYINPUT92), .B(new_n435), .C1(new_n461), .C2(new_n462), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n650), .B(new_n679), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT103), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n466), .A2(new_n715), .A3(new_n650), .A4(new_n679), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n710), .A2(new_n630), .A3(new_n686), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  NOR2_X1   g534(.A1(new_n625), .A2(new_n626), .ZN(new_n721));
  INV_X1    g535(.A(new_n627), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n600), .A2(new_n603), .A3(new_n271), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n603), .B1(new_n600), .B2(new_n271), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n591), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n721), .A2(new_n722), .B1(new_n725), .B2(new_n595), .ZN(new_n726));
  OAI21_X1  g540(.A(G469), .B1(new_n726), .B2(G902), .ZN(new_n727));
  INV_X1    g541(.A(new_n580), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n629), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT104), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n727), .A2(new_n731), .A3(new_n728), .A4(new_n629), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n401), .B1(new_n699), .B2(new_n325), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n659), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  NAND3_X1  g552(.A1(new_n734), .A2(new_n735), .A3(new_n665), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND4_X1  g554(.A1(new_n710), .A2(new_n734), .A3(new_n516), .A4(new_n686), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  INV_X1    g556(.A(new_n695), .ZN(new_n743));
  INV_X1    g557(.A(new_n336), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n288), .A2(new_n296), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n316), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n744), .B1(new_n746), .B2(new_n334), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n636), .A2(new_n401), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n734), .A2(new_n658), .A3(new_n743), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  NAND3_X1  g564(.A1(new_n730), .A2(new_n686), .A3(new_n732), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n335), .A2(new_n298), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n747), .B1(new_n752), .B2(G472), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n714), .A3(new_n716), .A4(new_n672), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n342), .ZN(G27));
  INV_X1    g570(.A(KEYINPUT105), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(KEYINPUT42), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n577), .B1(new_n572), .B2(new_n574), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n630), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n341), .A2(new_n402), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n758), .B1(new_n761), .B2(new_n717), .ZN(new_n762));
  INV_X1    g576(.A(new_n758), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n735), .A2(new_n718), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  XNOR2_X1  g580(.A(new_n682), .B(KEYINPUT106), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n735), .A2(new_n760), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  OR2_X1    g583(.A1(new_n616), .A2(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n616), .A2(KEYINPUT45), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(G469), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n582), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n629), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT46), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n728), .B(new_n691), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT107), .ZN(new_n778));
  INV_X1    g592(.A(new_n650), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n466), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT43), .Z(new_n781));
  OR2_X1    g595(.A1(new_n637), .A2(new_n709), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n783), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n778), .A2(new_n759), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  OAI21_X1  g601(.A(new_n728), .B1(new_n775), .B2(new_n776), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n718), .A3(new_n759), .A4(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n341), .A3(new_n402), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n371), .ZN(G42));
  NAND2_X1  g607(.A1(new_n381), .A2(G952), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n781), .A2(new_n512), .ZN(new_n795));
  INV_X1    g609(.A(new_n759), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n733), .A2(new_n796), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n672), .A2(new_n795), .A3(new_n753), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n705), .A2(new_n512), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n797), .A3(new_n402), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n466), .A3(new_n650), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n748), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n781), .A2(new_n512), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT111), .B1(new_n733), .B2(new_n576), .ZN(new_n805));
  OR3_X1    g619(.A1(new_n733), .A2(KEYINPUT111), .A3(new_n576), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n689), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n802), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT51), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n807), .B(new_n808), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(KEYINPUT112), .A3(new_n802), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n727), .A2(new_n629), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n728), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n789), .B2(new_n790), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n796), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n804), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(KEYINPUT110), .A3(new_n804), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n813), .A2(new_n815), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n820), .B1(KEYINPUT113), .B2(new_n802), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n802), .A2(KEYINPUT113), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n814), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT51), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n794), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n653), .A2(new_n654), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n800), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n730), .A2(new_n686), .A3(new_n732), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n804), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  INV_X1    g648(.A(new_n575), .ZN(new_n835));
  INV_X1    g649(.A(new_n657), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n651), .B1(new_n466), .B2(new_n510), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n640), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n632), .A2(new_n673), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n341), .A2(new_n510), .A3(new_n681), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n753), .A2(new_n714), .A3(new_n716), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n709), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n764), .A2(new_n762), .B1(new_n842), .B2(new_n760), .ZN(new_n843));
  INV_X1    g657(.A(new_n659), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n341), .A2(new_n402), .A3(new_n732), .A4(new_n730), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n341), .A2(new_n516), .A3(new_n672), .A4(new_n686), .ZN(new_n846));
  OAI22_X1  g660(.A1(new_n844), .A2(new_n845), .B1(new_n846), .B2(new_n733), .ZN(new_n847));
  INV_X1    g661(.A(new_n665), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n748), .A2(new_n730), .A3(new_n743), .A4(new_n732), .ZN(new_n849));
  OAI22_X1  g663(.A1(new_n845), .A2(new_n848), .B1(new_n849), .B2(new_n664), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n839), .A2(new_n843), .A3(new_n851), .A4(new_n768), .ZN(new_n852));
  INV_X1    g666(.A(new_n754), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n832), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n394), .B(new_n671), .C1(KEYINPUT109), .C2(new_n679), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n679), .A2(KEYINPUT109), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n695), .A2(new_n855), .A3(new_n685), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n705), .A3(new_n630), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n719), .A2(new_n854), .A3(new_n687), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n341), .A2(new_n684), .A3(new_n672), .A4(new_n686), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n755), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n862), .A2(new_n863), .A3(new_n719), .A4(new_n858), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n834), .B1(new_n852), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n840), .A2(new_n841), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n672), .A3(new_n760), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n765), .A2(new_n768), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n741), .A2(new_n749), .A3(new_n736), .A4(new_n739), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n632), .A2(new_n673), .A3(new_n838), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n860), .A2(new_n864), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT53), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n866), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT54), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n829), .A2(new_n831), .A3(new_n833), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n795), .A2(new_n735), .A3(new_n797), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT48), .Z(new_n883));
  OAI22_X1  g697(.A1(new_n881), .A2(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n639), .A2(new_n576), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT108), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(new_n780), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n816), .B(KEYINPUT49), .Z(new_n888));
  AOI21_X1  g702(.A(new_n705), .B1(new_n885), .B2(KEYINPUT108), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n887), .A2(new_n689), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n884), .A2(new_n890), .ZN(G75));
  NOR2_X1   g705(.A1(new_n381), .A2(G952), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT115), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n876), .A2(new_n298), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(G210), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n554), .A2(new_n556), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n524), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n894), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT114), .B1(new_n875), .B2(G902), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT114), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n902), .B(new_n298), .C1(new_n866), .C2(new_n874), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n518), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n900), .B1(new_n904), .B2(new_n906), .ZN(G51));
  XOR2_X1   g721(.A(new_n772), .B(KEYINPUT116), .Z(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n901), .B2(new_n903), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT117), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n911), .B(new_n908), .C1(new_n901), .C2(new_n903), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n773), .A2(KEYINPUT57), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n773), .A2(KEYINPUT57), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n879), .A2(new_n877), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n910), .B(new_n912), .C1(new_n915), .C2(new_n726), .ZN(new_n916));
  INV_X1    g730(.A(new_n892), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(G54));
  AND2_X1   g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n901), .B2(new_n903), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n450), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n457), .B(new_n919), .C1(new_n901), .C2(new_n903), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n917), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n921), .A2(KEYINPUT118), .A3(new_n917), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(G60));
  XNOR2_X1  g741(.A(new_n649), .B(KEYINPUT119), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n642), .B(new_n645), .C1(new_n880), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n642), .A2(new_n645), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n877), .A2(new_n932), .A3(new_n879), .A4(new_n929), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n893), .B1(new_n931), .B2(new_n933), .ZN(G63));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n875), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n669), .A2(new_n670), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT120), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n894), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n395), .B(KEYINPUT121), .Z(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g757(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n943), .B(new_n944), .Z(G66));
  NAND2_X1  g759(.A1(new_n513), .A2(G224), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(G953), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n871), .A2(new_n870), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(G953), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n897), .B1(G898), .B2(new_n381), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G69));
  OAI21_X1  g765(.A(new_n313), .B1(new_n312), .B2(new_n266), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n440), .A2(new_n441), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n862), .A2(new_n719), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n707), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n957), .A2(new_n707), .A3(KEYINPUT62), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n792), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n964));
  AOI211_X1 g778(.A(new_n796), .B(new_n692), .C1(new_n964), .C2(new_n837), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n837), .A2(new_n964), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(new_n405), .A3(new_n406), .A4(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n786), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n962), .A2(new_n963), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n963), .B1(new_n962), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n955), .B1(new_n971), .B2(G953), .ZN(new_n972));
  NAND2_X1  g786(.A1(G227), .A2(G900), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(G953), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n381), .A2(G900), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT125), .Z(new_n976));
  NOR2_X1   g790(.A1(new_n792), .A2(new_n956), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n784), .A2(new_n759), .A3(new_n785), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n735), .A2(new_n686), .A3(new_n743), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI22_X1  g794(.A1(new_n980), .A2(new_n778), .B1(new_n764), .B2(new_n762), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n977), .A2(new_n768), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n976), .B1(new_n982), .B2(G953), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n954), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n972), .A2(new_n974), .A3(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(G953), .B(new_n973), .C1(new_n983), .C2(new_n955), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(G72));
  NOR4_X1   g801(.A1(new_n969), .A2(new_n970), .A3(new_n870), .A4(new_n871), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n702), .B(KEYINPUT63), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n294), .B(new_n315), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n977), .A2(new_n981), .A3(new_n768), .A4(new_n948), .ZN(new_n992));
  INV_X1    g806(.A(new_n989), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n294), .B(new_n315), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n991), .B1(new_n994), .B2(new_n892), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n993), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n316), .ZN(new_n997));
  OAI211_X1 g811(.A(KEYINPUT126), .B(new_n917), .C1(new_n997), .C2(new_n315), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n317), .A2(new_n330), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n875), .A2(new_n993), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT127), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n990), .A2(new_n999), .A3(new_n1002), .ZN(G57));
endmodule


