

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U555 ( .A1(n587), .A2(G2104), .ZN(n932) );
  INV_X1 U556 ( .A(n695), .ZN(n673) );
  NAND2_X1 U557 ( .A1(n695), .A2(G8), .ZN(n694) );
  NOR2_X1 U558 ( .A1(n661), .A2(n660), .ZN(n1030) );
  NAND2_X1 U559 ( .A1(n560), .A2(n734), .ZN(n695) );
  NAND2_X1 U560 ( .A1(n537), .A2(n536), .ZN(n530) );
  NAND2_X1 U561 ( .A1(n530), .A2(n525), .ZN(n677) );
  XNOR2_X1 U562 ( .A(n733), .B(KEYINPUT91), .ZN(n560) );
  NOR2_X1 U563 ( .A1(n544), .A2(n729), .ZN(n543) );
  INV_X1 U564 ( .A(n1017), .ZN(n544) );
  INV_X1 U565 ( .A(KEYINPUT102), .ZN(n554) );
  NAND2_X1 U566 ( .A1(n553), .A2(n550), .ZN(n549) );
  NAND2_X1 U567 ( .A1(n780), .A2(n551), .ZN(n550) );
  NAND2_X1 U568 ( .A1(n555), .A2(n554), .ZN(n553) );
  NAND2_X1 U569 ( .A1(n552), .A2(n554), .ZN(n551) );
  NOR2_X1 U570 ( .A1(n533), .A2(n532), .ZN(n531) );
  INV_X1 U571 ( .A(n534), .ZN(n532) );
  XNOR2_X1 U572 ( .A(n703), .B(KEYINPUT31), .ZN(n704) );
  INV_X1 U573 ( .A(KEYINPUT96), .ZN(n703) );
  NAND2_X1 U574 ( .A1(n565), .A2(n564), .ZN(n566) );
  INV_X1 U575 ( .A(n571), .ZN(n552) );
  INV_X1 U576 ( .A(n780), .ZN(n555) );
  NAND2_X1 U577 ( .A1(n542), .A2(n540), .ZN(n539) );
  NOR2_X1 U578 ( .A1(n694), .A2(n541), .ZN(n540) );
  NOR2_X1 U579 ( .A1(n1017), .A2(KEYINPUT99), .ZN(n541) );
  NAND2_X1 U580 ( .A1(n526), .A2(n558), .ZN(n733) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n834) );
  INV_X1 U582 ( .A(KEYINPUT65), .ZN(n577) );
  XNOR2_X1 U583 ( .A(KEYINPUT23), .B(KEYINPUT67), .ZN(n588) );
  INV_X1 U584 ( .A(KEYINPUT17), .ZN(n591) );
  NOR2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n592) );
  INV_X1 U586 ( .A(G2105), .ZN(n587) );
  AND2_X1 U587 ( .A1(n556), .A2(n549), .ZN(n548) );
  AND2_X1 U588 ( .A1(n780), .A2(n554), .ZN(n523) );
  NOR2_X1 U589 ( .A1(n567), .A2(KEYINPUT29), .ZN(n524) );
  XNOR2_X2 U590 ( .A(n592), .B(n591), .ZN(n739) );
  AND2_X1 U591 ( .A1(n534), .A2(n535), .ZN(n525) );
  NOR2_X1 U592 ( .A1(n599), .A2(n559), .ZN(n526) );
  XOR2_X1 U593 ( .A(n699), .B(n698), .Z(n527) );
  AND2_X1 U594 ( .A1(n562), .A2(n561), .ZN(n528) );
  INV_X1 U595 ( .A(n732), .ZN(n557) );
  AND2_X1 U596 ( .A1(n571), .A2(KEYINPUT102), .ZN(n529) );
  INV_X1 U597 ( .A(KEYINPUT99), .ZN(n729) );
  NAND2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n535), .A2(n942), .ZN(n533) );
  NAND2_X1 U600 ( .A1(n664), .A2(KEYINPUT64), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n665), .A2(KEYINPUT64), .ZN(n535) );
  INV_X1 U602 ( .A(n665), .ZN(n536) );
  NOR2_X1 U603 ( .A1(n664), .A2(KEYINPUT64), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n676), .ZN(n679) );
  NOR2_X1 U605 ( .A1(n545), .A2(n539), .ZN(n730) );
  NAND2_X1 U606 ( .A1(n546), .A2(n543), .ZN(n542) );
  NOR2_X1 U607 ( .A1(n546), .A2(KEYINPUT99), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n728), .B(KEYINPUT98), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n782) );
  NAND2_X1 U610 ( .A1(n732), .A2(n523), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n557), .A2(n529), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n599), .A2(n600), .ZN(G160) );
  INV_X1 U613 ( .A(n600), .ZN(n558) );
  INV_X1 U614 ( .A(G40), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n684), .A2(n524), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n563), .A2(n689), .ZN(n562) );
  INV_X1 U617 ( .A(n688), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n684), .A2(n683), .ZN(n564) );
  AND2_X1 U619 ( .A1(n688), .A2(KEYINPUT29), .ZN(n565) );
  NAND2_X1 U620 ( .A1(n528), .A2(n566), .ZN(n568) );
  INV_X1 U621 ( .A(n683), .ZN(n567) );
  NAND2_X1 U622 ( .A1(n568), .A2(n693), .ZN(n707) );
  NAND2_X1 U623 ( .A1(n715), .A2(n714), .ZN(n717) );
  OR2_X1 U624 ( .A1(n694), .A2(n767), .ZN(n569) );
  XOR2_X1 U625 ( .A(KEYINPUT6), .B(n584), .Z(n570) );
  AND2_X1 U626 ( .A1(n768), .A2(n569), .ZN(n571) );
  XNOR2_X1 U627 ( .A(KEYINPUT30), .B(KEYINPUT95), .ZN(n698) );
  INV_X1 U628 ( .A(KEYINPUT32), .ZN(n716) );
  NAND2_X1 U629 ( .A1(n825), .A2(G54), .ZN(n667) );
  INV_X1 U630 ( .A(G2104), .ZN(n595) );
  XOR2_X1 U631 ( .A(n672), .B(KEYINPUT15), .Z(n942) );
  NAND2_X1 U632 ( .A1(n739), .A2(G137), .ZN(n593) );
  XNOR2_X1 U633 ( .A(KEYINPUT7), .B(n586), .ZN(G168) );
  NAND2_X1 U634 ( .A1(n834), .A2(G89), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  XOR2_X1 U636 ( .A(G543), .B(KEYINPUT0), .Z(n576) );
  INV_X1 U637 ( .A(G651), .ZN(n580) );
  NOR2_X2 U638 ( .A1(n576), .A2(n580), .ZN(n830) );
  NAND2_X1 U639 ( .A1(G76), .A2(n830), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT5), .B(n575), .ZN(n585) );
  NOR2_X1 U642 ( .A1(G651), .A2(n576), .ZN(n578) );
  XNOR2_X2 U643 ( .A(n578), .B(n577), .ZN(n825) );
  NAND2_X1 U644 ( .A1(n825), .A2(G51), .ZN(n579) );
  XOR2_X1 U645 ( .A(KEYINPUT75), .B(n579), .Z(n583) );
  NOR2_X1 U646 ( .A1(G543), .A2(n580), .ZN(n581) );
  XOR2_X2 U647 ( .A(KEYINPUT1), .B(n581), .Z(n826) );
  NAND2_X1 U648 ( .A1(n826), .A2(G63), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n570), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G101), .A2(n932), .ZN(n590) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT66), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n590), .B(n589), .ZN(n594) );
  NAND2_X1 U654 ( .A1(n594), .A2(n593), .ZN(n600) );
  AND2_X1 U655 ( .A1(n595), .A2(G2105), .ZN(n926) );
  NAND2_X1 U656 ( .A1(n926), .A2(G125), .ZN(n598) );
  NAND2_X1 U657 ( .A1(G2105), .A2(G2104), .ZN(n596) );
  XOR2_X1 U658 ( .A(KEYINPUT68), .B(n596), .Z(n735) );
  NAND2_X1 U659 ( .A1(G113), .A2(n735), .ZN(n597) );
  NAND2_X1 U660 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G138), .A2(n739), .ZN(n602) );
  NAND2_X1 U662 ( .A1(G102), .A2(n932), .ZN(n601) );
  NAND2_X1 U663 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U664 ( .A1(n926), .A2(G126), .ZN(n604) );
  NAND2_X1 U665 ( .A1(G114), .A2(n735), .ZN(n603) );
  NAND2_X1 U666 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U667 ( .A1(n606), .A2(n605), .ZN(G164) );
  NAND2_X1 U668 ( .A1(n830), .A2(G78), .ZN(n607) );
  XNOR2_X1 U669 ( .A(n607), .B(KEYINPUT72), .ZN(n609) );
  NAND2_X1 U670 ( .A1(G91), .A2(n834), .ZN(n608) );
  NAND2_X1 U671 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U672 ( .A(KEYINPUT73), .B(n610), .ZN(n614) );
  NAND2_X1 U673 ( .A1(G53), .A2(n825), .ZN(n612) );
  NAND2_X1 U674 ( .A1(G65), .A2(n826), .ZN(n611) );
  AND2_X1 U675 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U676 ( .A1(n614), .A2(n613), .ZN(G299) );
  NAND2_X1 U677 ( .A1(G90), .A2(n834), .ZN(n616) );
  NAND2_X1 U678 ( .A1(G77), .A2(n830), .ZN(n615) );
  NAND2_X1 U679 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U680 ( .A(KEYINPUT9), .B(n617), .ZN(n621) );
  NAND2_X1 U681 ( .A1(G52), .A2(n825), .ZN(n619) );
  NAND2_X1 U682 ( .A1(G64), .A2(n826), .ZN(n618) );
  AND2_X1 U683 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U684 ( .A1(n621), .A2(n620), .ZN(G301) );
  INV_X1 U685 ( .A(G301), .ZN(G171) );
  XOR2_X1 U686 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U687 ( .A1(n834), .A2(G88), .ZN(n624) );
  NAND2_X1 U688 ( .A1(G62), .A2(n826), .ZN(n622) );
  XOR2_X1 U689 ( .A(KEYINPUT83), .B(n622), .Z(n623) );
  NAND2_X1 U690 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U691 ( .A1(G50), .A2(n825), .ZN(n626) );
  NAND2_X1 U692 ( .A1(G75), .A2(n830), .ZN(n625) );
  NAND2_X1 U693 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U694 ( .A1(n628), .A2(n627), .ZN(G166) );
  INV_X1 U695 ( .A(G166), .ZN(G303) );
  NAND2_X1 U696 ( .A1(G49), .A2(n825), .ZN(n630) );
  NAND2_X1 U697 ( .A1(G87), .A2(n576), .ZN(n629) );
  NAND2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U699 ( .A1(n826), .A2(n631), .ZN(n634) );
  NAND2_X1 U700 ( .A1(G74), .A2(G651), .ZN(n632) );
  XOR2_X1 U701 ( .A(KEYINPUT81), .B(n632), .Z(n633) );
  NAND2_X1 U702 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U703 ( .A1(G73), .A2(n830), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n635), .B(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U705 ( .A1(G48), .A2(n825), .ZN(n637) );
  NAND2_X1 U706 ( .A1(G61), .A2(n826), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n834), .A2(G86), .ZN(n638) );
  XOR2_X1 U709 ( .A(KEYINPUT82), .B(n638), .Z(n639) );
  NOR2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U712 ( .A1(n825), .A2(G47), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n643), .B(KEYINPUT70), .ZN(n645) );
  NAND2_X1 U714 ( .A1(G60), .A2(n826), .ZN(n644) );
  NAND2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n650) );
  NAND2_X1 U716 ( .A1(G85), .A2(n834), .ZN(n647) );
  NAND2_X1 U717 ( .A1(G72), .A2(n830), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U719 ( .A(KEYINPUT69), .B(n648), .Z(n649) );
  NOR2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U721 ( .A(KEYINPUT71), .B(n651), .ZN(G290) );
  NOR2_X1 U722 ( .A1(G164), .A2(G1384), .ZN(n734) );
  NAND2_X1 U723 ( .A1(G1996), .A2(n673), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n652), .B(KEYINPUT26), .ZN(n662) );
  NAND2_X1 U725 ( .A1(n834), .A2(G81), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n653), .B(KEYINPUT12), .ZN(n655) );
  NAND2_X1 U727 ( .A1(G68), .A2(n830), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n656), .B(KEYINPUT13), .ZN(n658) );
  NAND2_X1 U730 ( .A1(G43), .A2(n825), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n826), .A2(G56), .ZN(n659) );
  XOR2_X1 U733 ( .A(KEYINPUT14), .B(n659), .Z(n660) );
  NAND2_X1 U734 ( .A1(n662), .A2(n1030), .ZN(n665) );
  NAND2_X1 U735 ( .A1(G1341), .A2(n695), .ZN(n663) );
  XNOR2_X1 U736 ( .A(KEYINPUT93), .B(n663), .ZN(n664) );
  NAND2_X1 U737 ( .A1(G66), .A2(n826), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U739 ( .A1(G92), .A2(n834), .ZN(n669) );
  NAND2_X1 U740 ( .A1(G79), .A2(n830), .ZN(n668) );
  NAND2_X1 U741 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  INV_X1 U743 ( .A(n942), .ZN(n1027) );
  NOR2_X1 U744 ( .A1(n673), .A2(G1348), .ZN(n675) );
  NOR2_X1 U745 ( .A1(n695), .A2(G2067), .ZN(n674) );
  NOR2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U747 ( .A1(n677), .A2(n1027), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n684) );
  INV_X1 U749 ( .A(G299), .ZN(n686) );
  NAND2_X1 U750 ( .A1(n673), .A2(G2072), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n680), .B(KEYINPUT27), .ZN(n682) );
  INV_X1 U752 ( .A(G1956), .ZN(n890) );
  NOR2_X1 U753 ( .A1(n890), .A2(n673), .ZN(n681) );
  NOR2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n683) );
  NOR2_X1 U756 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U757 ( .A(n687), .B(KEYINPUT28), .Z(n688) );
  INV_X1 U758 ( .A(KEYINPUT29), .ZN(n689) );
  XOR2_X1 U759 ( .A(KEYINPUT25), .B(G2078), .Z(n955) );
  NAND2_X1 U760 ( .A1(n673), .A2(n955), .ZN(n691) );
  NAND2_X1 U761 ( .A1(G1961), .A2(n695), .ZN(n690) );
  NAND2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U763 ( .A(KEYINPUT92), .B(n692), .Z(n700) );
  NAND2_X1 U764 ( .A1(n700), .A2(G171), .ZN(n693) );
  NOR2_X1 U765 ( .A1(G1966), .A2(n694), .ZN(n719) );
  NOR2_X1 U766 ( .A1(G2084), .A2(n695), .ZN(n721) );
  NOR2_X1 U767 ( .A1(n719), .A2(n721), .ZN(n696) );
  XNOR2_X1 U768 ( .A(n696), .B(KEYINPUT94), .ZN(n697) );
  NAND2_X1 U769 ( .A1(n697), .A2(G8), .ZN(n699) );
  NOR2_X1 U770 ( .A1(G168), .A2(n527), .ZN(n702) );
  NOR2_X1 U771 ( .A1(G171), .A2(n700), .ZN(n701) );
  NOR2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n705) );
  XNOR2_X1 U773 ( .A(n705), .B(n704), .ZN(n706) );
  NAND2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n718) );
  AND2_X1 U775 ( .A1(G286), .A2(G8), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n718), .A2(n708), .ZN(n715) );
  INV_X1 U777 ( .A(G8), .ZN(n713) );
  NOR2_X1 U778 ( .A1(G1971), .A2(n694), .ZN(n710) );
  NOR2_X1 U779 ( .A1(G2090), .A2(n695), .ZN(n709) );
  NOR2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U781 ( .A1(n711), .A2(G303), .ZN(n712) );
  OR2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U783 ( .A(n717), .B(n716), .ZN(n725) );
  XNOR2_X1 U784 ( .A(n718), .B(KEYINPUT97), .ZN(n720) );
  NOR2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U786 ( .A1(G8), .A2(n721), .ZN(n722) );
  NAND2_X1 U787 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U788 ( .A1(n725), .A2(n724), .ZN(n771) );
  NOR2_X1 U789 ( .A1(G1976), .A2(G288), .ZN(n1016) );
  NOR2_X1 U790 ( .A1(G1971), .A2(G303), .ZN(n726) );
  NOR2_X1 U791 ( .A1(n1016), .A2(n726), .ZN(n727) );
  NAND2_X1 U792 ( .A1(n771), .A2(n727), .ZN(n728) );
  NAND2_X1 U793 ( .A1(G1976), .A2(G288), .ZN(n1017) );
  NOR2_X1 U794 ( .A1(n730), .A2(KEYINPUT33), .ZN(n731) );
  XNOR2_X1 U795 ( .A(n731), .B(KEYINPUT100), .ZN(n732) );
  XOR2_X1 U796 ( .A(G1981), .B(G305), .Z(n1010) );
  NOR2_X1 U797 ( .A1(n734), .A2(n733), .ZN(n795) );
  NAND2_X1 U798 ( .A1(n926), .A2(G128), .ZN(n737) );
  BUF_X1 U799 ( .A(n735), .Z(n928) );
  NAND2_X1 U800 ( .A1(G116), .A2(n928), .ZN(n736) );
  NAND2_X1 U801 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U802 ( .A(KEYINPUT35), .B(n738), .ZN(n745) );
  NAND2_X1 U803 ( .A1(G140), .A2(n739), .ZN(n741) );
  NAND2_X1 U804 ( .A1(G104), .A2(n932), .ZN(n740) );
  NAND2_X1 U805 ( .A1(n741), .A2(n740), .ZN(n743) );
  XOR2_X1 U806 ( .A(KEYINPUT86), .B(KEYINPUT34), .Z(n742) );
  XNOR2_X1 U807 ( .A(n743), .B(n742), .ZN(n744) );
  NAND2_X1 U808 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U809 ( .A(KEYINPUT36), .B(n746), .Z(n909) );
  XNOR2_X1 U810 ( .A(G2067), .B(KEYINPUT37), .ZN(n793) );
  OR2_X1 U811 ( .A1(n909), .A2(n793), .ZN(n747) );
  XNOR2_X1 U812 ( .A(n747), .B(KEYINPUT87), .ZN(n987) );
  NAND2_X1 U813 ( .A1(n795), .A2(n987), .ZN(n791) );
  NAND2_X1 U814 ( .A1(n926), .A2(G119), .ZN(n748) );
  XNOR2_X1 U815 ( .A(n748), .B(KEYINPUT88), .ZN(n750) );
  NAND2_X1 U816 ( .A1(G107), .A2(n928), .ZN(n749) );
  NAND2_X1 U817 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U818 ( .A(n751), .B(KEYINPUT89), .ZN(n753) );
  NAND2_X1 U819 ( .A1(G131), .A2(n739), .ZN(n752) );
  NAND2_X1 U820 ( .A1(n753), .A2(n752), .ZN(n756) );
  NAND2_X1 U821 ( .A1(n932), .A2(G95), .ZN(n754) );
  XOR2_X1 U822 ( .A(KEYINPUT90), .B(n754), .Z(n755) );
  NOR2_X1 U823 ( .A1(n756), .A2(n755), .ZN(n908) );
  INV_X1 U824 ( .A(G1991), .ZN(n954) );
  NOR2_X1 U825 ( .A1(n908), .A2(n954), .ZN(n765) );
  NAND2_X1 U826 ( .A1(G141), .A2(n739), .ZN(n758) );
  NAND2_X1 U827 ( .A1(G117), .A2(n928), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n758), .A2(n757), .ZN(n761) );
  NAND2_X1 U829 ( .A1(n932), .A2(G105), .ZN(n759) );
  XOR2_X1 U830 ( .A(KEYINPUT38), .B(n759), .Z(n760) );
  NOR2_X1 U831 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U832 ( .A1(n926), .A2(G129), .ZN(n762) );
  NAND2_X1 U833 ( .A1(n763), .A2(n762), .ZN(n916) );
  AND2_X1 U834 ( .A1(G1996), .A2(n916), .ZN(n764) );
  NOR2_X1 U835 ( .A1(n765), .A2(n764), .ZN(n985) );
  INV_X1 U836 ( .A(n985), .ZN(n766) );
  NAND2_X1 U837 ( .A1(n766), .A2(n795), .ZN(n784) );
  AND2_X1 U838 ( .A1(n791), .A2(n784), .ZN(n779) );
  AND2_X1 U839 ( .A1(n1010), .A2(n779), .ZN(n768) );
  NAND2_X1 U840 ( .A1(n1016), .A2(KEYINPUT33), .ZN(n767) );
  NOR2_X1 U841 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U842 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U843 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U844 ( .A1(n694), .A2(n772), .ZN(n773) );
  XOR2_X1 U845 ( .A(KEYINPUT101), .B(n773), .Z(n777) );
  NOR2_X1 U846 ( .A1(G1981), .A2(G305), .ZN(n774) );
  XOR2_X1 U847 ( .A(n774), .B(KEYINPUT24), .Z(n775) );
  OR2_X1 U848 ( .A1(n694), .A2(n775), .ZN(n776) );
  NAND2_X1 U849 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U850 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U851 ( .A(G1986), .B(G290), .ZN(n1024) );
  NAND2_X1 U852 ( .A1(n1024), .A2(n795), .ZN(n781) );
  NAND2_X1 U853 ( .A1(n782), .A2(n781), .ZN(n798) );
  NOR2_X1 U854 ( .A1(G1996), .A2(n916), .ZN(n783) );
  XOR2_X1 U855 ( .A(KEYINPUT103), .B(n783), .Z(n979) );
  INV_X1 U856 ( .A(n784), .ZN(n787) );
  NOR2_X1 U857 ( .A1(G1986), .A2(G290), .ZN(n785) );
  AND2_X1 U858 ( .A1(n954), .A2(n908), .ZN(n975) );
  NOR2_X1 U859 ( .A1(n785), .A2(n975), .ZN(n786) );
  NOR2_X1 U860 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U861 ( .A(n788), .B(KEYINPUT104), .ZN(n789) );
  NOR2_X1 U862 ( .A1(n979), .A2(n789), .ZN(n790) );
  XNOR2_X1 U863 ( .A(n790), .B(KEYINPUT39), .ZN(n792) );
  NAND2_X1 U864 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U865 ( .A1(n793), .A2(n909), .ZN(n989) );
  NAND2_X1 U866 ( .A1(n794), .A2(n989), .ZN(n796) );
  NAND2_X1 U867 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U868 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U869 ( .A(n799), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U870 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U871 ( .A1(G135), .A2(n739), .ZN(n801) );
  NAND2_X1 U872 ( .A1(G111), .A2(n928), .ZN(n800) );
  NAND2_X1 U873 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U874 ( .A1(n926), .A2(G123), .ZN(n802) );
  XOR2_X1 U875 ( .A(KEYINPUT18), .B(n802), .Z(n803) );
  NOR2_X1 U876 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U877 ( .A1(n932), .A2(G99), .ZN(n805) );
  NAND2_X1 U878 ( .A1(n806), .A2(n805), .ZN(n976) );
  XNOR2_X1 U879 ( .A(G2096), .B(n976), .ZN(n807) );
  OR2_X1 U880 ( .A1(G2100), .A2(n807), .ZN(G156) );
  INV_X1 U881 ( .A(G57), .ZN(G237) );
  INV_X1 U882 ( .A(G132), .ZN(G219) );
  INV_X1 U883 ( .A(G82), .ZN(G220) );
  NAND2_X1 U884 ( .A1(G7), .A2(G661), .ZN(n808) );
  XOR2_X1 U885 ( .A(n808), .B(KEYINPUT10), .Z(n863) );
  NAND2_X1 U886 ( .A1(n863), .A2(G567), .ZN(n809) );
  XOR2_X1 U887 ( .A(KEYINPUT11), .B(n809), .Z(G234) );
  NAND2_X1 U888 ( .A1(n1030), .A2(G860), .ZN(G153) );
  INV_X1 U889 ( .A(G868), .ZN(n846) );
  NAND2_X1 U890 ( .A1(n1027), .A2(n846), .ZN(n810) );
  XNOR2_X1 U891 ( .A(n810), .B(KEYINPUT74), .ZN(n812) );
  NAND2_X1 U892 ( .A1(G868), .A2(G301), .ZN(n811) );
  NAND2_X1 U893 ( .A1(n812), .A2(n811), .ZN(G284) );
  NOR2_X1 U894 ( .A1(G868), .A2(G299), .ZN(n813) );
  XNOR2_X1 U895 ( .A(n813), .B(KEYINPUT76), .ZN(n815) );
  NOR2_X1 U896 ( .A1(n846), .A2(G286), .ZN(n814) );
  NOR2_X1 U897 ( .A1(n815), .A2(n814), .ZN(G297) );
  INV_X1 U898 ( .A(G860), .ZN(n824) );
  NAND2_X1 U899 ( .A1(G559), .A2(n824), .ZN(n816) );
  XOR2_X1 U900 ( .A(KEYINPUT77), .B(n816), .Z(n817) );
  NAND2_X1 U901 ( .A1(n817), .A2(n942), .ZN(n818) );
  XNOR2_X1 U902 ( .A(n818), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U903 ( .A1(n1030), .A2(n846), .ZN(n819) );
  XOR2_X1 U904 ( .A(KEYINPUT78), .B(n819), .Z(n822) );
  NAND2_X1 U905 ( .A1(G868), .A2(n942), .ZN(n820) );
  NOR2_X1 U906 ( .A1(G559), .A2(n820), .ZN(n821) );
  NOR2_X1 U907 ( .A1(n822), .A2(n821), .ZN(G282) );
  NAND2_X1 U908 ( .A1(G559), .A2(n942), .ZN(n823) );
  XNOR2_X1 U909 ( .A(n823), .B(n1030), .ZN(n844) );
  NAND2_X1 U910 ( .A1(n824), .A2(n844), .ZN(n837) );
  NAND2_X1 U911 ( .A1(G55), .A2(n825), .ZN(n828) );
  NAND2_X1 U912 ( .A1(G67), .A2(n826), .ZN(n827) );
  NAND2_X1 U913 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U914 ( .A(KEYINPUT80), .B(n829), .ZN(n833) );
  NAND2_X1 U915 ( .A1(G80), .A2(n830), .ZN(n831) );
  XNOR2_X1 U916 ( .A(KEYINPUT79), .B(n831), .ZN(n832) );
  NOR2_X1 U917 ( .A1(n833), .A2(n832), .ZN(n836) );
  NAND2_X1 U918 ( .A1(n834), .A2(G93), .ZN(n835) );
  NAND2_X1 U919 ( .A1(n836), .A2(n835), .ZN(n847) );
  XNOR2_X1 U920 ( .A(n837), .B(n847), .ZN(G145) );
  XNOR2_X1 U921 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n839) );
  XOR2_X1 U922 ( .A(G288), .B(G303), .Z(n838) );
  XNOR2_X1 U923 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U924 ( .A(n840), .B(G305), .ZN(n841) );
  XNOR2_X1 U925 ( .A(n841), .B(n847), .ZN(n842) );
  XOR2_X1 U926 ( .A(G299), .B(n842), .Z(n843) );
  XNOR2_X1 U927 ( .A(n843), .B(G290), .ZN(n945) );
  XNOR2_X1 U928 ( .A(n844), .B(n945), .ZN(n845) );
  NOR2_X1 U929 ( .A1(n846), .A2(n845), .ZN(n849) );
  NOR2_X1 U930 ( .A1(G868), .A2(n847), .ZN(n848) );
  NOR2_X1 U931 ( .A1(n849), .A2(n848), .ZN(G295) );
  NAND2_X1 U932 ( .A1(G2084), .A2(G2078), .ZN(n850) );
  XOR2_X1 U933 ( .A(KEYINPUT20), .B(n850), .Z(n851) );
  NAND2_X1 U934 ( .A1(G2090), .A2(n851), .ZN(n852) );
  XNOR2_X1 U935 ( .A(KEYINPUT21), .B(n852), .ZN(n853) );
  NAND2_X1 U936 ( .A1(n853), .A2(G2072), .ZN(G158) );
  XOR2_X1 U937 ( .A(KEYINPUT85), .B(G44), .Z(n854) );
  XNOR2_X1 U938 ( .A(KEYINPUT3), .B(n854), .ZN(G218) );
  NOR2_X1 U939 ( .A1(G220), .A2(G219), .ZN(n855) );
  XOR2_X1 U940 ( .A(KEYINPUT22), .B(n855), .Z(n856) );
  NOR2_X1 U941 ( .A1(G218), .A2(n856), .ZN(n857) );
  NAND2_X1 U942 ( .A1(G96), .A2(n857), .ZN(n868) );
  NAND2_X1 U943 ( .A1(n868), .A2(G2106), .ZN(n861) );
  NAND2_X1 U944 ( .A1(G69), .A2(G120), .ZN(n858) );
  NOR2_X1 U945 ( .A1(G237), .A2(n858), .ZN(n859) );
  NAND2_X1 U946 ( .A1(G108), .A2(n859), .ZN(n867) );
  NAND2_X1 U947 ( .A1(n867), .A2(G567), .ZN(n860) );
  NAND2_X1 U948 ( .A1(n861), .A2(n860), .ZN(n880) );
  NAND2_X1 U949 ( .A1(G483), .A2(G661), .ZN(n862) );
  NOR2_X1 U950 ( .A1(n880), .A2(n862), .ZN(n866) );
  NAND2_X1 U951 ( .A1(n866), .A2(G36), .ZN(G176) );
  NAND2_X1 U952 ( .A1(G2106), .A2(n863), .ZN(G217) );
  INV_X1 U953 ( .A(n863), .ZN(G223) );
  AND2_X1 U954 ( .A1(G15), .A2(G2), .ZN(n864) );
  NAND2_X1 U955 ( .A1(G661), .A2(n864), .ZN(G259) );
  NAND2_X1 U956 ( .A1(G3), .A2(G1), .ZN(n865) );
  NAND2_X1 U957 ( .A1(n866), .A2(n865), .ZN(G188) );
  INV_X1 U959 ( .A(G120), .ZN(G236) );
  INV_X1 U960 ( .A(G96), .ZN(G221) );
  INV_X1 U961 ( .A(G69), .ZN(G235) );
  NOR2_X1 U962 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U963 ( .A(n869), .B(KEYINPUT107), .Z(G325) );
  INV_X1 U964 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U965 ( .A(G1341), .B(G2454), .ZN(n870) );
  XNOR2_X1 U966 ( .A(n870), .B(G2430), .ZN(n871) );
  XNOR2_X1 U967 ( .A(n871), .B(G1348), .ZN(n877) );
  XOR2_X1 U968 ( .A(G2443), .B(G2427), .Z(n873) );
  XNOR2_X1 U969 ( .A(G2438), .B(G2446), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n875) );
  XOR2_X1 U971 ( .A(G2451), .B(G2435), .Z(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U973 ( .A(n877), .B(n876), .ZN(n878) );
  NAND2_X1 U974 ( .A1(n878), .A2(G14), .ZN(n879) );
  XNOR2_X1 U975 ( .A(KEYINPUT105), .B(n879), .ZN(n951) );
  XNOR2_X1 U976 ( .A(n951), .B(KEYINPUT106), .ZN(G401) );
  INV_X1 U977 ( .A(n880), .ZN(G319) );
  XOR2_X1 U978 ( .A(G2096), .B(KEYINPUT43), .Z(n882) );
  XNOR2_X1 U979 ( .A(G2090), .B(G2678), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U981 ( .A(n883), .B(KEYINPUT108), .Z(n885) );
  XNOR2_X1 U982 ( .A(G2067), .B(G2072), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U984 ( .A(KEYINPUT42), .B(G2100), .Z(n887) );
  XNOR2_X1 U985 ( .A(G2084), .B(G2078), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(G227) );
  XNOR2_X1 U988 ( .A(n890), .B(G1971), .ZN(n892) );
  XNOR2_X1 U989 ( .A(G1986), .B(G1976), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U991 ( .A(n893), .B(G2474), .Z(n895) );
  XNOR2_X1 U992 ( .A(G1981), .B(G1966), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U994 ( .A(KEYINPUT41), .B(G1961), .Z(n897) );
  XOR2_X1 U995 ( .A(G1996), .B(n954), .Z(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(G229) );
  NAND2_X1 U998 ( .A1(n928), .A2(G112), .ZN(n906) );
  NAND2_X1 U999 ( .A1(G136), .A2(n739), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(G100), .A2(n932), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(n926), .A2(G124), .ZN(n902) );
  XOR2_X1 U1003 ( .A(KEYINPUT44), .B(n902), .Z(n903) );
  NOR2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n907), .B(KEYINPUT109), .ZN(G162) );
  XOR2_X1 U1007 ( .A(G162), .B(n908), .Z(n911) );
  XOR2_X1 U1008 ( .A(G160), .B(n909), .Z(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n976), .B(KEYINPUT46), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1013 ( .A(n915), .B(n914), .Z(n918) );
  XOR2_X1 U1014 ( .A(G164), .B(n916), .Z(n917) );
  XNOR2_X1 U1015 ( .A(n918), .B(n917), .ZN(n940) );
  NAND2_X1 U1016 ( .A1(G139), .A2(n739), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(G103), .A2(n932), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n925) );
  NAND2_X1 U1019 ( .A1(n926), .A2(G127), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(G115), .A2(n928), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT47), .B(n923), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n992) );
  NAND2_X1 U1024 ( .A1(G130), .A2(n926), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n927), .B(KEYINPUT110), .ZN(n931) );
  NAND2_X1 U1026 ( .A1(n928), .A2(G118), .ZN(n929) );
  XOR2_X1 U1027 ( .A(KEYINPUT111), .B(n929), .Z(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(G142), .A2(n739), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(G106), .A2(n932), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT45), .B(n935), .Z(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(n992), .B(n938), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(n940), .B(n939), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(G37), .A2(n941), .ZN(G395) );
  XOR2_X1 U1037 ( .A(G286), .B(n1030), .Z(n944) );
  XOR2_X1 U1038 ( .A(G301), .B(n942), .Z(n943) );
  XNOR2_X1 U1039 ( .A(n944), .B(n943), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(n946), .B(n945), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(G37), .A2(n947), .ZN(G397) );
  NOR2_X1 U1042 ( .A1(G227), .A2(G229), .ZN(n948) );
  XOR2_X1 U1043 ( .A(KEYINPUT49), .B(n948), .Z(n949) );
  NAND2_X1 U1044 ( .A1(G319), .A2(n949), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n953) );
  NOR2_X1 U1046 ( .A1(G395), .A2(G397), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(G225) );
  INV_X1 U1048 ( .A(G225), .ZN(G308) );
  INV_X1 U1049 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1050 ( .A(n954), .B(G25), .Z(n965) );
  XOR2_X1 U1051 ( .A(G32), .B(G1996), .Z(n959) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(G27), .B(n955), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT116), .B(G2072), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(G33), .B(n960), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(KEYINPUT117), .B(n963), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(G28), .A2(n966), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n967), .B(KEYINPUT53), .ZN(n970) );
  XOR2_X1 U1063 ( .A(G2084), .B(G34), .Z(n968) );
  XNOR2_X1 U1064 ( .A(KEYINPUT54), .B(n968), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G35), .B(G2090), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n1002) );
  NAND2_X1 U1068 ( .A1(KEYINPUT55), .A2(n1002), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(G11), .A2(n973), .ZN(n1008) );
  XOR2_X1 U1070 ( .A(G160), .B(G2084), .Z(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n983) );
  XOR2_X1 U1073 ( .A(G2090), .B(G162), .Z(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1075 ( .A(KEYINPUT113), .B(n980), .Z(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT51), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(n988), .B(KEYINPUT114), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1082 ( .A(KEYINPUT115), .B(n991), .Z(n997) );
  XOR2_X1 U1083 ( .A(G2072), .B(n992), .Z(n994) );
  XOR2_X1 U1084 ( .A(G164), .B(G2078), .Z(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1086 ( .A(KEYINPUT50), .B(n995), .Z(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(KEYINPUT52), .B(n998), .ZN(n1000) );
  INV_X1 U1089 ( .A(KEYINPUT55), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(G29), .ZN(n1006) );
  INV_X1 U1092 ( .A(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1067) );
  XOR2_X1 U1097 ( .A(G16), .B(KEYINPUT56), .Z(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT118), .B(n1009), .ZN(n1037) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G168), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1012), .B(KEYINPUT57), .ZN(n1026) );
  XOR2_X1 U1102 ( .A(G1971), .B(G303), .Z(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT120), .B(n1013), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(G299), .B(G1956), .Z(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1021) );
  INV_X1 U1106 ( .A(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(KEYINPUT119), .B(n1019), .Z(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(n1022), .B(KEYINPUT121), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1035) );
  XNOR2_X1 U1113 ( .A(G1348), .B(n1027), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(G301), .B(G1961), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(n1030), .B(G1341), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(n1031), .B(KEYINPUT122), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1120 ( .A1(n1037), .A2(n1036), .ZN(n1064) );
  XOR2_X1 U1121 ( .A(G20), .B(G1956), .Z(n1041) );
  XNOR2_X1 U1122 ( .A(G1981), .B(G6), .ZN(n1039) );
  XNOR2_X1 U1123 ( .A(G19), .B(G1341), .ZN(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1044) );
  XOR2_X1 U1126 ( .A(KEYINPUT59), .B(G1348), .Z(n1042) );
  XNOR2_X1 U1127 ( .A(G4), .B(n1042), .ZN(n1043) );
  NOR2_X1 U1128 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1129 ( .A(KEYINPUT60), .B(n1045), .ZN(n1046) );
  XNOR2_X1 U1130 ( .A(n1046), .B(KEYINPUT124), .ZN(n1050) );
  XNOR2_X1 U1131 ( .A(G1966), .B(G21), .ZN(n1048) );
  XNOR2_X1 U1132 ( .A(G5), .B(G1961), .ZN(n1047) );
  NOR2_X1 U1133 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NAND2_X1 U1134 ( .A1(n1050), .A2(n1049), .ZN(n1059) );
  XNOR2_X1 U1135 ( .A(G1986), .B(G24), .ZN(n1055) );
  XNOR2_X1 U1136 ( .A(G1976), .B(G23), .ZN(n1052) );
  XNOR2_X1 U1137 ( .A(G1971), .B(G22), .ZN(n1051) );
  NOR2_X1 U1138 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  XNOR2_X1 U1139 ( .A(KEYINPUT125), .B(n1053), .ZN(n1054) );
  NOR2_X1 U1140 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  XOR2_X1 U1141 ( .A(KEYINPUT126), .B(n1056), .Z(n1057) );
  XNOR2_X1 U1142 ( .A(KEYINPUT58), .B(n1057), .ZN(n1058) );
  NOR2_X1 U1143 ( .A1(n1059), .A2(n1058), .ZN(n1060) );
  XOR2_X1 U1144 ( .A(KEYINPUT61), .B(n1060), .Z(n1062) );
  XOR2_X1 U1145 ( .A(G16), .B(KEYINPUT123), .Z(n1061) );
  NOR2_X1 U1146 ( .A1(n1062), .A2(n1061), .ZN(n1063) );
  NOR2_X1 U1147 ( .A1(n1064), .A2(n1063), .ZN(n1065) );
  XOR2_X1 U1148 ( .A(KEYINPUT127), .B(n1065), .Z(n1066) );
  NAND2_X1 U1149 ( .A1(n1067), .A2(n1066), .ZN(n1068) );
  XNOR2_X1 U1150 ( .A(KEYINPUT62), .B(n1068), .ZN(G150) );
  INV_X1 U1151 ( .A(G150), .ZN(G311) );
endmodule

