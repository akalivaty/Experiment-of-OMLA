

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U550 ( .A(n599), .Z(G164) );
  NOR2_X1 U551 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U552 ( .A1(n656), .A2(n655), .ZN(n669) );
  NOR2_X1 U553 ( .A1(G168), .A2(n661), .ZN(n662) );
  NOR2_X1 U554 ( .A1(n658), .A2(n684), .ZN(n660) );
  NOR2_X1 U555 ( .A1(n709), .A2(G1966), .ZN(n657) );
  XNOR2_X1 U556 ( .A(n621), .B(KEYINPUT26), .ZN(n623) );
  AND2_X1 U557 ( .A1(n516), .A2(n536), .ZN(n599) );
  AND2_X1 U558 ( .A1(n534), .A2(n519), .ZN(n516) );
  XNOR2_X1 U559 ( .A(n718), .B(n517), .ZN(n530) );
  INV_X1 U560 ( .A(KEYINPUT17), .ZN(n517) );
  NAND2_X1 U561 ( .A1(n530), .A2(G138), .ZN(n531) );
  NAND2_X1 U562 ( .A1(n632), .A2(n978), .ZN(n631) );
  NOR2_X1 U563 ( .A1(n624), .A2(n769), .ZN(n632) );
  NOR2_X2 U564 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X4 U565 ( .A1(G2104), .A2(G2105), .ZN(n718) );
  BUF_X2 U566 ( .A(n625), .Z(n627) );
  AND2_X2 U567 ( .A1(n524), .A2(G2104), .ZN(n888) );
  AND2_X2 U568 ( .A1(n526), .A2(G2105), .ZN(n885) );
  XOR2_X1 U569 ( .A(G543), .B(KEYINPUT0), .Z(n555) );
  INV_X1 U570 ( .A(G651), .ZN(n541) );
  INV_X1 U571 ( .A(G2105), .ZN(n524) );
  NOR2_X1 U572 ( .A1(n555), .A2(n541), .ZN(n538) );
  AND2_X1 U573 ( .A1(G125), .A2(n885), .ZN(n518) );
  AND2_X1 U574 ( .A1(n533), .A2(n532), .ZN(n519) );
  INV_X1 U575 ( .A(KEYINPUT30), .ZN(n659) );
  XNOR2_X1 U576 ( .A(KEYINPUT29), .B(KEYINPUT104), .ZN(n649) );
  INV_X1 U577 ( .A(KEYINPUT31), .ZN(n666) );
  XNOR2_X1 U578 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U579 ( .A1(n600), .A2(n735), .ZN(n625) );
  NAND2_X2 U580 ( .A1(G8), .A2(n627), .ZN(n709) );
  INV_X1 U581 ( .A(G2104), .ZN(n526) );
  NOR2_X1 U582 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U583 ( .A(n617), .B(KEYINPUT71), .ZN(n619) );
  XNOR2_X1 U584 ( .A(n543), .B(n542), .ZN(n792) );
  NAND2_X1 U585 ( .A1(n619), .A2(n618), .ZN(n769) );
  BUF_X1 U586 ( .A(n769), .Z(n992) );
  AND2_X1 U587 ( .A1(n529), .A2(n528), .ZN(G160) );
  NAND2_X1 U588 ( .A1(n530), .A2(G137), .ZN(n522) );
  AND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U590 ( .A1(G113), .A2(n884), .ZN(n521) );
  NAND2_X1 U591 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n523), .B(KEYINPUT65), .ZN(n529) );
  NAND2_X1 U593 ( .A1(G101), .A2(n888), .ZN(n525) );
  XNOR2_X1 U594 ( .A(KEYINPUT23), .B(n525), .ZN(n527) );
  NOR2_X1 U595 ( .A1(n527), .A2(n518), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT88), .ZN(n534) );
  NAND2_X1 U597 ( .A1(G114), .A2(n884), .ZN(n533) );
  NAND2_X1 U598 ( .A1(G102), .A2(n888), .ZN(n532) );
  NAND2_X1 U599 ( .A1(G126), .A2(n885), .ZN(n535) );
  XOR2_X1 U600 ( .A(KEYINPUT87), .B(n535), .Z(n536) );
  XOR2_X1 U601 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n540) );
  XNOR2_X2 U602 ( .A(n538), .B(KEYINPUT66), .ZN(n796) );
  NAND2_X1 U603 ( .A1(G73), .A2(n796), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n547) );
  NOR2_X1 U605 ( .A1(G543), .A2(n541), .ZN(n543) );
  XNOR2_X1 U606 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n542) );
  NAND2_X1 U607 ( .A1(G61), .A2(n792), .ZN(n545) );
  NOR2_X1 U608 ( .A1(G651), .A2(G543), .ZN(n793) );
  NAND2_X1 U609 ( .A1(G86), .A2(n793), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n550) );
  NOR2_X1 U612 ( .A1(G651), .A2(n555), .ZN(n548) );
  XNOR2_X2 U613 ( .A(KEYINPUT64), .B(n548), .ZN(n797) );
  NAND2_X1 U614 ( .A1(G48), .A2(n797), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(G305) );
  NAND2_X1 U616 ( .A1(G651), .A2(G74), .ZN(n552) );
  NAND2_X1 U617 ( .A1(G49), .A2(n797), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U619 ( .A1(n792), .A2(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(KEYINPUT78), .ZN(n557) );
  NAND2_X1 U621 ( .A1(G87), .A2(n555), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT79), .B(n558), .Z(G288) );
  NAND2_X1 U624 ( .A1(G65), .A2(n792), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G91), .A2(n793), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G78), .A2(n796), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G53), .A2(n797), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  OR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(G299) );
  NAND2_X1 U631 ( .A1(G64), .A2(n792), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G52), .A2(n797), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G77), .A2(n796), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT68), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G90), .A2(n793), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U639 ( .A1(n572), .A2(n571), .ZN(G171) );
  INV_X1 U640 ( .A(G171), .ZN(G301) );
  NAND2_X1 U641 ( .A1(G63), .A2(n792), .ZN(n574) );
  NAND2_X1 U642 ( .A1(G51), .A2(n797), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U644 ( .A(KEYINPUT6), .B(n575), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n793), .A2(G89), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n576), .B(KEYINPUT4), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G76), .A2(n796), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U649 ( .A(KEYINPUT5), .B(n579), .Z(n580) );
  XNOR2_X1 U650 ( .A(KEYINPUT72), .B(n580), .ZN(n581) );
  NOR2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U652 ( .A(KEYINPUT7), .B(n583), .Z(G168) );
  XOR2_X1 U653 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U654 ( .A1(G75), .A2(n796), .ZN(n584) );
  XOR2_X1 U655 ( .A(KEYINPUT81), .B(n584), .Z(n586) );
  NAND2_X1 U656 ( .A1(n793), .A2(G88), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U658 ( .A(KEYINPUT82), .B(n587), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G62), .A2(n792), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G50), .A2(n797), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U662 ( .A1(n591), .A2(n590), .ZN(G166) );
  INV_X1 U663 ( .A(G166), .ZN(G303) );
  AND2_X1 U664 ( .A1(n793), .A2(G85), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G60), .A2(n792), .ZN(n593) );
  NAND2_X1 U666 ( .A1(G47), .A2(n797), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G72), .A2(n796), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(G290) );
  XOR2_X1 U671 ( .A(G1981), .B(G305), .Z(n975) );
  NAND2_X1 U672 ( .A1(G160), .A2(G40), .ZN(n734) );
  INV_X1 U673 ( .A(n734), .ZN(n600) );
  NOR2_X1 U674 ( .A1(n599), .A2(G1384), .ZN(n735) );
  NOR2_X1 U675 ( .A1(G1976), .A2(G288), .ZN(n690) );
  NAND2_X1 U676 ( .A1(n690), .A2(KEYINPUT33), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n709), .A2(n601), .ZN(n699) );
  NAND2_X1 U678 ( .A1(G66), .A2(n792), .ZN(n603) );
  NAND2_X1 U679 ( .A1(G92), .A2(n793), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G79), .A2(n796), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G54), .A2(n797), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X2 U685 ( .A(KEYINPUT15), .B(n608), .Z(n978) );
  NAND2_X1 U686 ( .A1(n792), .A2(G56), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n609), .B(KEYINPUT14), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n796), .A2(G68), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n793), .A2(G81), .ZN(n610) );
  XNOR2_X1 U690 ( .A(n610), .B(KEYINPUT12), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n614) );
  XNOR2_X1 U692 ( .A(KEYINPUT70), .B(KEYINPUT13), .ZN(n613) );
  XNOR2_X1 U693 ( .A(n614), .B(n613), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G43), .A2(n797), .ZN(n618) );
  INV_X1 U696 ( .A(n625), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n620), .A2(G1996), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n627), .A2(G1341), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  INV_X1 U700 ( .A(n625), .ZN(n637) );
  AND2_X1 U701 ( .A1(n637), .A2(G2067), .ZN(n626) );
  XNOR2_X1 U702 ( .A(n626), .B(KEYINPUT101), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n627), .A2(G1348), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n634) );
  OR2_X1 U706 ( .A1(n978), .A2(n632), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n636) );
  INV_X1 U708 ( .A(KEYINPUT102), .ZN(n635) );
  XNOR2_X1 U709 ( .A(n636), .B(n635), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n627), .A2(G1956), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n637), .A2(G2072), .ZN(n638) );
  XOR2_X1 U712 ( .A(KEYINPUT27), .B(n638), .Z(n639) );
  NAND2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n641), .B(KEYINPUT100), .ZN(n645) );
  NOR2_X1 U715 ( .A1(n645), .A2(G299), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n644), .B(KEYINPUT103), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n645), .A2(G299), .ZN(n646) );
  XNOR2_X1 U718 ( .A(KEYINPUT28), .B(n646), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n650), .B(n649), .ZN(n656) );
  XOR2_X1 U721 ( .A(KEYINPUT25), .B(G2078), .Z(n960) );
  NOR2_X1 U722 ( .A1(n960), .A2(n627), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n651), .B(KEYINPUT98), .ZN(n653) );
  NOR2_X1 U724 ( .A1(n637), .A2(G1961), .ZN(n652) );
  NOR2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U726 ( .A(KEYINPUT99), .B(n654), .Z(n663) );
  NOR2_X1 U727 ( .A1(G301), .A2(n663), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n657), .B(KEYINPUT97), .ZN(n681) );
  NAND2_X1 U729 ( .A1(G8), .A2(n681), .ZN(n658) );
  NOR2_X1 U730 ( .A1(G2084), .A2(n627), .ZN(n684) );
  XNOR2_X1 U731 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n662), .B(KEYINPUT105), .ZN(n665) );
  NAND2_X1 U733 ( .A1(n663), .A2(G301), .ZN(n664) );
  NAND2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n671) );
  INV_X1 U736 ( .A(KEYINPUT106), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n671), .B(n670), .ZN(n682) );
  AND2_X1 U738 ( .A1(G286), .A2(G8), .ZN(n672) );
  AND2_X1 U739 ( .A1(n682), .A2(n672), .ZN(n679) );
  INV_X1 U740 ( .A(G8), .ZN(n677) );
  NOR2_X1 U741 ( .A1(G1971), .A2(n709), .ZN(n674) );
  NOR2_X1 U742 ( .A1(G2090), .A2(n627), .ZN(n673) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n675), .A2(G303), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n680), .B(KEYINPUT32), .ZN(n688) );
  NAND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n683), .B(KEYINPUT107), .ZN(n686) );
  NAND2_X1 U749 ( .A1(n684), .A2(G8), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n703) );
  NOR2_X1 U752 ( .A1(G1971), .A2(G303), .ZN(n689) );
  NOR2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n985) );
  INV_X1 U754 ( .A(KEYINPUT33), .ZN(n691) );
  AND2_X1 U755 ( .A1(n985), .A2(n691), .ZN(n692) );
  NAND2_X1 U756 ( .A1(n703), .A2(n692), .ZN(n697) );
  INV_X1 U757 ( .A(n709), .ZN(n694) );
  NAND2_X1 U758 ( .A1(G288), .A2(G1976), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n693), .B(KEYINPUT108), .ZN(n986) );
  AND2_X1 U760 ( .A1(n694), .A2(n986), .ZN(n695) );
  OR2_X1 U761 ( .A1(KEYINPUT33), .A2(n695), .ZN(n696) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n700) );
  AND2_X1 U764 ( .A1(n975), .A2(n700), .ZN(n715) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n701) );
  NAND2_X1 U766 ( .A1(G8), .A2(n701), .ZN(n702) );
  NAND2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n705) );
  INV_X1 U768 ( .A(KEYINPUT109), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n705), .B(n704), .ZN(n706) );
  NAND2_X1 U770 ( .A1(n706), .A2(n709), .ZN(n713) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n707), .B(KEYINPUT24), .ZN(n708) );
  XNOR2_X1 U773 ( .A(n708), .B(KEYINPUT95), .ZN(n710) );
  NOR2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U775 ( .A(n711), .B(KEYINPUT96), .Z(n712) );
  NAND2_X1 U776 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U777 ( .A1(n715), .A2(n714), .ZN(n749) );
  NAND2_X1 U778 ( .A1(G95), .A2(n888), .ZN(n717) );
  NAND2_X1 U779 ( .A1(G119), .A2(n885), .ZN(n716) );
  NAND2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n721) );
  XOR2_X1 U781 ( .A(n718), .B(KEYINPUT17), .Z(n889) );
  NAND2_X1 U782 ( .A1(n889), .A2(G131), .ZN(n719) );
  XOR2_X1 U783 ( .A(KEYINPUT90), .B(n719), .Z(n720) );
  NOR2_X1 U784 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U785 ( .A1(n884), .A2(G107), .ZN(n722) );
  NAND2_X1 U786 ( .A1(n723), .A2(n722), .ZN(n897) );
  XOR2_X1 U787 ( .A(KEYINPUT91), .B(G1991), .Z(n951) );
  AND2_X1 U788 ( .A1(n897), .A2(n951), .ZN(n724) );
  XNOR2_X1 U789 ( .A(n724), .B(KEYINPUT92), .ZN(n733) );
  NAND2_X1 U790 ( .A1(G117), .A2(n884), .ZN(n726) );
  NAND2_X1 U791 ( .A1(G129), .A2(n885), .ZN(n725) );
  NAND2_X1 U792 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U793 ( .A1(n888), .A2(G105), .ZN(n727) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n727), .Z(n728) );
  NOR2_X1 U795 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U796 ( .A1(n889), .A2(G141), .ZN(n730) );
  NAND2_X1 U797 ( .A1(n731), .A2(n730), .ZN(n880) );
  AND2_X1 U798 ( .A1(G1996), .A2(n880), .ZN(n732) );
  NOR2_X1 U799 ( .A1(n733), .A2(n732), .ZN(n936) );
  NOR2_X1 U800 ( .A1(n735), .A2(n734), .ZN(n762) );
  XNOR2_X1 U801 ( .A(KEYINPUT93), .B(n762), .ZN(n736) );
  NOR2_X1 U802 ( .A1(n936), .A2(n736), .ZN(n755) );
  XOR2_X1 U803 ( .A(KEYINPUT94), .B(n755), .Z(n747) );
  XNOR2_X1 U804 ( .A(G2067), .B(KEYINPUT37), .ZN(n760) );
  NAND2_X1 U805 ( .A1(G104), .A2(n888), .ZN(n738) );
  NAND2_X1 U806 ( .A1(G140), .A2(n889), .ZN(n737) );
  NAND2_X1 U807 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U808 ( .A(KEYINPUT34), .B(n739), .ZN(n745) );
  NAND2_X1 U809 ( .A1(n885), .A2(G128), .ZN(n740) );
  XOR2_X1 U810 ( .A(KEYINPUT89), .B(n740), .Z(n742) );
  NAND2_X1 U811 ( .A1(n884), .A2(G116), .ZN(n741) );
  NAND2_X1 U812 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U813 ( .A(KEYINPUT35), .B(n743), .Z(n744) );
  NOR2_X1 U814 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U815 ( .A(KEYINPUT36), .B(n746), .ZN(n881) );
  NOR2_X1 U816 ( .A1(n760), .A2(n881), .ZN(n934) );
  NAND2_X1 U817 ( .A1(n762), .A2(n934), .ZN(n758) );
  NAND2_X1 U818 ( .A1(n747), .A2(n758), .ZN(n748) );
  XNOR2_X1 U819 ( .A(n750), .B(KEYINPUT110), .ZN(n752) );
  XNOR2_X1 U820 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U821 ( .A1(n984), .A2(n762), .ZN(n751) );
  NAND2_X1 U822 ( .A1(n752), .A2(n751), .ZN(n765) );
  NOR2_X1 U823 ( .A1(G1996), .A2(n880), .ZN(n925) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n753) );
  NOR2_X1 U825 ( .A1(n951), .A2(n897), .ZN(n930) );
  NOR2_X1 U826 ( .A1(n753), .A2(n930), .ZN(n754) );
  NOR2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U828 ( .A1(n925), .A2(n756), .ZN(n757) );
  XNOR2_X1 U829 ( .A(KEYINPUT39), .B(n757), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U831 ( .A1(n760), .A2(n881), .ZN(n938) );
  NAND2_X1 U832 ( .A1(n761), .A2(n938), .ZN(n763) );
  NAND2_X1 U833 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U834 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U835 ( .A(n766), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U836 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U837 ( .A(G132), .ZN(G219) );
  INV_X1 U838 ( .A(G82), .ZN(G220) );
  NAND2_X1 U839 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U840 ( .A(n767), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U841 ( .A(G223), .ZN(n829) );
  NAND2_X1 U842 ( .A1(n829), .A2(G567), .ZN(n768) );
  XOR2_X1 U843 ( .A(KEYINPUT11), .B(n768), .Z(G234) );
  INV_X1 U844 ( .A(G860), .ZN(n838) );
  OR2_X1 U845 ( .A1(n992), .A2(n838), .ZN(G153) );
  NAND2_X1 U846 ( .A1(G868), .A2(G301), .ZN(n771) );
  OR2_X1 U847 ( .A1(n978), .A2(G868), .ZN(n770) );
  NAND2_X1 U848 ( .A1(n771), .A2(n770), .ZN(G284) );
  INV_X1 U849 ( .A(G868), .ZN(n810) );
  NOR2_X1 U850 ( .A1(G286), .A2(n810), .ZN(n772) );
  XOR2_X1 U851 ( .A(KEYINPUT73), .B(n772), .Z(n774) );
  NOR2_X1 U852 ( .A1(G868), .A2(G299), .ZN(n773) );
  NOR2_X1 U853 ( .A1(n774), .A2(n773), .ZN(G297) );
  NAND2_X1 U854 ( .A1(n838), .A2(G559), .ZN(n775) );
  NAND2_X1 U855 ( .A1(n775), .A2(n978), .ZN(n776) );
  XNOR2_X1 U856 ( .A(n776), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U857 ( .A1(G868), .A2(n992), .ZN(n779) );
  NAND2_X1 U858 ( .A1(G868), .A2(n978), .ZN(n777) );
  NOR2_X1 U859 ( .A1(G559), .A2(n777), .ZN(n778) );
  NOR2_X1 U860 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U861 ( .A1(G111), .A2(n884), .ZN(n781) );
  NAND2_X1 U862 ( .A1(G99), .A2(n888), .ZN(n780) );
  NAND2_X1 U863 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U864 ( .A(KEYINPUT74), .B(n782), .ZN(n785) );
  NAND2_X1 U865 ( .A1(n885), .A2(G123), .ZN(n783) );
  XOR2_X1 U866 ( .A(KEYINPUT18), .B(n783), .Z(n784) );
  NOR2_X1 U867 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U868 ( .A1(n889), .A2(G135), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n787), .A2(n786), .ZN(n927) );
  XOR2_X1 U870 ( .A(n927), .B(G2096), .Z(n789) );
  XNOR2_X1 U871 ( .A(G2100), .B(KEYINPUT75), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n789), .A2(n788), .ZN(G156) );
  NAND2_X1 U873 ( .A1(G559), .A2(n978), .ZN(n790) );
  XOR2_X1 U874 ( .A(KEYINPUT76), .B(n790), .Z(n791) );
  XNOR2_X1 U875 ( .A(n992), .B(n791), .ZN(n837) );
  XNOR2_X1 U876 ( .A(G166), .B(G288), .ZN(n808) );
  NAND2_X1 U877 ( .A1(G67), .A2(n792), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G93), .A2(n793), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n801) );
  NAND2_X1 U880 ( .A1(G80), .A2(n796), .ZN(n799) );
  NAND2_X1 U881 ( .A1(G55), .A2(n797), .ZN(n798) );
  NAND2_X1 U882 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U883 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U884 ( .A(KEYINPUT77), .B(n802), .ZN(n839) );
  XOR2_X1 U885 ( .A(KEYINPUT83), .B(n839), .Z(n804) );
  XNOR2_X1 U886 ( .A(G299), .B(KEYINPUT19), .ZN(n803) );
  XNOR2_X1 U887 ( .A(n804), .B(n803), .ZN(n805) );
  XOR2_X1 U888 ( .A(n805), .B(G290), .Z(n806) );
  XNOR2_X1 U889 ( .A(G305), .B(n806), .ZN(n807) );
  XNOR2_X1 U890 ( .A(n808), .B(n807), .ZN(n902) );
  XNOR2_X1 U891 ( .A(n837), .B(n902), .ZN(n809) );
  NAND2_X1 U892 ( .A1(n809), .A2(G868), .ZN(n812) );
  NAND2_X1 U893 ( .A1(n810), .A2(n839), .ZN(n811) );
  NAND2_X1 U894 ( .A1(n812), .A2(n811), .ZN(G295) );
  XOR2_X1 U895 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n814) );
  NAND2_X1 U896 ( .A1(G2078), .A2(G2084), .ZN(n813) );
  XNOR2_X1 U897 ( .A(n814), .B(n813), .ZN(n815) );
  NAND2_X1 U898 ( .A1(n815), .A2(G2090), .ZN(n816) );
  XOR2_X1 U899 ( .A(KEYINPUT85), .B(n816), .Z(n817) );
  XNOR2_X1 U900 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U901 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U902 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U903 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U904 ( .A1(G120), .A2(G108), .ZN(n819) );
  NOR2_X1 U905 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U906 ( .A1(G69), .A2(n820), .ZN(n835) );
  NAND2_X1 U907 ( .A1(G567), .A2(n835), .ZN(n825) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n821) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n821), .Z(n822) );
  NOR2_X1 U910 ( .A1(G218), .A2(n822), .ZN(n823) );
  NAND2_X1 U911 ( .A1(G96), .A2(n823), .ZN(n836) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n836), .ZN(n824) );
  NAND2_X1 U913 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U914 ( .A(KEYINPUT86), .B(n826), .Z(G319) );
  INV_X1 U915 ( .A(G319), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G661), .A2(G483), .ZN(n827) );
  NOR2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n834) );
  NAND2_X1 U918 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n829), .ZN(G217) );
  NAND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n831) );
  INV_X1 U921 ( .A(G661), .ZN(n830) );
  NOR2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U923 ( .A(n832), .B(KEYINPUT113), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U925 ( .A1(n834), .A2(n833), .ZN(G188) );
  XOR2_X1 U926 ( .A(G96), .B(KEYINPUT114), .Z(G221) );
  XOR2_X1 U927 ( .A(G108), .B(KEYINPUT120), .Z(G238) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  NAND2_X1 U933 ( .A1(n838), .A2(n837), .ZN(n840) );
  XNOR2_X1 U934 ( .A(n840), .B(n839), .ZN(G145) );
  XOR2_X1 U935 ( .A(KEYINPUT42), .B(G2090), .Z(n842) );
  XNOR2_X1 U936 ( .A(G2084), .B(G2072), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U938 ( .A(n843), .B(G2100), .Z(n845) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2078), .ZN(n844) );
  XNOR2_X1 U940 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U942 ( .A(G2678), .B(KEYINPUT115), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U944 ( .A(n849), .B(n848), .Z(G227) );
  XNOR2_X1 U945 ( .A(G1961), .B(G2474), .ZN(n859) );
  XOR2_X1 U946 ( .A(G1966), .B(G1976), .Z(n851) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1981), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U949 ( .A(G1956), .B(G1971), .Z(n853) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U953 ( .A(KEYINPUT116), .B(KEYINPUT41), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G124), .A2(n885), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U958 ( .A1(n884), .A2(G112), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U960 ( .A1(G100), .A2(n888), .ZN(n864) );
  NAND2_X1 U961 ( .A1(G136), .A2(n889), .ZN(n863) );
  NAND2_X1 U962 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U963 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U964 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n868) );
  XNOR2_X1 U965 ( .A(G164), .B(KEYINPUT48), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n879) );
  NAND2_X1 U967 ( .A1(G103), .A2(n888), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G139), .A2(n889), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G115), .A2(n884), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G127), .A2(n885), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT47), .B(n873), .ZN(n874) );
  XNOR2_X1 U974 ( .A(KEYINPUT117), .B(n874), .ZN(n875) );
  NOR2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n940) );
  XNOR2_X1 U976 ( .A(G160), .B(n940), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(G162), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n883) );
  XOR2_X1 U979 ( .A(n881), .B(n880), .Z(n882) );
  XNOR2_X1 U980 ( .A(n883), .B(n882), .ZN(n899) );
  NAND2_X1 U981 ( .A1(G118), .A2(n884), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G130), .A2(n885), .ZN(n886) );
  NAND2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n894) );
  NAND2_X1 U984 ( .A1(G106), .A2(n888), .ZN(n891) );
  NAND2_X1 U985 ( .A1(G142), .A2(n889), .ZN(n890) );
  NAND2_X1 U986 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U987 ( .A(n892), .B(KEYINPUT45), .Z(n893) );
  NOR2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n895), .B(n927), .ZN(n896) );
  XOR2_X1 U990 ( .A(n897), .B(n896), .Z(n898) );
  XNOR2_X1 U991 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U992 ( .A1(G37), .A2(n900), .ZN(n901) );
  XOR2_X1 U993 ( .A(KEYINPUT119), .B(n901), .Z(G395) );
  XOR2_X1 U994 ( .A(n902), .B(G286), .Z(n904) );
  XNOR2_X1 U995 ( .A(G171), .B(n978), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U997 ( .A(n905), .B(n992), .Z(n906) );
  NOR2_X1 U998 ( .A1(G37), .A2(n906), .ZN(G397) );
  XNOR2_X1 U999 ( .A(G2454), .B(G2443), .ZN(n916) );
  XOR2_X1 U1000 ( .A(G2430), .B(KEYINPUT112), .Z(n908) );
  XNOR2_X1 U1001 ( .A(G2446), .B(KEYINPUT111), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n912) );
  XOR2_X1 U1003 ( .A(G2451), .B(G2427), .Z(n910) );
  XNOR2_X1 U1004 ( .A(G1341), .B(G1348), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1006 ( .A(n912), .B(n911), .Z(n914) );
  XNOR2_X1 U1007 ( .A(G2435), .B(G2438), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1010 ( .A1(n917), .A2(G14), .ZN(n923) );
  NAND2_X1 U1011 ( .A1(n923), .A2(G319), .ZN(n920) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(n923), .ZN(G401) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(n926), .Z(n932) );
  XNOR2_X1 U1022 ( .A(G160), .B(G2084), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1026 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1027 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1028 ( .A(n937), .B(KEYINPUT121), .ZN(n939) );
  NAND2_X1 U1029 ( .A1(n939), .A2(n938), .ZN(n947) );
  XOR2_X1 U1030 ( .A(n940), .B(KEYINPUT122), .Z(n941) );
  XOR2_X1 U1031 ( .A(G2072), .B(n941), .Z(n943) );
  XNOR2_X1 U1032 ( .A(G164), .B(G2078), .ZN(n942) );
  NAND2_X1 U1033 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1034 ( .A(KEYINPUT123), .B(n944), .Z(n945) );
  XNOR2_X1 U1035 ( .A(KEYINPUT50), .B(n945), .ZN(n946) );
  NOR2_X1 U1036 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n948), .ZN(n949) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1039 ( .A1(n949), .A2(n970), .ZN(n950) );
  NAND2_X1 U1040 ( .A1(n950), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1041 ( .A(G2090), .B(G35), .ZN(n965) );
  XOR2_X1 U1042 ( .A(G25), .B(n951), .Z(n959) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(G1996), .B(G32), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(G28), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(KEYINPUT124), .B(G2072), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(G33), .B(n955), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n962) );
  XNOR2_X1 U1051 ( .A(G27), .B(n960), .ZN(n961) );
  NOR2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n963), .ZN(n964) );
  NOR2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1055 ( .A(G2084), .B(G34), .Z(n966) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(n966), .ZN(n967) );
  NAND2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(n970), .B(n969), .ZN(n972) );
  INV_X1 U1059 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1060 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n973), .ZN(n1025) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XOR2_X1 U1063 ( .A(G1966), .B(G168), .Z(n974) );
  XNOR2_X1 U1064 ( .A(KEYINPUT125), .B(n974), .ZN(n976) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(n977), .B(KEYINPUT57), .ZN(n996) );
  XNOR2_X1 U1067 ( .A(n978), .B(G1348), .ZN(n982) );
  XNOR2_X1 U1068 ( .A(G301), .B(G1961), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G299), .B(G1956), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n991) );
  AND2_X1 U1073 ( .A1(G303), .A2(G1971), .ZN(n988) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(n989), .B(KEYINPUT126), .ZN(n990) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n994) );
  XNOR2_X1 U1078 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1080 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1081 ( .A1(n998), .A2(n997), .ZN(n1023) );
  INV_X1 U1082 ( .A(G16), .ZN(n1021) );
  XNOR2_X1 U1083 ( .A(G1986), .B(G24), .ZN(n1003) );
  XNOR2_X1 U1084 ( .A(G1976), .B(G23), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(G22), .B(G1971), .ZN(n999) );
  NOR2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(KEYINPUT127), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(KEYINPUT58), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G21), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G1961), .B(G5), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1018) );
  XOR2_X1 U1094 ( .A(G1348), .B(KEYINPUT59), .Z(n1009) );
  XNOR2_X1 U1095 ( .A(G4), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(G20), .B(G1956), .ZN(n1010) );
  NOR2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(G1341), .B(G19), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT60), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1108 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

