//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT66), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n467), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n464), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n464), .ZN(new_n477));
  OAI21_X1  g052(.A(G137), .B1(new_n465), .B2(new_n466), .ZN(new_n478));
  INV_X1    g053(.A(G101), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n477), .A2(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n476), .A2(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(new_n465), .A2(new_n466), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT67), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(new_n480), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n485), .A2(new_n477), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n464), .C2(G112), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n480), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OAI22_X1  g071(.A1(new_n484), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n462), .A2(new_n463), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n499), .A2(new_n467), .A3(new_n473), .A4(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n502), .A2(G138), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT4), .B1(new_n504), .B2(new_n484), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n497), .B1(new_n501), .B2(new_n505), .ZN(G164));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n514), .A2(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n512), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n514), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n517), .A2(new_n516), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n513), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n511), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n514), .A2(new_n536), .B1(new_n520), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  AOI22_X1  g114(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n511), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n514), .A2(new_n542), .B1(new_n520), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND3_X1  g125(.A1(new_n513), .A2(G53), .A3(G543), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT68), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n529), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n518), .A2(new_n519), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n529), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(G651), .A2(new_n556), .B1(new_n558), .B2(G91), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n552), .A2(new_n553), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n553), .B1(new_n552), .B2(new_n559), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n558), .A2(G87), .ZN(new_n566));
  OAI211_X1 g141(.A(G49), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n529), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(KEYINPUT69), .B1(new_n572), .B2(G651), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n566), .B(new_n567), .C1(new_n570), .C2(new_n573), .ZN(G288));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n507), .B2(new_n508), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n509), .A2(new_n513), .A3(G86), .ZN(new_n580));
  OAI211_X1 g155(.A(G48), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n529), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n511), .B1(new_n585), .B2(KEYINPUT70), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(KEYINPUT70), .B2(new_n585), .ZN(new_n587));
  INV_X1    g162(.A(new_n514), .ZN(new_n588));
  XNOR2_X1  g163(.A(KEYINPUT71), .B(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n588), .A2(new_n589), .B1(new_n558), .B2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(G290));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(G301), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n529), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(G54), .A2(new_n588), .B1(new_n596), .B2(G651), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT72), .B(KEYINPUT10), .Z(new_n598));
  NAND3_X1  g173(.A1(new_n558), .A2(G92), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n598), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n520), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n597), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(KEYINPUT73), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(KEYINPUT73), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n593), .B1(new_n606), .B2(new_n592), .ZN(G284));
  AOI21_X1  g182(.A(new_n593), .B1(new_n606), .B2(new_n592), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI221_X1 g193(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n485), .A2(new_n477), .ZN(new_n620));
  INV_X1    g195(.A(G123), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(G135), .B2(new_n487), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT75), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT76), .B(G2096), .Z(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n467), .A2(new_n473), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(new_n481), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XOR2_X1   g205(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT77), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT78), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n644), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  OAI21_X1  g225(.A(G14), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(G401));
  XOR2_X1   g227(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n656), .B2(new_n653), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n667), .B2(new_n670), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n668), .A2(new_n669), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n676), .A2(new_n666), .A3(new_n670), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n674), .B(new_n677), .C1(new_n666), .C2(new_n676), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  XOR2_X1   g259(.A(KEYINPUT35), .B(G1991), .Z(new_n685));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n489), .A2(G119), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT84), .Z(new_n688));
  NOR2_X1   g263(.A1(G95), .A2(G2105), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT85), .Z(new_n690));
  OAI211_X1 g265(.A(new_n690), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT86), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n487), .A2(G131), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT83), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n686), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n686), .A2(G25), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT87), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n696), .A2(KEYINPUT87), .A3(new_n698), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n685), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(new_n685), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n703), .A2(new_n704), .A3(new_n699), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G6), .B(G305), .S(G16), .Z(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT32), .B(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT88), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n706), .A2(G23), .ZN(new_n715));
  INV_X1    g290(.A(G87), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n567), .B1(new_n520), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n568), .A2(new_n569), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n572), .A2(KEYINPUT69), .A3(G651), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n715), .B1(new_n720), .B2(new_n706), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n710), .A2(new_n714), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT34), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n706), .A2(G24), .ZN(new_n726));
  INV_X1    g301(.A(G290), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n706), .ZN(new_n728));
  INV_X1    g303(.A(G1986), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n702), .A2(new_n705), .A3(new_n725), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT36), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n725), .A2(new_n730), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n733), .A2(new_n702), .A3(new_n734), .A4(new_n705), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n686), .A2(G32), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n487), .A2(G141), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT92), .Z(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  INV_X1    g317(.A(G105), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n481), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n489), .B2(G129), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n738), .B1(new_n746), .B2(new_n686), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT30), .B(G28), .ZN(new_n750));
  OR2_X1    g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n750), .A2(new_n686), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n624), .B2(new_n686), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT94), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n686), .A2(G26), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT28), .Z(new_n757));
  OAI221_X1 g332(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n758));
  INV_X1    g333(.A(G140), .ZN(new_n759));
  INV_X1    g334(.A(G128), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n758), .B1(new_n486), .B2(new_n759), .C1(new_n760), .C2(new_n620), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT90), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(KEYINPUT90), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n757), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2067), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n706), .A2(G4), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n606), .B2(new_n706), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT89), .B(G1348), .Z(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n749), .A2(new_n755), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n706), .A2(G20), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT23), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n610), .B2(new_n706), .ZN(new_n774));
  INV_X1    g349(.A(G1956), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2072), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n686), .A2(G33), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  INV_X1    g355(.A(G139), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n486), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n783));
  INV_X1    g358(.A(new_n628), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n784), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(new_n464), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n782), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n783), .B2(new_n786), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n778), .B1(new_n788), .B2(G29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n686), .A2(G35), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G162), .B2(new_n686), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT29), .Z(new_n792));
  INV_X1    g367(.A(G2090), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n776), .B1(new_n777), .B2(new_n789), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n706), .A2(G5), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G171), .B2(new_n706), .ZN(new_n797));
  INV_X1    g372(.A(G1961), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n706), .A2(G21), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G168), .B2(new_n706), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT93), .B(G1966), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G34), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n804), .A2(KEYINPUT24), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(KEYINPUT24), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n686), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G160), .B2(new_n686), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n799), .B(new_n803), .C1(G2084), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G2084), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n706), .A2(G19), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n545), .B2(new_n706), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(G1341), .ZN(new_n813));
  NOR2_X1   g388(.A1(G27), .A2(G29), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G164), .B2(G29), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G2078), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(G2078), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n812), .A2(G1341), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n813), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n768), .B2(new_n769), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n789), .A2(new_n777), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n795), .A2(new_n810), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n771), .A2(new_n794), .A3(new_n822), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n736), .A2(new_n737), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n737), .B1(new_n736), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(G311));
  NAND2_X1  g401(.A1(new_n736), .A2(new_n823), .ZN(G150));
  AOI22_X1  g402(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n511), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT97), .B(G93), .Z(new_n831));
  OAI22_X1  g406(.A1(new_n514), .A2(new_n830), .B1(new_n520), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT99), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n606), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n837), .B(new_n838), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n833), .A2(KEYINPUT98), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n829), .A2(new_n832), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n840), .A2(new_n545), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n545), .B1(new_n840), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n839), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n836), .B1(new_n850), .B2(new_n852), .ZN(G145));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n746), .B(new_n788), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n693), .A2(new_n695), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n630), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n630), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n740), .A2(new_n745), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n788), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n863), .A3(new_n857), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n764), .B(G164), .ZN(new_n866));
  OAI221_X1 g441(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n867));
  INV_X1    g442(.A(G142), .ZN(new_n868));
  INV_X1    g443(.A(G130), .ZN(new_n869));
  OAI221_X1 g444(.A(new_n867), .B1(new_n486), .B2(new_n868), .C1(new_n869), .C2(new_n620), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n866), .A2(new_n870), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n624), .B(G160), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n492), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n860), .A2(new_n864), .A3(new_n871), .A4(new_n872), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n876), .B1(new_n874), .B2(new_n877), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n854), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n874), .A2(new_n877), .ZN(new_n883));
  INV_X1    g458(.A(new_n876), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n885), .A2(KEYINPUT40), .A3(new_n879), .A4(new_n878), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n882), .A2(new_n886), .ZN(G395));
  XNOR2_X1  g462(.A(G290), .B(G303), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n720), .B(G305), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(KEYINPUT42), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n892), .A2(KEYINPUT42), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n846), .B(new_n615), .Z(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n561), .B2(new_n562), .ZN(new_n899));
  INV_X1    g474(.A(new_n562), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(KEYINPUT100), .A3(new_n560), .ZN(new_n901));
  INV_X1    g476(.A(new_n603), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(G299), .A2(KEYINPUT100), .A3(new_n603), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT41), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n903), .A2(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n896), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n895), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n895), .B1(new_n909), .B2(new_n911), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n841), .A2(G868), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(G295));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n919), .A3(new_n917), .ZN(new_n920));
  INV_X1    g495(.A(new_n895), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n909), .A2(new_n911), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n592), .B1(new_n923), .B2(new_n912), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT102), .B1(new_n924), .B2(new_n916), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n920), .A2(new_n925), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  XNOR2_X1  g502(.A(G171), .B(G168), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n844), .B2(new_n845), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n840), .A2(new_n843), .ZN(new_n930));
  INV_X1    g505(.A(new_n545), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n840), .A2(new_n545), .A3(new_n843), .ZN(new_n933));
  XNOR2_X1  g508(.A(G286), .B(G171), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n904), .A3(new_n903), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n929), .B2(new_n935), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT103), .B1(new_n846), .B2(new_n934), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n891), .B(new_n937), .C1(new_n908), .C2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n942), .B2(KEYINPUT104), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n906), .B(new_n907), .C1(new_n939), .C2(new_n940), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n891), .A4(new_n937), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n937), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n890), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n943), .A2(new_n944), .A3(new_n947), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n942), .A2(KEYINPUT104), .ZN(new_n951));
  INV_X1    g526(.A(new_n907), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n952), .A2(new_n936), .A3(new_n905), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n939), .A2(new_n940), .A3(new_n910), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n890), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n951), .A2(new_n879), .A3(new_n955), .A4(new_n947), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n950), .A2(KEYINPUT106), .B1(new_n956), .B2(KEYINPUT43), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n951), .A2(new_n879), .A3(new_n947), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n944), .A4(new_n949), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n927), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n951), .A2(new_n949), .A3(new_n879), .A4(new_n947), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n962), .A2(new_n963), .A3(KEYINPUT43), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n962), .B2(KEYINPUT43), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n961), .B1(new_n927), .B2(new_n967), .ZN(G397));
  INV_X1    g543(.A(G40), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n476), .A2(new_n969), .A3(new_n482), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  XOR2_X1   g547(.A(KEYINPUT107), .B(G1384), .Z(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(G164), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT109), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n862), .A2(new_n976), .A3(G1996), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n856), .A2(new_n704), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n685), .B1(new_n693), .B2(new_n695), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n976), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n764), .A2(G2067), .ZN(new_n983));
  INV_X1    g558(.A(G2067), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n762), .A2(new_n984), .A3(new_n763), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1996), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n975), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT108), .Z(new_n989));
  AOI22_X1  g564(.A1(new_n986), .A2(new_n976), .B1(new_n989), .B2(new_n746), .ZN(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n975), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT48), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n979), .A2(new_n982), .A3(new_n990), .A4(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n989), .A2(KEYINPUT46), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n976), .B1(new_n986), .B2(new_n862), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n989), .A2(KEYINPUT46), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n998), .A2(KEYINPUT47), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(KEYINPUT47), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n979), .A2(new_n980), .A3(new_n990), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1002), .A2(new_n985), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT127), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1001), .B1(new_n1004), .B2(new_n976), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n501), .A2(new_n505), .ZN(new_n1007));
  INV_X1    g582(.A(new_n497), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n970), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G86), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n581), .B1(new_n520), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(G61), .B1(new_n517), .B2(new_n516), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n511), .B1(new_n1013), .B2(new_n577), .ZN(new_n1014));
  OAI21_X1  g589(.A(G1981), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT114), .B(G1981), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(new_n1017), .A3(KEYINPUT115), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n1019));
  NAND3_X1  g594(.A1(G305), .A2(new_n1019), .A3(G1981), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(new_n1022), .A3(new_n1020), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n1010), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT117), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1024), .A2(new_n1028), .A3(new_n1025), .A4(new_n1010), .ZN(new_n1029));
  AOI211_X1 g604(.A(G1976), .B(G288), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1017), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1010), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT113), .B1(new_n1009), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1035), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1038));
  NOR3_X1   g613(.A1(G164), .A2(G1384), .A3(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n971), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1037), .A2(new_n793), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1042));
  INV_X1    g617(.A(new_n973), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(KEYINPUT45), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n973), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(KEYINPUT111), .A3(KEYINPUT45), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n972), .B1(G164), .B2(G1384), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1050), .A2(new_n970), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1971), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1041), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n1006), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G303), .A2(G8), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT55), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n720), .A2(G1976), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1010), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  AOI221_X4 g636(.A(new_n1006), .B1(new_n720), .B2(G1976), .C1(new_n970), .C2(new_n1009), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1054), .A2(new_n1057), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1032), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1384), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1042), .A2(new_n1033), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1038), .B1(G164), .B2(G1384), .ZN(new_n1070));
  AND4_X1   g645(.A1(new_n793), .A2(new_n1069), .A3(new_n970), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT111), .B1(new_n1047), .B2(KEYINPUT45), .ZN(new_n1072));
  NOR4_X1   g647(.A1(G164), .A2(new_n1045), .A3(new_n972), .A4(new_n973), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n970), .B(new_n1050), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1074), .B2(new_n709), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT118), .B(new_n1056), .C1(new_n1075), .C2(new_n1006), .ZN(new_n1076));
  OAI211_X1 g651(.A(G8), .B(new_n1057), .C1(new_n1041), .C2(new_n1052), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1077), .A3(new_n1065), .ZN(new_n1078));
  OAI21_X1  g653(.A(G8), .B1(new_n1052), .B2(new_n1071), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT118), .B1(new_n1079), .B2(new_n1056), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G2084), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1037), .A2(new_n1082), .A3(new_n1040), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1050), .A2(new_n970), .ZN(new_n1084));
  NOR3_X1   g659(.A1(G164), .A2(new_n972), .A3(G1384), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n802), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(G168), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(G168), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT51), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1091), .A3(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1094));
  INV_X1    g669(.A(G2078), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1049), .A2(new_n1095), .A3(new_n1051), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1096), .A2(new_n1097), .B1(new_n1098), .B2(new_n798), .ZN(new_n1099));
  OR4_X1    g674(.A1(new_n1097), .A2(new_n1084), .A3(G2078), .A4(new_n1085), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1084), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT53), .B1(new_n1102), .B2(new_n1095), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1961), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n974), .A2(new_n970), .A3(KEYINPUT53), .A4(new_n1095), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1106));
  NOR4_X1   g681(.A1(new_n1103), .A2(new_n1104), .A3(G171), .A4(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1094), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1099), .A2(G301), .A3(new_n1100), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1109), .B(KEYINPUT54), .C1(G301), .C2(new_n1110), .ZN(new_n1111));
  AND4_X1   g686(.A1(new_n1081), .A2(new_n1093), .A3(new_n1108), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n552), .A2(new_n559), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1113), .B(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1102), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1069), .A2(new_n970), .A3(new_n1070), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n775), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1115), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1348), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1098), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n970), .A2(new_n984), .A3(new_n1009), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1122), .A2(new_n1123), .B1(new_n605), .B2(new_n604), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1117), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n970), .A2(new_n1009), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT58), .B(G1341), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT121), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n1131), .B(new_n1128), .C1(new_n970), .C2(new_n1009), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1051), .B(new_n987), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n545), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n545), .B(new_n1139), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1122), .A2(new_n1123), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1117), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n1120), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1115), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(KEYINPUT61), .A3(new_n1125), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1148), .A2(new_n1151), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1126), .B1(new_n1143), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1067), .B1(new_n1112), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1160), .A2(G8), .A3(G168), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1078), .A2(new_n1080), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1159), .B1(new_n1162), .B2(KEYINPUT63), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1077), .A2(new_n1065), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT118), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1075), .A2(new_n1006), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1167), .B2(new_n1057), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1168), .A3(new_n1076), .ZN(new_n1169));
  OAI211_X1 g744(.A(KEYINPUT119), .B(new_n1164), .C1(new_n1169), .C2(new_n1161), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1165), .B(new_n1171), .C1(new_n1057), .C2(new_n1054), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1163), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1090), .A2(new_n1174), .A3(new_n1092), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1165), .A2(new_n1168), .A3(new_n1076), .A4(new_n1101), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT125), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1081), .A2(new_n1175), .A3(new_n1179), .A4(new_n1101), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1093), .A2(KEYINPUT62), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1158), .A2(new_n1173), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n727), .A2(new_n729), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n975), .B1(new_n1185), .B2(new_n991), .ZN(new_n1186));
  AND4_X1   g761(.A1(new_n1186), .A2(new_n979), .A3(new_n982), .A4(new_n990), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1183), .A2(new_n1184), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1184), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1005), .B1(new_n1188), .B2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g765(.A1(G227), .A2(new_n460), .ZN(new_n1192));
  NOR3_X1   g766(.A1(G229), .A2(G401), .A3(new_n1192), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n885), .A2(new_n879), .A3(new_n878), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1195), .A2(new_n967), .ZN(G308));
  OR2_X1    g770(.A1(new_n965), .A2(new_n966), .ZN(new_n1197));
  OAI211_X1 g771(.A(new_n1194), .B(new_n1193), .C1(new_n1197), .C2(new_n964), .ZN(G225));
endmodule


