

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756;

  NOR2_X1 U371 ( .A1(n540), .A2(n355), .ZN(n542) );
  INV_X1 U372 ( .A(G953), .ZN(n746) );
  XNOR2_X2 U373 ( .A(n520), .B(n519), .ZN(n585) );
  XNOR2_X2 U374 ( .A(n390), .B(n531), .ZN(n540) );
  NOR2_X2 U375 ( .A1(n518), .A2(n719), .ZN(n520) );
  XNOR2_X2 U376 ( .A(n437), .B(n436), .ZN(n742) );
  XNOR2_X2 U377 ( .A(n424), .B(n423), .ZN(n453) );
  XNOR2_X2 U378 ( .A(KEYINPUT78), .B(G143), .ZN(n424) );
  AND2_X1 U379 ( .A1(n611), .A2(n610), .ZN(n745) );
  INV_X1 U380 ( .A(n604), .ZN(n373) );
  AND2_X2 U381 ( .A1(n661), .A2(n619), .ZN(n650) );
  NAND2_X1 U382 ( .A1(n378), .A2(n377), .ZN(n661) );
  XNOR2_X1 U383 ( .A(n394), .B(n392), .ZN(n473) );
  AND2_X1 U384 ( .A1(n386), .A2(n385), .ZN(n382) );
  XNOR2_X1 U385 ( .A(n584), .B(KEYINPUT42), .ZN(n755) );
  NOR2_X1 U386 ( .A1(n672), .A2(n561), .ZN(n708) );
  XNOR2_X1 U387 ( .A(n360), .B(n356), .ZN(n664) );
  XNOR2_X1 U388 ( .A(n473), .B(n411), .ZN(n736) );
  XNOR2_X1 U389 ( .A(n395), .B(G116), .ZN(n394) );
  NOR2_X1 U390 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U391 ( .A(G125), .B(G146), .ZN(n435) );
  XNOR2_X1 U392 ( .A(n366), .B(n365), .ZN(n364) );
  INV_X1 U393 ( .A(KEYINPUT46), .ZN(n365) );
  XNOR2_X1 U394 ( .A(n369), .B(n457), .ZN(n474) );
  INV_X1 U395 ( .A(G137), .ZN(n455) );
  AND2_X1 U396 ( .A1(n664), .A2(n663), .ZN(n666) );
  XNOR2_X1 U397 ( .A(n453), .B(G134), .ZN(n369) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n493) );
  XNOR2_X1 U399 ( .A(KEYINPUT18), .B(KEYINPUT4), .ZN(n417) );
  AND2_X1 U400 ( .A1(n397), .A2(KEYINPUT44), .ZN(n569) );
  INV_X1 U401 ( .A(KEYINPUT45), .ZN(n387) );
  XNOR2_X1 U402 ( .A(n393), .B(G119), .ZN(n392) );
  INV_X1 U403 ( .A(KEYINPUT86), .ZN(n393) );
  INV_X1 U404 ( .A(KEYINPUT10), .ZN(n436) );
  INV_X1 U405 ( .A(KEYINPUT65), .ZN(n454) );
  XNOR2_X1 U406 ( .A(G122), .B(G140), .ZN(n497) );
  INV_X1 U407 ( .A(G128), .ZN(n423) );
  XNOR2_X1 U408 ( .A(n363), .B(n362), .ZN(n611) );
  INV_X1 U409 ( .A(KEYINPUT48), .ZN(n362) );
  NAND2_X1 U410 ( .A1(n354), .A2(n364), .ZN(n363) );
  XNOR2_X1 U411 ( .A(n504), .B(n503), .ZN(n546) );
  XNOR2_X1 U412 ( .A(n502), .B(G475), .ZN(n503) );
  XNOR2_X1 U413 ( .A(n388), .B(G478), .ZN(n545) );
  NAND2_X1 U414 ( .A1(n621), .A2(n513), .ZN(n388) );
  NAND2_X1 U415 ( .A1(n571), .A2(n663), .ZN(n391) );
  OR2_X1 U416 ( .A1(n654), .A2(G902), .ZN(n396) );
  XOR2_X1 U417 ( .A(G101), .B(G110), .Z(n407) );
  XNOR2_X1 U418 ( .A(G128), .B(G119), .ZN(n441) );
  XNOR2_X1 U419 ( .A(n742), .B(KEYINPUT23), .ZN(n440) );
  XNOR2_X1 U420 ( .A(n474), .B(n459), .ZN(n743) );
  XNOR2_X1 U421 ( .A(n401), .B(n400), .ZN(n399) );
  INV_X1 U422 ( .A(KEYINPUT81), .ZN(n400) );
  NAND2_X1 U423 ( .A1(n379), .A2(KEYINPUT74), .ZN(n378) );
  NAND2_X1 U424 ( .A1(n358), .A2(n351), .ZN(n377) );
  NAND2_X1 U425 ( .A1(n357), .A2(n382), .ZN(n379) );
  NOR2_X1 U426 ( .A1(n690), .A2(n559), .ZN(n368) );
  AND2_X1 U427 ( .A1(n487), .A2(n486), .ZN(n598) );
  XNOR2_X1 U428 ( .A(n431), .B(n430), .ZN(n432) );
  INV_X1 U429 ( .A(KEYINPUT89), .ZN(n430) );
  OR2_X1 U430 ( .A1(n647), .A2(G902), .ZN(n360) );
  NAND2_X1 U431 ( .A1(n383), .A2(n384), .ZN(n381) );
  NOR2_X1 U432 ( .A1(n569), .A2(n387), .ZN(n383) );
  NOR2_X1 U433 ( .A1(G902), .A2(G237), .ZN(n429) );
  XOR2_X1 U434 ( .A(KEYINPUT72), .B(KEYINPUT95), .Z(n467) );
  XNOR2_X1 U435 ( .A(G146), .B(G101), .ZN(n468) );
  XOR2_X1 U436 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n469) );
  XNOR2_X1 U437 ( .A(n361), .B(KEYINPUT66), .ZN(n458) );
  INV_X1 U438 ( .A(G140), .ZN(n361) );
  XNOR2_X1 U439 ( .A(n420), .B(n419), .ZN(n421) );
  INV_X1 U440 ( .A(KEYINPUT17), .ZN(n419) );
  NAND2_X1 U441 ( .A1(n666), .A2(n376), .ZN(n375) );
  INV_X1 U442 ( .A(n666), .ZN(n402) );
  XNOR2_X1 U443 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U444 ( .A(n501), .B(n500), .ZN(n640) );
  XNOR2_X1 U445 ( .A(n499), .B(n403), .ZN(n500) );
  XNOR2_X1 U446 ( .A(n745), .B(KEYINPUT73), .ZN(n613) );
  XNOR2_X1 U447 ( .A(n593), .B(n522), .ZN(n586) );
  NAND2_X1 U448 ( .A1(n666), .A2(n465), .ZN(n558) );
  XNOR2_X1 U449 ( .A(n530), .B(KEYINPUT22), .ZN(n531) );
  XNOR2_X1 U450 ( .A(n446), .B(n447), .ZN(n647) );
  XNOR2_X1 U451 ( .A(n512), .B(n389), .ZN(n621) );
  XNOR2_X1 U452 ( .A(n743), .B(n463), .ZN(n654) );
  XNOR2_X1 U453 ( .A(n398), .B(KEYINPUT79), .ZN(n662) );
  NAND2_X1 U454 ( .A1(n399), .A2(n353), .ZN(n398) );
  AND2_X1 U455 ( .A1(n595), .A2(n373), .ZN(n727) );
  AND2_X1 U456 ( .A1(n367), .A2(n597), .ZN(n548) );
  AND2_X1 U457 ( .A1(n591), .A2(n374), .ZN(n350) );
  AND2_X1 U458 ( .A1(n381), .A2(n380), .ZN(n351) );
  AND2_X1 U459 ( .A1(n611), .A2(n359), .ZN(n352) );
  OR2_X1 U460 ( .A1(n745), .A2(KEYINPUT2), .ZN(n353) );
  AND2_X1 U461 ( .A1(n601), .A2(n600), .ZN(n354) );
  NAND2_X1 U462 ( .A1(n539), .A2(n373), .ZN(n355) );
  XOR2_X1 U463 ( .A(n449), .B(KEYINPUT25), .Z(n356) );
  AND2_X1 U464 ( .A1(n352), .A2(n381), .ZN(n357) );
  AND2_X1 U465 ( .A1(n382), .A2(n352), .ZN(n358) );
  AND2_X1 U466 ( .A1(n610), .A2(KEYINPUT2), .ZN(n359) );
  INV_X1 U467 ( .A(KEYINPUT104), .ZN(n376) );
  INV_X1 U468 ( .A(KEYINPUT74), .ZN(n380) );
  NAND2_X1 U469 ( .A1(n585), .A2(n755), .ZN(n366) );
  XNOR2_X1 U470 ( .A(n368), .B(KEYINPUT34), .ZN(n367) );
  XNOR2_X1 U471 ( .A(n369), .B(n511), .ZN(n389) );
  NAND2_X1 U472 ( .A1(n350), .A2(n370), .ZN(n544) );
  NAND2_X1 U473 ( .A1(n372), .A2(n371), .ZN(n370) );
  NAND2_X1 U474 ( .A1(n604), .A2(n376), .ZN(n371) );
  NAND2_X1 U475 ( .A1(n373), .A2(n375), .ZN(n372) );
  NOR2_X1 U476 ( .A1(n604), .A2(n402), .ZN(n556) );
  NAND2_X1 U477 ( .A1(n402), .A2(KEYINPUT104), .ZN(n374) );
  XNOR2_X2 U478 ( .A(n582), .B(KEYINPUT1), .ZN(n604) );
  NAND2_X1 U479 ( .A1(n382), .A2(n381), .ZN(n660) );
  INV_X1 U480 ( .A(n568), .ZN(n384) );
  NAND2_X1 U481 ( .A1(n569), .A2(n387), .ZN(n385) );
  NAND2_X1 U482 ( .A1(n568), .A2(n387), .ZN(n386) );
  OR2_X2 U483 ( .A1(n559), .A2(n391), .ZN(n390) );
  XNOR2_X1 U484 ( .A(n528), .B(n527), .ZN(n559) );
  XNOR2_X2 U485 ( .A(G113), .B(KEYINPUT3), .ZN(n395) );
  XNOR2_X2 U486 ( .A(n396), .B(n464), .ZN(n582) );
  NAND2_X1 U487 ( .A1(n553), .A2(n549), .ZN(n397) );
  XNOR2_X2 U488 ( .A(n548), .B(n547), .ZN(n553) );
  NAND2_X1 U489 ( .A1(n660), .A2(n659), .ZN(n401) );
  AND2_X1 U490 ( .A1(n604), .A2(n664), .ZN(n533) );
  AND2_X1 U491 ( .A1(n604), .A2(n402), .ZN(n667) );
  NOR2_X1 U492 ( .A1(n586), .A2(n526), .ZN(n528) );
  XOR2_X1 U493 ( .A(n498), .B(n497), .Z(n403) );
  NOR2_X1 U494 ( .A1(KEYINPUT44), .A2(KEYINPUT85), .ZN(n404) );
  XNOR2_X1 U495 ( .A(n422), .B(n421), .ZN(n426) );
  XNOR2_X1 U496 ( .A(G134), .B(KEYINPUT116), .ZN(n515) );
  INV_X1 U497 ( .A(KEYINPUT15), .ZN(n405) );
  XNOR2_X1 U498 ( .A(n405), .B(G902), .ZN(n615) );
  XNOR2_X1 U499 ( .A(G107), .B(G104), .ZN(n406) );
  XNOR2_X1 U500 ( .A(n407), .B(n406), .ZN(n735) );
  INV_X1 U501 ( .A(KEYINPUT67), .ZN(n408) );
  XNOR2_X1 U502 ( .A(n735), .B(n408), .ZN(n462) );
  XOR2_X1 U503 ( .A(KEYINPUT70), .B(KEYINPUT16), .Z(n410) );
  INV_X1 U504 ( .A(G122), .ZN(n409) );
  XNOR2_X1 U505 ( .A(n462), .B(n736), .ZN(n428) );
  INV_X1 U506 ( .A(KEYINPUT88), .ZN(n412) );
  NAND2_X1 U507 ( .A1(KEYINPUT87), .A2(n412), .ZN(n415) );
  INV_X1 U508 ( .A(KEYINPUT87), .ZN(n413) );
  NAND2_X1 U509 ( .A1(n413), .A2(KEYINPUT88), .ZN(n414) );
  NAND2_X1 U510 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U511 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U512 ( .A(n435), .B(n418), .ZN(n422) );
  NAND2_X1 U513 ( .A1(G224), .A2(n746), .ZN(n420) );
  XOR2_X1 U514 ( .A(KEYINPUT75), .B(n453), .Z(n425) );
  XNOR2_X1 U515 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U516 ( .A(n428), .B(n427), .ZN(n632) );
  NOR2_X2 U517 ( .A1(n615), .A2(n632), .ZN(n433) );
  XNOR2_X1 U518 ( .A(n429), .B(KEYINPUT71), .ZN(n477) );
  NAND2_X1 U519 ( .A1(G210), .A2(n477), .ZN(n431) );
  XNOR2_X2 U520 ( .A(n433), .B(n432), .ZN(n596) );
  INV_X1 U521 ( .A(KEYINPUT38), .ZN(n434) );
  XNOR2_X1 U522 ( .A(n596), .B(n434), .ZN(n682) );
  INV_X1 U523 ( .A(n435), .ZN(n437) );
  NAND2_X1 U524 ( .A1(G234), .A2(n746), .ZN(n438) );
  XOR2_X1 U525 ( .A(KEYINPUT8), .B(n438), .Z(n506) );
  AND2_X1 U526 ( .A1(n506), .A2(G221), .ZN(n439) );
  XNOR2_X1 U527 ( .A(n440), .B(n439), .ZN(n447) );
  XNOR2_X1 U528 ( .A(G110), .B(n458), .ZN(n444) );
  XOR2_X1 U529 ( .A(KEYINPUT92), .B(G137), .Z(n442) );
  XNOR2_X1 U530 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U531 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U532 ( .A(n445), .B(KEYINPUT24), .Z(n446) );
  INV_X1 U533 ( .A(n615), .ZN(n612) );
  NAND2_X1 U534 ( .A1(n612), .A2(G234), .ZN(n448) );
  XNOR2_X1 U535 ( .A(n448), .B(KEYINPUT20), .ZN(n450) );
  NAND2_X1 U536 ( .A1(G217), .A2(n450), .ZN(n449) );
  NAND2_X1 U537 ( .A1(G221), .A2(n450), .ZN(n452) );
  INV_X1 U538 ( .A(KEYINPUT21), .ZN(n451) );
  XNOR2_X1 U539 ( .A(n452), .B(n451), .ZN(n663) );
  XNOR2_X1 U540 ( .A(n454), .B(G131), .ZN(n496) );
  XNOR2_X1 U541 ( .A(n455), .B(KEYINPUT4), .ZN(n456) );
  XNOR2_X1 U542 ( .A(n496), .B(n456), .ZN(n457) );
  XNOR2_X1 U543 ( .A(n458), .B(KEYINPUT91), .ZN(n459) );
  NAND2_X1 U544 ( .A1(n746), .A2(G227), .ZN(n460) );
  XNOR2_X1 U545 ( .A(n460), .B(G146), .ZN(n461) );
  XNOR2_X1 U546 ( .A(n462), .B(n461), .ZN(n463) );
  INV_X1 U547 ( .A(G469), .ZN(n464) );
  INV_X1 U548 ( .A(n582), .ZN(n465) );
  XNOR2_X1 U549 ( .A(n558), .B(KEYINPUT107), .ZN(n487) );
  NAND2_X1 U550 ( .A1(G210), .A2(n493), .ZN(n466) );
  XNOR2_X1 U551 ( .A(n467), .B(n466), .ZN(n471) );
  XNOR2_X1 U552 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U553 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U554 ( .A(n473), .B(n472), .ZN(n475) );
  XNOR2_X1 U555 ( .A(n475), .B(n474), .ZN(n624) );
  OR2_X1 U556 ( .A1(n624), .A2(G902), .ZN(n476) );
  XNOR2_X2 U557 ( .A(n476), .B(G472), .ZN(n672) );
  NAND2_X1 U558 ( .A1(G214), .A2(n477), .ZN(n681) );
  AND2_X1 U559 ( .A1(n672), .A2(n681), .ZN(n478) );
  XNOR2_X1 U560 ( .A(n478), .B(KEYINPUT30), .ZN(n485) );
  NAND2_X1 U561 ( .A1(G237), .A2(G234), .ZN(n479) );
  XNOR2_X1 U562 ( .A(n479), .B(KEYINPUT90), .ZN(n480) );
  XNOR2_X1 U563 ( .A(KEYINPUT14), .B(n480), .ZN(n482) );
  AND2_X1 U564 ( .A1(n482), .A2(G953), .ZN(n481) );
  NAND2_X1 U565 ( .A1(G902), .A2(n481), .ZN(n523) );
  OR2_X1 U566 ( .A1(n523), .A2(G900), .ZN(n484) );
  NAND2_X1 U567 ( .A1(G952), .A2(n482), .ZN(n695) );
  NOR2_X1 U568 ( .A1(n695), .A2(G953), .ZN(n524) );
  INV_X1 U569 ( .A(n524), .ZN(n483) );
  NAND2_X1 U570 ( .A1(n484), .A2(n483), .ZN(n574) );
  AND2_X1 U571 ( .A1(n485), .A2(n574), .ZN(n486) );
  NAND2_X1 U572 ( .A1(n682), .A2(n598), .ZN(n489) );
  XNOR2_X1 U573 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U574 ( .A(n489), .B(n488), .ZN(n518) );
  XOR2_X1 U575 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n491) );
  XNOR2_X1 U576 ( .A(G143), .B(KEYINPUT11), .ZN(n490) );
  XNOR2_X1 U577 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U578 ( .A(n742), .B(n492), .Z(n495) );
  NAND2_X1 U579 ( .A1(n493), .A2(G214), .ZN(n494) );
  XNOR2_X1 U580 ( .A(n495), .B(n494), .ZN(n501) );
  XNOR2_X1 U581 ( .A(n496), .B(KEYINPUT97), .ZN(n499) );
  XOR2_X1 U582 ( .A(G113), .B(G104), .Z(n498) );
  NOR2_X1 U583 ( .A1(G902), .A2(n640), .ZN(n504) );
  XNOR2_X1 U584 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n502) );
  INV_X1 U585 ( .A(KEYINPUT99), .ZN(n505) );
  XNOR2_X1 U586 ( .A(n546), .B(n505), .ZN(n517) );
  XOR2_X1 U587 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n508) );
  NAND2_X1 U588 ( .A1(G217), .A2(n506), .ZN(n507) );
  XNOR2_X1 U589 ( .A(n508), .B(n507), .ZN(n512) );
  XOR2_X1 U590 ( .A(KEYINPUT7), .B(G122), .Z(n510) );
  XNOR2_X1 U591 ( .A(G107), .B(G116), .ZN(n509) );
  XNOR2_X1 U592 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U593 ( .A(G902), .ZN(n513) );
  INV_X1 U594 ( .A(n545), .ZN(n516) );
  OR2_X1 U595 ( .A1(n517), .A2(n516), .ZN(n707) );
  XNOR2_X1 U596 ( .A(n707), .B(KEYINPUT101), .ZN(n555) );
  INV_X1 U597 ( .A(n555), .ZN(n514) );
  NOR2_X1 U598 ( .A1(n518), .A2(n514), .ZN(n609) );
  XOR2_X1 U599 ( .A(n515), .B(n609), .Z(G36) );
  AND2_X1 U600 ( .A1(n517), .A2(n516), .ZN(n721) );
  INV_X1 U601 ( .A(n721), .ZN(n719) );
  XNOR2_X1 U602 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n519) );
  XNOR2_X1 U603 ( .A(n585), .B(G131), .ZN(G33) );
  INV_X1 U604 ( .A(KEYINPUT6), .ZN(n521) );
  XNOR2_X1 U605 ( .A(n672), .B(n521), .ZN(n591) );
  INV_X1 U606 ( .A(n663), .ZN(n576) );
  NAND2_X1 U607 ( .A1(n596), .A2(n681), .ZN(n593) );
  INV_X1 U608 ( .A(KEYINPUT19), .ZN(n522) );
  NOR2_X1 U609 ( .A1(G898), .A2(n523), .ZN(n525) );
  NOR2_X1 U610 ( .A1(n525), .A2(n524), .ZN(n526) );
  INV_X1 U611 ( .A(KEYINPUT0), .ZN(n527) );
  NOR2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n529) );
  XOR2_X1 U613 ( .A(n529), .B(KEYINPUT103), .Z(n571) );
  XOR2_X1 U614 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n530) );
  INV_X1 U615 ( .A(n540), .ZN(n535) );
  NOR2_X1 U616 ( .A1(n591), .A2(n540), .ZN(n532) );
  XNOR2_X1 U617 ( .A(n532), .B(KEYINPUT84), .ZN(n534) );
  INV_X1 U618 ( .A(n664), .ZN(n578) );
  AND2_X1 U619 ( .A1(n534), .A2(n533), .ZN(n565) );
  XOR2_X1 U620 ( .A(n565), .B(G101), .Z(G3) );
  AND2_X1 U621 ( .A1(n535), .A2(n578), .ZN(n537) );
  INV_X1 U622 ( .A(n672), .ZN(n579) );
  AND2_X1 U623 ( .A1(n604), .A2(n579), .ZN(n536) );
  NAND2_X1 U624 ( .A1(n537), .A2(n536), .ZN(n713) );
  XNOR2_X1 U625 ( .A(KEYINPUT77), .B(n591), .ZN(n538) );
  AND2_X1 U626 ( .A1(n578), .A2(n538), .ZN(n539) );
  INV_X1 U627 ( .A(KEYINPUT32), .ZN(n541) );
  XNOR2_X1 U628 ( .A(n542), .B(n541), .ZN(n756) );
  NAND2_X1 U629 ( .A1(n713), .A2(n756), .ZN(n550) );
  XNOR2_X1 U630 ( .A(KEYINPUT105), .B(KEYINPUT33), .ZN(n543) );
  XNOR2_X1 U631 ( .A(n544), .B(n543), .ZN(n690) );
  AND2_X1 U632 ( .A1(n546), .A2(n545), .ZN(n597) );
  XNOR2_X1 U633 ( .A(KEYINPUT76), .B(KEYINPUT35), .ZN(n547) );
  INV_X1 U634 ( .A(n550), .ZN(n549) );
  NAND2_X1 U635 ( .A1(n549), .A2(n404), .ZN(n552) );
  NAND2_X1 U636 ( .A1(n550), .A2(KEYINPUT85), .ZN(n551) );
  NAND2_X1 U637 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U638 ( .A1(n554), .A2(n553), .ZN(n567) );
  NOR2_X1 U639 ( .A1(n555), .A2(n721), .ZN(n685) );
  NAND2_X1 U640 ( .A1(n556), .A2(n672), .ZN(n674) );
  OR2_X1 U641 ( .A1(n559), .A2(n674), .ZN(n557) );
  XNOR2_X1 U642 ( .A(n557), .B(KEYINPUT31), .ZN(n724) );
  NOR2_X1 U643 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U644 ( .A(n560), .B(KEYINPUT93), .ZN(n561) );
  NOR2_X1 U645 ( .A1(n724), .A2(n708), .ZN(n562) );
  NOR2_X1 U646 ( .A1(n685), .A2(n562), .ZN(n563) );
  XNOR2_X1 U647 ( .A(n563), .B(KEYINPUT102), .ZN(n564) );
  NOR2_X1 U648 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U649 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U650 ( .A1(n681), .A2(n682), .ZN(n570) );
  XNOR2_X1 U651 ( .A(n570), .B(KEYINPUT110), .ZN(n686) );
  INV_X1 U652 ( .A(n571), .ZN(n684) );
  NOR2_X1 U653 ( .A1(n686), .A2(n684), .ZN(n573) );
  XNOR2_X1 U654 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n572) );
  XNOR2_X1 U655 ( .A(n573), .B(n572), .ZN(n698) );
  XOR2_X1 U656 ( .A(KEYINPUT28), .B(KEYINPUT108), .Z(n581) );
  INV_X1 U657 ( .A(n574), .ZN(n575) );
  NOR2_X1 U658 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U659 ( .A1(n578), .A2(n577), .ZN(n590) );
  OR2_X1 U660 ( .A1(n579), .A2(n590), .ZN(n580) );
  XOR2_X1 U661 ( .A(n581), .B(n580), .Z(n583) );
  NOR2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n698), .A2(n587), .ZN(n584) );
  INV_X1 U664 ( .A(n586), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n588), .A2(n587), .ZN(n718) );
  NOR2_X1 U666 ( .A1(n718), .A2(n685), .ZN(n589) );
  XNOR2_X1 U667 ( .A(n589), .B(KEYINPUT47), .ZN(n601) );
  NOR2_X1 U668 ( .A1(n719), .A2(n590), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n603) );
  NOR2_X1 U670 ( .A1(n603), .A2(n593), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n594), .B(KEYINPUT36), .ZN(n595) );
  AND2_X1 U672 ( .A1(n596), .A2(n597), .ZN(n599) );
  AND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n716) );
  NOR2_X1 U674 ( .A1(n727), .A2(n716), .ZN(n600) );
  INV_X1 U675 ( .A(n681), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n606) );
  XNOR2_X1 U679 ( .A(n607), .B(n606), .ZN(n608) );
  NOR2_X1 U680 ( .A1(n608), .A2(n596), .ZN(n729) );
  NOR2_X1 U681 ( .A1(n609), .A2(n729), .ZN(n610) );
  INV_X1 U682 ( .A(n660), .ZN(n730) );
  NAND2_X1 U683 ( .A1(n730), .A2(n614), .ZN(n618) );
  XNOR2_X1 U684 ( .A(n615), .B(KEYINPUT82), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n616), .A2(KEYINPUT2), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n618), .A2(n617), .ZN(n619) );
  AND2_X1 U687 ( .A1(n650), .A2(G478), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n621), .B(n620), .ZN(n623) );
  INV_X1 U689 ( .A(G952), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n622), .A2(G953), .ZN(n643) );
  INV_X1 U691 ( .A(n643), .ZN(n657) );
  NOR2_X1 U692 ( .A1(n623), .A2(n657), .ZN(G63) );
  NAND2_X1 U693 ( .A1(n650), .A2(G472), .ZN(n626) );
  XOR2_X1 U694 ( .A(n624), .B(KEYINPUT62), .Z(n625) );
  XNOR2_X1 U695 ( .A(n626), .B(n625), .ZN(n627) );
  NAND2_X1 U696 ( .A1(n627), .A2(n643), .ZN(n629) );
  XNOR2_X1 U697 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n629), .B(n628), .ZN(G57) );
  NAND2_X1 U699 ( .A1(n650), .A2(G210), .ZN(n634) );
  XNOR2_X1 U700 ( .A(KEYINPUT80), .B(KEYINPUT54), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n630), .B(KEYINPUT55), .ZN(n631) );
  XNOR2_X1 U702 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U704 ( .A1(n635), .A2(n643), .ZN(n637) );
  INV_X1 U705 ( .A(KEYINPUT56), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(G51) );
  XNOR2_X1 U707 ( .A(n553), .B(G122), .ZN(G24) );
  NAND2_X1 U708 ( .A1(n650), .A2(G475), .ZN(n642) );
  XNOR2_X1 U709 ( .A(KEYINPUT64), .B(KEYINPUT123), .ZN(n638) );
  XOR2_X1 U710 ( .A(n638), .B(KEYINPUT59), .Z(n639) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U712 ( .A(n642), .B(n641), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n646) );
  INV_X1 U714 ( .A(KEYINPUT60), .ZN(n645) );
  XNOR2_X1 U715 ( .A(n646), .B(n645), .ZN(G60) );
  NAND2_X1 U716 ( .A1(n650), .A2(G217), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X1 U718 ( .A1(n649), .A2(n657), .ZN(G66) );
  NAND2_X1 U719 ( .A1(n650), .A2(G469), .ZN(n656) );
  XOR2_X1 U720 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n652) );
  XNOR2_X1 U721 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n651) );
  XOR2_X1 U722 ( .A(n652), .B(n651), .Z(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(n658) );
  NOR2_X1 U725 ( .A1(n658), .A2(n657), .ZN(G54) );
  INV_X1 U726 ( .A(KEYINPUT2), .ZN(n659) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n703) );
  NOR2_X1 U728 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U729 ( .A(KEYINPUT49), .B(n665), .ZN(n670) );
  XOR2_X1 U730 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n668) );
  XOR2_X1 U731 ( .A(n668), .B(n667), .Z(n669) );
  NAND2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U734 ( .A(n673), .B(KEYINPUT118), .ZN(n676) );
  INV_X1 U735 ( .A(n674), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U737 ( .A(n677), .B(KEYINPUT119), .ZN(n678) );
  XNOR2_X1 U738 ( .A(n678), .B(KEYINPUT51), .ZN(n680) );
  INV_X1 U739 ( .A(n698), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n693) );
  NOR2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n684), .A2(n683), .ZN(n689) );
  NOR2_X1 U743 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U744 ( .A(n687), .B(KEYINPUT120), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X1 U746 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U747 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n694), .B(KEYINPUT52), .ZN(n696) );
  NOR2_X1 U749 ( .A1(n696), .A2(n695), .ZN(n701) );
  INV_X1 U750 ( .A(n690), .ZN(n697) );
  NAND2_X1 U751 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U752 ( .A1(n699), .A2(n746), .ZN(n700) );
  NOR2_X1 U753 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U754 ( .A1(n703), .A2(n702), .ZN(n705) );
  INV_X1 U755 ( .A(KEYINPUT53), .ZN(n704) );
  XNOR2_X1 U756 ( .A(n705), .B(n704), .ZN(G75) );
  NAND2_X1 U757 ( .A1(n708), .A2(n721), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n706), .B(G104), .ZN(G6) );
  XOR2_X1 U759 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n710) );
  INV_X1 U760 ( .A(n707), .ZN(n723) );
  NAND2_X1 U761 ( .A1(n708), .A2(n723), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U763 ( .A(G107), .B(n711), .ZN(G9) );
  XOR2_X1 U764 ( .A(G110), .B(KEYINPUT113), .Z(n712) );
  XNOR2_X1 U765 ( .A(n713), .B(n712), .ZN(G12) );
  NOR2_X1 U766 ( .A1(n707), .A2(n718), .ZN(n715) );
  XNOR2_X1 U767 ( .A(G128), .B(KEYINPUT29), .ZN(n714) );
  XNOR2_X1 U768 ( .A(n715), .B(n714), .ZN(G30) );
  XOR2_X1 U769 ( .A(G143), .B(n716), .Z(n717) );
  XNOR2_X1 U770 ( .A(KEYINPUT114), .B(n717), .ZN(G45) );
  NOR2_X1 U771 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U772 ( .A(G146), .B(n720), .Z(G48) );
  NAND2_X1 U773 ( .A1(n724), .A2(n721), .ZN(n722) );
  XNOR2_X1 U774 ( .A(n722), .B(G113), .ZN(G15) );
  XOR2_X1 U775 ( .A(G116), .B(KEYINPUT115), .Z(n726) );
  NAND2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U777 ( .A(n726), .B(n725), .ZN(G18) );
  XNOR2_X1 U778 ( .A(n727), .B(G125), .ZN(n728) );
  XNOR2_X1 U779 ( .A(n728), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U780 ( .A(G140), .B(n729), .Z(G42) );
  NAND2_X1 U781 ( .A1(n730), .A2(n746), .ZN(n734) );
  NAND2_X1 U782 ( .A1(G953), .A2(G224), .ZN(n731) );
  XNOR2_X1 U783 ( .A(KEYINPUT61), .B(n731), .ZN(n732) );
  NAND2_X1 U784 ( .A1(n732), .A2(G898), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n734), .A2(n733), .ZN(n740) );
  XNOR2_X1 U786 ( .A(n736), .B(n735), .ZN(n738) );
  NOR2_X1 U787 ( .A1(n746), .A2(G898), .ZN(n737) );
  NOR2_X1 U788 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U790 ( .A(KEYINPUT124), .B(n741), .ZN(G69) );
  XOR2_X1 U791 ( .A(n743), .B(n742), .Z(n749) );
  XNOR2_X1 U792 ( .A(n749), .B(KEYINPUT125), .ZN(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n747) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U795 ( .A(KEYINPUT126), .B(n748), .ZN(n754) );
  XNOR2_X1 U796 ( .A(n749), .B(G227), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n750), .A2(G900), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(G953), .ZN(n752) );
  XOR2_X1 U799 ( .A(KEYINPUT127), .B(n752), .Z(n753) );
  NAND2_X1 U800 ( .A1(n754), .A2(n753), .ZN(G72) );
  XNOR2_X1 U801 ( .A(G137), .B(n755), .ZN(G39) );
  XNOR2_X1 U802 ( .A(G119), .B(n756), .ZN(G21) );
endmodule

