//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT67), .A2(G116), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT67), .A2(G116), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G119), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT2), .B(G113), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n193), .B(new_n190), .C1(new_n191), .C2(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n201), .A3(G143), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n198), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n205), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n199), .A2(new_n201), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(new_n209), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n207), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(G134), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT65), .A3(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n220), .B2(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n217), .A2(KEYINPUT11), .A3(G134), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(G137), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(KEYINPUT69), .B(new_n207), .C1(new_n208), .C2(new_n212), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n215), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n211), .A2(new_n209), .ZN(new_n237));
  INV_X1    g051(.A(new_n210), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n202), .A2(new_n204), .A3(new_n233), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT68), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n225), .A2(new_n228), .A3(new_n226), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n229), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT64), .B(G146), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n238), .B1(new_n246), .B2(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n235), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(new_n240), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n242), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n232), .A2(KEYINPUT30), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n213), .A2(new_n230), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n245), .A2(new_n248), .A3(new_n240), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT30), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI211_X1 g072(.A(KEYINPUT66), .B(KEYINPUT30), .C1(new_n254), .C2(new_n255), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n197), .B(new_n252), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n261), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n197), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n232), .A2(new_n268), .A3(new_n251), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n260), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n260), .A2(KEYINPUT31), .A3(new_n267), .A4(new_n269), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n269), .A2(new_n274), .B1(new_n197), .B2(new_n256), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n232), .A2(new_n268), .A3(new_n251), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT28), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n272), .A2(new_n273), .B1(new_n266), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(G472), .A2(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n187), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n272), .A2(new_n273), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n266), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT32), .A3(new_n280), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n260), .A2(new_n287), .A3(new_n266), .A4(new_n269), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT29), .B1(new_n275), .B2(new_n277), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n269), .A2(new_n293), .A3(new_n274), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n269), .B2(new_n274), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n294), .A2(new_n295), .A3(new_n287), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n268), .B1(new_n232), .B2(new_n251), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n269), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI211_X1 g113(.A(KEYINPUT71), .B(new_n268), .C1(new_n232), .C2(new_n251), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT28), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n292), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n291), .B1(new_n302), .B2(new_n266), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n303), .A2(KEYINPUT73), .A3(G472), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT73), .B1(new_n303), .B2(G472), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n282), .B(new_n286), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT16), .ZN(new_n307));
  INV_X1    g121(.A(G125), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G140), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT76), .ZN(new_n312));
  OR3_X1    g126(.A1(new_n310), .A2(KEYINPUT76), .A3(G125), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n307), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n198), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n315), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n310), .A2(KEYINPUT76), .A3(G125), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(KEYINPUT76), .ZN(new_n320));
  OAI211_X1 g134(.A(G146), .B(new_n317), .C1(new_n320), .C2(new_n307), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n322));
  AOI21_X1  g136(.A(G143), .B1(new_n262), .B2(G214), .ZN(new_n323));
  OAI21_X1  g137(.A(G131), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT17), .ZN(new_n325));
  INV_X1    g139(.A(G237), .ZN(new_n326));
  INV_X1    g140(.A(G953), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G214), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n209), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n227), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n324), .A2(new_n325), .A3(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(KEYINPUT17), .B(G131), .C1(new_n322), .C2(new_n323), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n316), .A2(new_n321), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G113), .B(G122), .ZN(new_n335));
  INV_X1    g149(.A(G104), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n335), .B(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n320), .A2(G146), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n319), .A2(new_n246), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT18), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n322), .A2(new_n323), .B1(new_n341), .B2(new_n227), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n329), .A2(KEYINPUT18), .A3(G131), .A4(new_n330), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n334), .A2(new_n337), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT89), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n334), .A2(KEYINPUT89), .A3(new_n337), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n334), .A2(new_n345), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n337), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n289), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n353), .A2(G475), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n348), .A2(new_n349), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT87), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n357), .A2(KEYINPUT19), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(KEYINPUT19), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n319), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT86), .B1(new_n320), .B2(KEYINPUT19), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT86), .A4(KEYINPUT19), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n246), .B(new_n360), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT88), .ZN(new_n365));
  INV_X1    g179(.A(new_n360), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT19), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT86), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n369), .B2(new_n362), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT88), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n246), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n324), .A2(new_n331), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n321), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n365), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n337), .B1(new_n376), .B2(new_n345), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n355), .B1(new_n356), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(G475), .A2(G902), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n374), .B1(new_n364), .B2(KEYINPUT88), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n380), .A2(new_n372), .B1(new_n340), .B2(new_n344), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n350), .B(KEYINPUT90), .C1(new_n381), .C2(new_n337), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  XOR2_X1   g197(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT91), .ZN(new_n387));
  NOR3_X1   g201(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n387), .B(new_n388), .C1(new_n356), .C2(new_n377), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n350), .B1(new_n381), .B2(new_n337), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n387), .B1(new_n391), .B2(new_n388), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n354), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G214), .B1(G237), .B2(G902), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT82), .ZN(new_n396));
  OAI21_X1  g210(.A(G210), .B1(G237), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT3), .B1(new_n336), .B2(G107), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT3), .ZN(new_n401));
  INV_X1    g215(.A(G107), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(G104), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n336), .A2(G107), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n399), .B1(new_n405), .B2(G101), .ZN(new_n406));
  INV_X1    g220(.A(G101), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n400), .A2(new_n403), .A3(new_n407), .A4(new_n404), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n408), .A2(KEYINPUT79), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(KEYINPUT79), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n405), .A2(new_n399), .A3(G101), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n412), .A2(KEYINPUT80), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(KEYINPUT80), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n411), .A2(new_n197), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n403), .A2(new_n404), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n407), .A4(new_n400), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(KEYINPUT79), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n402), .A2(G104), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n404), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G101), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n190), .B(KEYINPUT5), .C1(new_n191), .C2(G119), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n191), .A2(KEYINPUT5), .A3(G119), .ZN(new_n425));
  INV_X1    g239(.A(G113), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n420), .A2(new_n196), .A3(new_n423), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n415), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G122), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n415), .A2(new_n429), .A3(new_n431), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G224), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(G953), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G125), .B1(new_n239), .B2(new_n241), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n308), .B(new_n207), .C1(new_n208), .C2(new_n212), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n438), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n437), .A3(new_n442), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n430), .A2(new_n449), .A3(new_n432), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n435), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n431), .B(KEYINPUT8), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n423), .B1(new_n409), .B2(new_n410), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n428), .A2(new_n196), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n457), .B2(new_n429), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT84), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n460));
  AOI211_X1 g274(.A(new_n460), .B(new_n454), .C1(new_n457), .C2(new_n429), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n439), .A2(new_n441), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT7), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(new_n437), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n439), .A2(KEYINPUT7), .A3(new_n438), .A4(new_n441), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n434), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n289), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n398), .B1(new_n452), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n455), .A2(new_n456), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n420), .A2(new_n423), .B1(new_n428), .B2(new_n196), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n453), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n458), .A2(KEYINPUT84), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n434), .A2(new_n465), .A3(new_n466), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n451), .A3(new_n397), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n396), .B1(new_n469), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n327), .A2(G952), .ZN(new_n480));
  INV_X1    g294(.A(G234), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n480), .B1(new_n481), .B2(new_n326), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n289), .B(new_n327), .C1(G234), .C2(G237), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT21), .B(G898), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n209), .A2(G128), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n205), .A2(G143), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(new_n220), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n209), .A2(KEYINPUT13), .A3(G128), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT13), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(KEYINPUT92), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT13), .B1(new_n209), .B2(G128), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT92), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n490), .B(new_n493), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n492), .B1(new_n499), .B2(G134), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n188), .A2(G122), .A3(new_n189), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n191), .A2(G122), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n402), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n502), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G107), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n489), .A2(new_n490), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G134), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n503), .A2(new_n402), .B1(new_n491), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n188), .A2(KEYINPUT14), .A3(G122), .A4(new_n189), .ZN(new_n512));
  OAI211_X1 g326(.A(G107), .B(new_n512), .C1(new_n505), .C2(KEYINPUT14), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT93), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT9), .B(G234), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(G217), .A3(new_n327), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n500), .A2(new_n507), .B1(new_n513), .B2(new_n511), .ZN(new_n521));
  INV_X1    g335(.A(new_n519), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT93), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G478), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n289), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n525), .B2(new_n289), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n488), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n525), .A2(new_n289), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n527), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT94), .A3(new_n529), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n394), .A2(new_n479), .A3(new_n487), .A4(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G221), .B1(new_n517), .B2(G902), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n203), .B1(new_n246), .B2(G143), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n205), .B1(new_n238), .B2(KEYINPUT1), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n207), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n420), .A2(new_n423), .A3(new_n541), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n418), .A2(new_n419), .B1(G101), .B2(new_n422), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n213), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n544), .A2(KEYINPUT12), .A3(new_n245), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT12), .B1(new_n544), .B2(new_n245), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT80), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n412), .B(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n549), .A2(new_n242), .A3(new_n250), .A4(new_n411), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n215), .A2(KEYINPUT10), .A3(new_n543), .A4(new_n231), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n542), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n245), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n550), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G110), .B(G140), .ZN(new_n556));
  INV_X1    g370(.A(G227), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G953), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n556), .B(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n547), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT81), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n563), .A2(new_n564), .A3(new_n245), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(new_n563), .B2(new_n245), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n555), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n562), .B1(new_n567), .B2(new_n559), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n568), .A2(G469), .A3(G902), .ZN(new_n569));
  INV_X1    g383(.A(G469), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n555), .B(new_n560), .C1(new_n565), .C2(new_n566), .ZN(new_n571));
  INV_X1    g385(.A(new_n555), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n559), .B1(new_n547), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n570), .B1(new_n574), .B2(new_n289), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n538), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n537), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT78), .ZN(new_n578));
  INV_X1    g392(.A(new_n321), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT24), .B(G110), .Z(new_n580));
  INV_X1    g394(.A(G119), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G128), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n205), .A2(G119), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT75), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n205), .A2(G119), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(G128), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n580), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n586), .B(new_n590), .C1(new_n582), .C2(KEYINPUT23), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(G110), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n339), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT77), .B1(new_n579), .B2(new_n593), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n589), .A2(new_n592), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT77), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n321), .A4(new_n339), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n316), .A2(new_n321), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n584), .A2(new_n588), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n599), .A2(new_n580), .B1(G110), .B2(new_n591), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n594), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n327), .A2(G221), .A3(G234), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT22), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G137), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n594), .A2(new_n597), .A3(new_n601), .A4(new_n605), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G217), .B1(new_n481), .B2(G902), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT74), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n611), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n607), .A2(new_n289), .A3(new_n608), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n614), .B2(KEYINPUT25), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT25), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n607), .A2(new_n616), .A3(new_n289), .A4(new_n608), .ZN(new_n617));
  AOI221_X4 g431(.A(new_n578), .B1(new_n609), .B2(new_n612), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n609), .A2(new_n612), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT78), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n306), .A2(new_n577), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT95), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  OR3_X1    g439(.A1(new_n521), .A2(KEYINPUT98), .A3(new_n522), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n522), .B1(new_n521), .B2(KEYINPUT98), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT33), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n525), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n525), .A2(KEYINPUT97), .A3(new_n630), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n526), .A2(G902), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT99), .B(G478), .Z(new_n637));
  AOI22_X1  g451(.A1(new_n635), .A2(new_n636), .B1(new_n533), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n394), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT100), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n633), .A2(new_n634), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n641), .A2(new_n628), .A3(new_n636), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n533), .A2(new_n637), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n376), .A2(new_n345), .ZN(new_n645));
  INV_X1    g459(.A(new_n337), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n645), .A2(new_n646), .B1(new_n348), .B2(new_n349), .ZN(new_n647));
  INV_X1    g461(.A(new_n388), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT91), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n389), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n383), .B2(new_n385), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n644), .B1(new_n651), .B2(new_n354), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n640), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n622), .B(new_n538), .C1(new_n569), .C2(new_n575), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n279), .B2(G902), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n285), .A2(new_n280), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n469), .A2(new_n478), .ZN(new_n663));
  INV_X1    g477(.A(new_n396), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI211_X1 g479(.A(KEYINPUT96), .B(new_n396), .C1(new_n469), .C2(new_n478), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n487), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n656), .A2(new_n661), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT34), .B(G104), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G6));
  NAND4_X1  g484(.A1(new_n378), .A2(new_n379), .A3(new_n382), .A4(new_n384), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n354), .B1(new_n386), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n532), .A2(new_n535), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n661), .A2(new_n667), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT35), .B(G107), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NOR2_X1   g492(.A1(new_n537), .A2(new_n660), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n606), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n602), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n612), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n619), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n576), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT102), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G12));
  NAND2_X1  g504(.A1(new_n286), .A2(new_n282), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT73), .ZN(new_n692));
  INV_X1    g506(.A(new_n292), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n232), .A2(new_n251), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n197), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n276), .B1(new_n695), .B2(KEYINPUT71), .ZN(new_n696));
  INV_X1    g510(.A(new_n300), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n274), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n295), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n269), .A2(new_n293), .A3(new_n274), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(KEYINPUT29), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n693), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n290), .B1(new_n702), .B2(new_n267), .ZN(new_n703));
  INV_X1    g517(.A(G472), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n692), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n303), .A2(KEYINPUT73), .A3(G472), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n691), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(G900), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n483), .B1(new_n484), .B2(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n707), .A2(new_n675), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n477), .A2(new_n397), .A3(new_n451), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n397), .B1(new_n477), .B2(new_n451), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n664), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT96), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n663), .A2(new_n662), .A3(new_n664), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n685), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  XNOR2_X1  g533(.A(new_n663), .B(KEYINPUT38), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n721), .A2(new_n396), .A3(new_n683), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n260), .A2(new_n269), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n267), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n696), .A2(new_n266), .A3(new_n697), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n289), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G472), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT103), .Z(new_n728));
  OR2_X1    g542(.A1(new_n728), .A2(new_n691), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n394), .A2(new_n536), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n722), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n569), .A2(new_n575), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n709), .B(KEYINPUT104), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n733), .B(KEYINPUT39), .Z(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n538), .A3(new_n734), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT105), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT40), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n736), .A2(KEYINPUT40), .A3(new_n737), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n731), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n209), .ZN(G45));
  NOR3_X1   g557(.A1(new_n394), .A2(new_n638), .A3(new_n709), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n717), .A2(new_n306), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G146), .ZN(G48));
  INV_X1    g560(.A(new_n622), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n705), .A2(new_n706), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n286), .A2(new_n282), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n667), .ZN(new_n751));
  OAI21_X1  g565(.A(G469), .B1(new_n568), .B2(G902), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n563), .A2(new_n245), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT81), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n563), .A2(new_n564), .A3(new_n245), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n560), .B1(new_n756), .B2(new_n555), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n570), .B(new_n289), .C1(new_n757), .C2(new_n562), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n752), .A2(new_n758), .A3(new_n538), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n750), .A2(new_n655), .A3(new_n751), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G15));
  NOR2_X1   g576(.A1(new_n667), .A2(new_n675), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n750), .A3(new_n759), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G116), .ZN(G18));
  NAND2_X1  g579(.A1(new_n386), .A2(new_n393), .ZN(new_n766));
  INV_X1    g580(.A(new_n354), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n768), .A2(new_n486), .A3(new_n673), .A4(new_n684), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n752), .A2(new_n758), .A3(new_n538), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n714), .B2(new_n715), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n306), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G119), .ZN(G21));
  AND2_X1   g587(.A1(new_n272), .A2(new_n273), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n294), .A2(new_n295), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n267), .B1(new_n301), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n280), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n619), .A2(new_n620), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n658), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n394), .A2(new_n536), .A3(new_n486), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n716), .A4(new_n759), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n771), .A2(KEYINPUT106), .A3(new_n780), .A4(new_n781), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G122), .ZN(G24));
  AND2_X1   g601(.A1(new_n771), .A2(new_n744), .ZN(new_n788));
  AOI21_X1  g602(.A(G902), .B1(new_n283), .B2(new_n284), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n301), .A2(new_n775), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n266), .A2(new_n790), .B1(new_n272), .B2(new_n273), .ZN(new_n791));
  OAI22_X1  g605(.A1(new_n789), .A2(new_n704), .B1(new_n791), .B2(new_n281), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n684), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT107), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n308), .ZN(G27));
  NOR3_X1   g610(.A1(new_n711), .A2(new_n712), .A3(new_n396), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n573), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(KEYINPUT109), .B(new_n559), .C1(new_n547), .C2(new_n572), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n799), .A2(G469), .A3(new_n571), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(G469), .A2(G902), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT108), .Z(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n538), .B(new_n797), .C1(new_n804), .C2(new_n569), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n306), .A2(new_n622), .A3(new_n806), .A4(new_n744), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT42), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n778), .B1(new_n748), .B2(new_n749), .ZN(new_n810));
  INV_X1    g624(.A(new_n709), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n768), .A2(KEYINPUT42), .A3(new_n644), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n805), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n810), .A2(KEYINPUT110), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT110), .B1(new_n810), .B2(new_n813), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n809), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G131), .ZN(G33));
  AND2_X1   g631(.A1(new_n674), .A2(new_n811), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(new_n306), .A3(new_n622), .A4(new_n806), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G134), .ZN(G36));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n570), .B1(new_n574), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n799), .A2(new_n571), .A3(new_n800), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n822), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n824), .A2(new_n803), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  OR3_X1    g640(.A1(new_n825), .A2(new_n826), .A3(KEYINPUT46), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n825), .B2(KEYINPUT46), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n569), .B1(new_n825), .B2(KEYINPUT46), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n538), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(new_n734), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n394), .A2(new_n644), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT43), .Z(new_n834));
  AOI21_X1  g648(.A(new_n684), .B1(new_n658), .B2(new_n659), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n834), .A2(KEYINPUT44), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT44), .B1(new_n834), .B2(new_n835), .ZN(new_n837));
  INV_X1    g651(.A(new_n797), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G137), .ZN(G39));
  XNOR2_X1  g655(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n831), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT47), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(KEYINPUT112), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n830), .A2(new_n538), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n707), .A2(new_n747), .A3(new_n744), .A4(new_n797), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n843), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT113), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n310), .ZN(G42));
  NOR2_X1   g664(.A1(G952), .A2(G953), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT121), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n834), .A2(new_n483), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n780), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n721), .A2(new_n396), .A3(new_n759), .ZN(new_n856));
  OR4_X1    g670(.A1(KEYINPUT119), .A2(new_n855), .A3(KEYINPUT50), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n729), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n770), .A2(new_n838), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n622), .A3(new_n483), .A4(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n768), .A3(new_n644), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n854), .A2(new_n859), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n862), .B2(new_n793), .ZN(new_n863));
  XOR2_X1   g677(.A(KEYINPUT119), .B(KEYINPUT50), .Z(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n855), .B2(new_n856), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n857), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n752), .A2(new_n758), .ZN(new_n867));
  INV_X1    g681(.A(new_n538), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n843), .B2(new_n846), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n838), .B(new_n855), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n853), .B(new_n866), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n862), .A2(new_n810), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT48), .Z(new_n876));
  NAND3_X1  g690(.A1(new_n854), .A2(new_n771), .A3(new_n780), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n480), .C1(new_n656), .C2(new_n860), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n855), .A2(new_n838), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n866), .B1(new_n870), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n879), .B1(new_n881), .B2(KEYINPUT51), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n652), .A2(new_n792), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n801), .A2(new_n803), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n868), .B1(new_n885), .B2(new_n758), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n530), .A2(new_n531), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n672), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n576), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n891), .B2(new_n707), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n797), .A2(new_n683), .A3(new_n811), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n707), .A2(new_n747), .A3(new_n805), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n892), .A2(new_n894), .B1(new_n895), .B2(new_n818), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n816), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n623), .A2(new_n772), .A3(new_n686), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n667), .B1(new_n654), .B2(new_n640), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n750), .B(new_n759), .C1(new_n899), .C2(new_n763), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n479), .A2(new_n487), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n657), .A2(new_n901), .A3(new_n660), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT115), .B1(new_n768), .B2(new_n888), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT115), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n394), .B(new_n904), .C1(new_n531), .C2(new_n530), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT114), .B1(new_n768), .B2(new_n644), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT114), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n394), .A2(new_n638), .A3(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n903), .B(new_n905), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n898), .A2(new_n900), .A3(new_n786), .A4(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT116), .B1(new_n897), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n786), .A2(new_n760), .A3(new_n764), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(new_n623), .A3(new_n686), .A4(new_n772), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n306), .A2(new_n890), .B1(new_n884), .B2(new_n886), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n819), .B1(new_n916), .B2(new_n893), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT110), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n304), .A2(new_n305), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n779), .B1(new_n919), .B2(new_n691), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n886), .A2(new_n744), .A3(KEYINPUT42), .A4(new_n797), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n810), .A2(KEYINPUT110), .A3(new_n813), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n924), .B2(new_n809), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT116), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n915), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n716), .A2(new_n730), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n683), .A2(new_n709), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT117), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n729), .A2(new_n886), .A3(new_n928), .A4(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n718), .A2(new_n931), .A3(new_n745), .A4(new_n794), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT52), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n710), .A2(new_n717), .B1(new_n788), .B2(new_n793), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n935), .A2(KEYINPUT52), .A3(new_n745), .A4(new_n931), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n912), .A2(new_n927), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT53), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT54), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT54), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n937), .A2(KEYINPUT53), .A3(new_n915), .A4(new_n925), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n938), .A2(KEYINPUT118), .A3(new_n939), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT118), .B1(new_n938), .B2(new_n939), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n942), .B(new_n943), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n852), .B1(new_n883), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n664), .A2(new_n538), .ZN(new_n949));
  NOR4_X1   g763(.A1(new_n720), .A2(new_n833), .A3(new_n778), .A4(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n867), .B(KEYINPUT49), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n858), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n948), .A2(new_n952), .ZN(G75));
  OAI21_X1  g767(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(G210), .A3(G902), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT56), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n435), .A2(new_n450), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n448), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT55), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n955), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n955), .B2(new_n956), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n327), .A2(G952), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G51));
  XOR2_X1   g777(.A(new_n803), .B(KEYINPUT57), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n938), .A2(new_n939), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT118), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n938), .A2(KEYINPUT118), .A3(new_n939), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n942), .B1(new_n969), .B2(new_n943), .ZN(new_n970));
  INV_X1    g784(.A(new_n946), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n568), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n954), .A2(G902), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n975), .A2(new_n824), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n962), .B1(new_n974), .B2(new_n976), .ZN(G54));
  NAND2_X1  g791(.A1(new_n378), .A2(new_n382), .ZN(new_n978));
  NAND2_X1  g792(.A1(KEYINPUT58), .A2(G475), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n962), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(G60));
  NAND2_X1  g798(.A1(G478), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT59), .Z(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n635), .B1(new_n947), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n635), .A2(new_n987), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n954), .A2(KEYINPUT54), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n946), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n988), .A2(new_n991), .A3(new_n962), .ZN(G63));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT60), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n954), .A2(new_n681), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n969), .B2(new_n943), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n609), .B(KEYINPUT122), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n996), .B(new_n981), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT61), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n954), .A2(new_n995), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n962), .B1(new_n1003), .B2(new_n998), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(KEYINPUT61), .A3(new_n996), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(new_n1005), .ZN(G66));
  NOR3_X1   g820(.A1(new_n485), .A2(new_n436), .A3(new_n327), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(new_n915), .B2(new_n327), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT123), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n957), .B1(G898), .B2(new_n327), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1009), .B(new_n1010), .Z(G69));
  OAI21_X1  g825(.A(new_n252), .B1(new_n258), .B2(new_n259), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT124), .Z(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(new_n370), .Z(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(G900), .B2(G953), .ZN(new_n1016));
  AND4_X1   g830(.A1(new_n745), .A2(new_n816), .A3(new_n819), .A4(new_n935), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n810), .A2(new_n928), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n832), .B1(new_n839), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n848), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1016), .B1(new_n1020), .B2(G953), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT125), .ZN(new_n1022));
  OAI21_X1  g836(.A(G953), .B1(new_n557), .B2(new_n708), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n707), .A2(new_n747), .A3(new_n838), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n736), .A2(new_n737), .A3(new_n909), .ZN(new_n1025));
  AOI22_X1  g839(.A1(new_n832), .A2(new_n839), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n935), .A2(new_n745), .ZN(new_n1027));
  OAI21_X1  g841(.A(KEYINPUT62), .B1(new_n742), .B2(new_n1027), .ZN(new_n1028));
  OR3_X1    g842(.A1(new_n742), .A2(KEYINPUT62), .A3(new_n1027), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n848), .A2(new_n1026), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1030), .A2(new_n327), .ZN(new_n1031));
  OAI221_X1 g845(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .C1(new_n1031), .C2(new_n1014), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1023), .A2(new_n1022), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1032), .B(new_n1033), .ZN(G72));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  OAI21_X1  g850(.A(new_n1036), .B1(new_n1020), .B2(new_n911), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n723), .A2(new_n267), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n962), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT126), .ZN(new_n1040));
  INV_X1    g854(.A(new_n724), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1040), .B1(new_n1041), .B2(new_n1038), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n723), .A2(KEYINPUT126), .A3(new_n266), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n940), .A2(new_n1042), .A3(new_n1036), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1036), .B1(new_n1030), .B2(new_n911), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1045), .A2(new_n1041), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1039), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g861(.A(KEYINPUT127), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1047), .B(new_n1048), .ZN(G57));
endmodule


