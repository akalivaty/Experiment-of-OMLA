//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n450), .B(new_n451), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT65), .Z(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(G137), .A3(new_n460), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n460), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(new_n468), .ZN(G160));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n460), .A2(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n472), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n460), .A2(G138), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n461), .A2(KEYINPUT4), .A3(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n460), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n485), .A2(new_n486), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  INV_X1    g067(.A(G651), .ZN(new_n493));
  NAND2_X1  g068(.A1(G75), .A2(G543), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT66), .Z(new_n495));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G62), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n493), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n504), .A2(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n502), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  INV_X1    g091(.A(G89), .ZN(new_n517));
  INV_X1    g092(.A(G51), .ZN(new_n518));
  OAI221_X1 g093(.A(new_n516), .B1(new_n510), .B2(new_n517), .C1(new_n518), .C2(new_n504), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT67), .B1(new_n507), .B2(new_n506), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n498), .A2(new_n521), .A3(new_n499), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G63), .ZN(new_n524));
  NOR3_X1   g099(.A1(new_n523), .A2(new_n524), .A3(new_n493), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G168));
  NAND3_X1  g101(.A1(new_n520), .A2(new_n522), .A3(G64), .ZN(new_n527));
  NAND2_X1  g102(.A1(G77), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT68), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n527), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(G651), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n504), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT69), .B(G52), .ZN(new_n535));
  INV_X1    g110(.A(new_n510), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n534), .A2(new_n535), .B1(new_n536), .B2(G90), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n533), .A2(KEYINPUT70), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT70), .B1(new_n533), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND3_X1  g116(.A1(new_n520), .A2(new_n522), .A3(G56), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n493), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n504), .A2(new_n545), .B1(new_n510), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n504), .A2(KEYINPUT9), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n504), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n510), .A2(KEYINPUT71), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n500), .A2(new_n503), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(G91), .A3(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n500), .A2(G65), .ZN(new_n562));
  AND2_X1   g137(.A1(G78), .A2(G543), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n557), .A2(new_n561), .A3(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(new_n523), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n567), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n558), .A2(G87), .A3(new_n560), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n534), .A2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n558), .A2(G86), .A3(new_n560), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n503), .A2(G48), .A3(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G61), .B1(new_n507), .B2(new_n506), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n575), .A2(new_n576), .B1(G73), .B2(G543), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n500), .A2(KEYINPUT72), .A3(G61), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n493), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n582));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n523), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n493), .B1(new_n585), .B2(new_n586), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n504), .A2(new_n590), .B1(new_n510), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n582), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  AOI211_X1 g169(.A(KEYINPUT74), .B(new_n592), .C1(new_n587), .C2(new_n588), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NOR2_X1   g173(.A1(G301), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n558), .A2(G92), .A3(new_n560), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n500), .A2(G66), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT76), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n493), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n534), .A2(KEYINPUT75), .ZN(new_n607));
  INV_X1    g182(.A(G54), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n504), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n606), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n599), .B1(new_n598), .B2(new_n614), .ZN(G284));
  AOI21_X1  g190(.A(new_n599), .B1(new_n598), .B2(new_n614), .ZN(G321));
  NAND2_X1  g191(.A1(G299), .A2(new_n598), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n598), .B2(G168), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(new_n598), .B2(G168), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n614), .B1(new_n620), .B2(G860), .ZN(G148));
  INV_X1    g196(.A(new_n548), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n598), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n612), .B(KEYINPUT77), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n623), .B1(new_n625), .B2(new_n598), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n461), .A2(new_n466), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT13), .Z(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n477), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n460), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G123), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n461), .A2(G2105), .ZN(new_n638));
  OAI221_X1 g213(.A(new_n634), .B1(new_n635), .B2(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT78), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(G401));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n631), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n640), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n672), .A2(new_n673), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n674), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(KEYINPUT79), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(new_n677), .B2(new_n678), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT80), .ZN(new_n687));
  XOR2_X1   g262(.A(G1981), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n687), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  NOR2_X1   g269(.A1(G16), .A2(G19), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n548), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1341), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G26), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n473), .A2(G128), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT84), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(G116), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G2105), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G140), .B2(new_n477), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n700), .B1(new_n707), .B2(G29), .ZN(new_n708));
  INV_X1    g283(.A(G2067), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n698), .A2(G35), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G162), .B2(new_n698), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT29), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n697), .B(new_n710), .C1(G2090), .C2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G20), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT23), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n557), .A2(new_n561), .A3(new_n564), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n715), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1956), .ZN(new_n720));
  INV_X1    g295(.A(G2078), .ZN(new_n721));
  NAND2_X1  g296(.A1(G164), .A2(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G27), .B2(G29), .ZN(new_n723));
  INV_X1    g298(.A(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n724), .B2(KEYINPUT24), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(KEYINPUT24), .B2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G160), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n698), .ZN(new_n728));
  INV_X1    g303(.A(G2084), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n721), .A2(new_n723), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n730), .B(new_n731), .C1(new_n721), .C2(new_n723), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n698), .A2(G33), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n477), .A2(G139), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n461), .A2(G127), .ZN(new_n738));
  NAND2_X1  g313(.A1(G115), .A2(G2104), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n460), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n733), .B1(new_n741), .B2(new_n698), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2072), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n720), .A2(new_n732), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n713), .A2(G2090), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT91), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n698), .A2(G32), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n466), .A2(G105), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT26), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n748), .B(new_n750), .C1(G129), .C2(new_n473), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n477), .A2(G141), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT85), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT86), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n747), .B1(new_n756), .B2(new_n698), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT27), .B(G1996), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT87), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n757), .B(new_n759), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n714), .A2(new_n744), .A3(new_n746), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n715), .A2(G4), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n614), .B2(new_n715), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1348), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(G301), .A2(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n715), .A2(G5), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT88), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G16), .B2(G21), .ZN(new_n771));
  NAND2_X1  g346(.A1(G168), .A2(G16), .ZN(new_n772));
  MUX2_X1   g347(.A(new_n770), .B(new_n771), .S(new_n772), .Z(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT89), .B(G28), .Z(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n778), .B2(KEYINPUT30), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(KEYINPUT30), .B2(new_n778), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n777), .B(new_n780), .C1(new_n639), .C2(new_n698), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n769), .A2(new_n775), .A3(new_n776), .A4(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT90), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(KEYINPUT90), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n767), .A2(new_n766), .A3(new_n768), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n765), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G23), .B(G288), .S(G16), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT33), .B(G1976), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT82), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n787), .B(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT83), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(KEYINPUT83), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n715), .A2(G6), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n580), .B2(new_n715), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT32), .B(G1981), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n715), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n715), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1971), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n794), .A2(new_n795), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n791), .A2(new_n792), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n698), .A2(G25), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n477), .A2(G131), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n460), .A2(G107), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  INV_X1    g382(.A(G119), .ZN(new_n808));
  OAI221_X1 g383(.A(new_n805), .B1(new_n806), .B2(new_n807), .C1(new_n808), .C2(new_n638), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT81), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n804), .B1(new_n811), .B2(new_n698), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  XOR2_X1   g388(.A(new_n812), .B(new_n813), .Z(new_n814));
  NOR2_X1   g389(.A1(new_n596), .A2(new_n715), .ZN(new_n815));
  INV_X1    g390(.A(G1986), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n715), .A2(G24), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n816), .B1(new_n815), .B2(new_n817), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n803), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n803), .A2(new_n824), .A3(new_n820), .A4(new_n821), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n786), .B1(new_n823), .B2(new_n825), .ZN(G311));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n825), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n765), .A2(new_n784), .A3(new_n785), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n827), .A2(new_n828), .A3(new_n783), .ZN(G150));
  XNOR2_X1  g404(.A(KEYINPUT94), .B(G55), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n534), .A2(new_n830), .B1(new_n536), .B2(G93), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT93), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n520), .A2(new_n522), .A3(G67), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n832), .B1(new_n835), .B2(G651), .ZN(new_n836));
  AOI211_X1 g411(.A(KEYINPUT93), .B(new_n493), .C1(new_n833), .C2(new_n834), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT97), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n614), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT92), .B(KEYINPUT38), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n835), .A2(G651), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT93), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n835), .A2(new_n832), .A3(G651), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT95), .B1(new_n544), .B2(new_n547), .ZN(new_n850));
  OR3_X1    g425(.A1(new_n544), .A2(KEYINPUT95), .A3(new_n547), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n831), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n838), .A2(KEYINPUT95), .A3(new_n622), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n845), .B(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  INV_X1    g431(.A(G860), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n842), .B1(new_n856), .B2(new_n858), .ZN(G145));
  XOR2_X1   g434(.A(new_n755), .B(KEYINPUT86), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n741), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n707), .B(new_n491), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n755), .A2(new_n741), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n741), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n756), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n862), .B1(new_n868), .B2(new_n864), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n809), .B(KEYINPUT99), .ZN(new_n871));
  INV_X1    g446(.A(new_n629), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  INV_X1    g451(.A(G118), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(G2105), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(G142), .B2(new_n477), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n473), .A2(KEYINPUT98), .A3(G130), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT98), .B1(new_n473), .B2(G130), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n874), .A2(new_n875), .A3(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n871), .A2(new_n872), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n885), .B2(new_n873), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n870), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT100), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n886), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n866), .A2(new_n890), .A3(new_n869), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n866), .A2(new_n890), .A3(new_n869), .A4(KEYINPUT101), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n870), .A2(new_n895), .A3(new_n887), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n889), .A2(new_n893), .A3(new_n894), .A4(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n639), .B(G160), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n481), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n866), .A2(new_n890), .A3(new_n869), .A4(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n888), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT40), .B1(new_n900), .B2(new_n906), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(G395));
  NAND2_X1  g484(.A1(new_n838), .A2(new_n598), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n612), .A2(new_n718), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n602), .A2(G299), .A3(new_n611), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(KEYINPUT103), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n913), .B(new_n914), .C1(KEYINPUT103), .C2(new_n911), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n912), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n854), .B1(new_n624), .B2(G559), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n614), .A2(new_n620), .A3(new_n853), .A4(new_n852), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT105), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n916), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n920), .A2(new_n923), .A3(new_n927), .A4(new_n922), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n589), .A2(new_n593), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT74), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n589), .A2(new_n582), .A3(new_n593), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(G305), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n580), .B1(new_n594), .B2(new_n595), .ZN(new_n934));
  XNOR2_X1  g509(.A(G288), .B(G303), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n938), .B(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n929), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n910), .B1(new_n941), .B2(new_n598), .ZN(G295));
  OAI21_X1  g517(.A(new_n910), .B1(new_n941), .B2(new_n598), .ZN(G331));
  INV_X1    g518(.A(new_n938), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n538), .B2(new_n539), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n533), .A2(new_n537), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT70), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n533), .A2(KEYINPUT70), .A3(new_n537), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT106), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n852), .A2(new_n853), .A3(G286), .ZN(new_n953));
  AOI21_X1  g528(.A(G286), .B1(new_n852), .B2(new_n853), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n854), .A2(G168), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n852), .A2(new_n853), .A3(G286), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n956), .A2(new_n946), .A3(new_n951), .A4(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n958), .A3(new_n918), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n916), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n913), .B1(KEYINPUT103), .B2(new_n911), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n955), .A2(new_n958), .A3(KEYINPUT41), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n944), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n956), .A2(new_n957), .B1(new_n946), .B2(new_n951), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n917), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n955), .A2(new_n958), .A3(new_n915), .A4(new_n919), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n938), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NOR4_X1   g544(.A1(new_n963), .A2(new_n968), .A3(new_n969), .A4(G37), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n967), .ZN(new_n971));
  AOI21_X1  g546(.A(G37), .B1(new_n971), .B2(new_n944), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n966), .A2(new_n967), .A3(new_n938), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT43), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT44), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  NOR4_X1   g551(.A1(new_n963), .A2(new_n968), .A3(KEYINPUT43), .A4(G37), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n979), .ZN(G397));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n491), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G125), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n463), .B1(new_n472), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G2105), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n477), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(G40), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1996), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT107), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n756), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n990), .A2(new_n755), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(new_n991), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT108), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n707), .B(new_n709), .ZN(new_n999));
  INV_X1    g574(.A(new_n990), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n809), .B(new_n813), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n990), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n995), .A2(new_n998), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G290), .A2(G1986), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n596), .A2(new_n816), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1000), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT124), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n989), .B1(new_n982), .B2(KEYINPUT50), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n491), .A2(new_n1015), .A3(new_n981), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n766), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(G2078), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n989), .B1(new_n982), .B2(new_n983), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n491), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n491), .A2(KEYINPUT117), .A3(KEYINPUT45), .A4(new_n981), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1018), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n984), .A2(KEYINPUT110), .ZN(new_n1029));
  INV_X1    g604(.A(G40), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n464), .A2(new_n468), .A3(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1023), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n982), .A2(new_n1033), .A3(new_n983), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1029), .A2(new_n1032), .A3(new_n721), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n1019), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT123), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(KEYINPUT123), .A3(new_n1019), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1028), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1013), .B1(new_n1040), .B2(G301), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1028), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1035), .A2(KEYINPUT123), .A3(new_n1019), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT123), .B1(new_n1035), .B2(new_n1019), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1022), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1018), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G301), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1012), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(G160), .A2(G40), .A3(new_n981), .A4(new_n491), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n568), .A2(G1976), .A3(new_n569), .A4(new_n570), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1054), .B(G8), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT52), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n982), .A2(new_n989), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n1069));
  INV_X1    g644(.A(G1981), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n500), .A2(new_n503), .A3(G86), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1071), .A2(new_n573), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1071), .B2(new_n573), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n577), .A2(new_n578), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G651), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n574), .A2(G1981), .A3(new_n579), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1069), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1077), .A2(new_n1070), .A3(new_n572), .A4(new_n573), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n579), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1081), .B(KEYINPUT49), .C1(new_n1082), .C2(new_n1070), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1083), .A3(new_n1063), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1080), .A2(KEYINPUT114), .A3(new_n1083), .A4(new_n1063), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1068), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G303), .A2(G8), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT55), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1014), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1016), .A2(new_n1092), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1016), .A2(new_n1092), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT111), .B(G2090), .Z(new_n1096));
  NAND3_X1  g671(.A1(new_n1029), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1097));
  INV_X1    g672(.A(G1971), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1095), .A2(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1090), .B1(new_n1099), .B2(new_n1062), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1090), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1103), .A2(new_n1031), .A3(new_n1016), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(new_n1096), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1101), .B(G8), .C1(new_n1102), .C2(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1088), .A2(new_n1100), .A3(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1042), .B(G301), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1108), .B(KEYINPUT54), .C1(new_n1050), .C2(G301), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT118), .B(G2084), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1027), .A2(new_n774), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(G8), .B1(new_n1113), .B2(G286), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1104), .A2(new_n1110), .B1(new_n1027), .B2(new_n774), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(G168), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1062), .B1(new_n1115), .B2(G168), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1107), .A2(new_n1109), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n718), .B(KEYINPUT57), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1016), .B(new_n1092), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1014), .ZN(new_n1125));
  INV_X1    g700(.A(G1956), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1029), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1123), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n982), .A2(new_n989), .A3(G2067), .ZN(new_n1132));
  INV_X1    g707(.A(G1348), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1132), .B1(new_n1017), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(KEYINPUT120), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1136), .B(new_n1132), .C1(new_n1017), .C2(new_n1133), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1135), .A2(new_n1137), .A3(new_n612), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1127), .A2(new_n1130), .A3(new_n1123), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1131), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT58), .B(G1341), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1097), .A2(G1996), .B1(new_n1061), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n548), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1144), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(new_n548), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n1149));
  INV_X1    g724(.A(new_n612), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(KEYINPUT60), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n612), .A2(KEYINPUT122), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n612), .A2(new_n1152), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1154), .B(new_n1156), .C1(new_n1137), .C2(new_n1135), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1148), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1129), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1097), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(G1956), .B1(new_n1124), .B2(new_n1014), .ZN(new_n1164));
  XNOR2_X1  g739(.A(G299), .B(KEYINPUT57), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1166), .B2(new_n1131), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1139), .A2(new_n1168), .A3(KEYINPUT61), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1140), .B1(new_n1160), .B2(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1053), .A2(new_n1122), .A3(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1088), .A2(new_n1100), .A3(new_n1106), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1113), .A2(G8), .A3(G168), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(G8), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n1090), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1178), .A2(new_n1180), .A3(new_n1088), .A4(new_n1106), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1113), .A2(G286), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1119), .B1(new_n1118), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1114), .A2(KEYINPUT51), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT62), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1117), .A2(new_n1187), .A3(new_n1120), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1047), .A2(new_n1186), .A3(new_n1107), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1190));
  NOR2_X1   g765(.A1(G288), .A2(G1976), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1081), .B(KEYINPUT115), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1106), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1194), .A2(new_n1063), .B1(new_n1195), .B2(new_n1088), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1182), .A2(new_n1189), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1011), .B1(new_n1172), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1005), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1005), .A2(new_n1199), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1007), .A2(new_n1000), .ZN(new_n1202));
  XNOR2_X1  g777(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1202), .B(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1200), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(new_n996), .ZN(new_n1206));
  OR3_X1    g781(.A1(new_n1001), .A2(KEYINPUT125), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n994), .A2(KEYINPUT46), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT46), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n993), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(KEYINPUT125), .B1(new_n1001), .B2(new_n1206), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1212), .B(KEYINPUT47), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n995), .A2(new_n998), .A3(new_n1002), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n811), .A2(new_n813), .ZN(new_n1215));
  OAI22_X1  g790(.A1(new_n1214), .A2(new_n1215), .B1(G2067), .B2(new_n707), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n990), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1205), .A2(new_n1213), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1198), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g794(.A1(new_n977), .A2(new_n978), .ZN(new_n1221));
  OR2_X1    g795(.A1(G227), .A2(new_n458), .ZN(new_n1222));
  NOR3_X1   g796(.A1(G229), .A2(G401), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g797(.A(new_n896), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n895), .B1(new_n870), .B2(new_n887), .ZN(new_n1225));
  NOR2_X1   g799(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AND2_X1   g800(.A1(new_n893), .A2(new_n894), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n901), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g802(.A(G37), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n888), .A2(new_n901), .A3(new_n903), .ZN(new_n1230));
  INV_X1    g804(.A(new_n905), .ZN(new_n1231));
  OAI21_X1  g805(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g806(.A(new_n1223), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1233));
  NOR2_X1   g807(.A1(new_n1221), .A2(new_n1233), .ZN(G308));
  OAI221_X1 g808(.A(new_n1223), .B1(new_n1228), .B2(new_n1232), .C1(new_n977), .C2(new_n978), .ZN(G225));
endmodule


