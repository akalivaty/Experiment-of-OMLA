//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n605, new_n606, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1114, new_n1115, new_n1116;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT68), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n468), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n468), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n471), .A2(G137), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n467), .B(new_n474), .C1(new_n472), .C2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n471), .A2(new_n473), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n472), .ZN(new_n488));
  AOI211_X1 g063(.A(new_n481), .B(new_n487), .C1(G124), .C2(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n492));
  AOI21_X1  g067(.A(KEYINPUT67), .B1(new_n492), .B2(G2104), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(G2104), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n473), .B(new_n491), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n471), .A2(new_n497), .A3(new_n473), .A4(new_n491), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n496), .A2(new_n498), .A3(new_n501), .A4(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n475), .A2(new_n503), .A3(new_n491), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(G114), .A2(G2104), .ZN(new_n506));
  INV_X1    g081(.A(G126), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n482), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G2105), .B1(G102), .B2(new_n465), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n521), .A2(G543), .ZN(new_n523));
  AOI22_X1  g098(.A1(G88), .A2(new_n522), .B1(new_n523), .B2(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n516), .A2(KEYINPUT73), .A3(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n513), .A2(new_n515), .ZN(new_n528));
  INV_X1    g103(.A(G62), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n525), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G651), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n524), .A2(new_n532), .ZN(G166));
  NAND2_X1  g108(.A1(new_n522), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n523), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n516), .A2(new_n521), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n521), .A2(G543), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT74), .B(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n517), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(G171));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n541), .A2(new_n549), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT75), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n517), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n523), .A2(G53), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n516), .A2(new_n521), .A3(G91), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT76), .Z(new_n565));
  AOI22_X1  g140(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n563), .B(new_n565), .C1(new_n517), .C2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G166), .ZN(G303));
  AOI22_X1  g144(.A1(G87), .A2(new_n522), .B1(new_n523), .B2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n528), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n522), .A2(G86), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n518), .A2(new_n520), .A3(G48), .A4(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G305));
  XNOR2_X1  g157(.A(KEYINPUT79), .B(G85), .ZN(new_n583));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n541), .A2(new_n583), .B1(new_n543), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n517), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n585), .A2(new_n587), .ZN(G290));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n541), .A2(KEYINPUT10), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n528), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n523), .A2(G54), .B1(new_n593), .B2(G651), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT10), .B1(new_n541), .B2(new_n589), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G171), .B2(new_n597), .ZN(G321));
  XNOR2_X1  g174(.A(G321), .B(KEYINPUT80), .ZN(G284));
  NAND2_X1  g175(.A1(G299), .A2(new_n597), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n597), .B2(G168), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n597), .B2(G168), .ZN(G280));
  INV_X1    g178(.A(new_n596), .ZN(new_n604));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G860), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT81), .ZN(G148));
  OAI21_X1  g182(.A(G868), .B1(new_n596), .B2(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n555), .B2(G868), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n488), .A2(G123), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n486), .A2(G135), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n472), .A2(G111), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2096), .Z(new_n616));
  NAND2_X1  g191(.A1(new_n475), .A2(new_n465), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT13), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT15), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2435), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(KEYINPUT14), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n629), .B(new_n630), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n628), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G1341), .B(G1348), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT83), .Z(new_n636));
  OR2_X1    g211(.A1(new_n632), .A2(new_n634), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n636), .A2(new_n638), .ZN(G401));
  XNOR2_X1  g214(.A(G2072), .B(G2078), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  OAI211_X1 g218(.A(KEYINPUT17), .B(new_n640), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n643), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT17), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n641), .ZN(new_n647));
  OAI221_X1 g222(.A(new_n644), .B1(new_n645), .B2(new_n641), .C1(new_n647), .C2(new_n640), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n642), .A2(new_n640), .A3(new_n643), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2096), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT85), .ZN(new_n656));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  AND2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n656), .A2(new_n657), .ZN(new_n663));
  AOI22_X1  g238(.A1(new_n661), .A2(new_n662), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  OR3_X1    g239(.A1(new_n658), .A2(new_n663), .A3(new_n660), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n665), .C1(new_n662), .C2(new_n661), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  INV_X1    g244(.A(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n668), .B(new_n672), .ZN(G229));
  NOR2_X1   g248(.A1(G5), .A2(G16), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(G171), .B2(G16), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(G1961), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G28), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT93), .Z(new_n679));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n679), .B(new_n680), .C1(new_n677), .C2(G28), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G11), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n681), .B(new_n682), .C1(new_n615), .C2(new_n680), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT94), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G21), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G168), .B2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(G1966), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n675), .A2(G1961), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT95), .Z(new_n692));
  NAND3_X1  g267(.A1(new_n685), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT96), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(G299), .A2(G16), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n686), .A2(KEYINPUT23), .A3(G20), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT23), .ZN(new_n698));
  INV_X1    g273(.A(G20), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G16), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n696), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT98), .ZN(new_n702));
  INV_X1    g277(.A(G1956), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(G29), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n488), .A2(G129), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n486), .A2(G141), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n465), .A2(G105), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT26), .Z(new_n710));
  NAND4_X1  g285(.A1(new_n706), .A2(new_n707), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(new_n680), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G1996), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n686), .A2(G4), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n604), .B2(new_n686), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT90), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT89), .B(G1348), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n704), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n702), .A2(new_n703), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n717), .A2(new_n719), .ZN(new_n723));
  OR2_X1    g298(.A1(KEYINPUT24), .A2(G34), .ZN(new_n724));
  NAND2_X1  g299(.A1(KEYINPUT24), .A2(G34), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n724), .A2(new_n680), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G160), .B2(new_n680), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT28), .ZN(new_n728));
  INV_X1    g303(.A(G26), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G29), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n488), .A2(G128), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n486), .A2(G140), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n472), .A2(G116), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(G29), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n730), .B1(new_n737), .B2(new_n728), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n723), .B1(G2084), .B2(new_n727), .C1(new_n738), .C2(G2067), .ZN(new_n739));
  NOR4_X1   g314(.A1(new_n695), .A2(new_n721), .A3(new_n722), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n686), .A2(G19), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n555), .B2(new_n686), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G1341), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n693), .A2(new_n694), .ZN(new_n744));
  AND4_X1   g319(.A1(new_n676), .A2(new_n740), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n686), .A2(G22), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G166), .B2(new_n686), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1971), .Z(new_n748));
  NOR2_X1   g323(.A1(G16), .A2(G23), .ZN(new_n749));
  INV_X1    g324(.A(G288), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT33), .B(G1976), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G6), .A2(G16), .ZN(new_n754));
  INV_X1    g329(.A(G305), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G16), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT32), .B(G1981), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n748), .A2(new_n753), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT34), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n488), .A2(G119), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n486), .A2(G131), .ZN(new_n762));
  OR2_X1    g337(.A1(G95), .A2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n763), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(new_n680), .ZN(new_n766));
  OR2_X1    g341(.A1(G25), .A2(G29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(KEYINPUT86), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(KEYINPUT86), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT35), .B(G1991), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OR3_X1    g347(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n686), .A2(G24), .ZN(new_n775));
  INV_X1    g350(.A(G290), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n686), .ZN(new_n777));
  MUX2_X1   g352(.A(new_n775), .B(new_n777), .S(KEYINPUT87), .Z(new_n778));
  INV_X1    g353(.A(G1986), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n760), .A2(new_n773), .A3(new_n774), .A4(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G27), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT97), .B1(new_n784), .B2(G29), .ZN(new_n785));
  OR3_X1    g360(.A1(new_n784), .A2(KEYINPUT97), .A3(G29), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n785), .B(new_n786), .C1(G164), .C2(new_n680), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G2078), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n738), .A2(G2067), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n745), .A2(new_n783), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n486), .A2(G139), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n465), .A2(G103), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  AOI22_X1  g368(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n791), .B(new_n793), .C1(new_n472), .C2(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G33), .B(new_n795), .S(G29), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT91), .B(G2072), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n712), .A2(new_n713), .B1(G2084), .B2(new_n727), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT92), .Z(new_n801));
  NOR2_X1   g376(.A1(new_n787), .A2(G2078), .ZN(new_n802));
  NOR2_X1   g377(.A1(G29), .A2(G35), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G162), .B2(G29), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT29), .B(G2090), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n790), .A2(new_n801), .A3(new_n802), .A4(new_n807), .ZN(G311));
  NOR2_X1   g383(.A1(new_n790), .A2(new_n807), .ZN(new_n809));
  INV_X1    g384(.A(new_n801), .ZN(new_n810));
  INV_X1    g385(.A(new_n802), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(G150));
  AOI22_X1  g387(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n517), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT99), .Z(new_n815));
  AOI22_X1  g390(.A1(G93), .A2(new_n522), .B1(new_n523), .B2(G55), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT101), .B(G860), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n817), .B(new_n555), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n596), .A2(new_n605), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT39), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n823), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n822), .B(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n821), .B1(new_n827), .B2(new_n818), .ZN(G145));
  INV_X1    g403(.A(G37), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n488), .A2(G130), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n486), .A2(G142), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n472), .A2(G118), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n765), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT105), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n618), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n505), .A2(new_n838), .A3(new_n509), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n505), .B2(new_n509), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n795), .A2(KEYINPUT104), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n736), .B(new_n711), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n843), .B(new_n844), .Z(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n837), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n836), .A2(new_n618), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n836), .A2(new_n618), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n615), .B(G160), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G162), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n847), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n847), .A2(KEYINPUT106), .A3(new_n850), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n852), .B1(new_n850), .B2(KEYINPUT106), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n829), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g433(.A1(new_n817), .A2(new_n597), .ZN(new_n859));
  XNOR2_X1  g434(.A(G166), .B(new_n755), .ZN(new_n860));
  XNOR2_X1  g435(.A(G288), .B(G290), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(KEYINPUT107), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(KEYINPUT107), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT108), .ZN(new_n865));
  MUX2_X1   g440(.A(new_n864), .B(new_n865), .S(KEYINPUT42), .Z(new_n866));
  NOR2_X1   g441(.A1(new_n596), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n822), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G299), .B(new_n596), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(KEYINPUT41), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n866), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n859), .B1(new_n873), .B2(new_n597), .ZN(G295));
  OAI21_X1  g449(.A(new_n859), .B1(new_n873), .B2(new_n597), .ZN(G331));
  INV_X1    g450(.A(new_n865), .ZN(new_n876));
  XOR2_X1   g451(.A(G171), .B(G286), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n822), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n869), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT110), .ZN(new_n881));
  INV_X1    g456(.A(new_n871), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(new_n878), .ZN(new_n883));
  INV_X1    g458(.A(new_n878), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(KEYINPUT110), .A3(new_n871), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n876), .A2(new_n880), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n880), .B1(new_n882), .B2(new_n878), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n865), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n829), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT111), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n886), .A2(KEYINPUT111), .A3(new_n829), .A4(new_n888), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(KEYINPUT43), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n883), .A2(new_n885), .A3(new_n880), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n865), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n886), .A3(new_n829), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n893), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(KEYINPUT43), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n886), .A2(new_n899), .A3(new_n829), .A4(new_n888), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n903), .ZN(G397));
  INV_X1    g479(.A(G1384), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT45), .B1(new_n841), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(G160), .A2(G40), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT113), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n908), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT113), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n736), .B(G2067), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(G1996), .B2(new_n711), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G1996), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(new_n711), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT114), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n911), .A2(new_n779), .A3(new_n776), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n911), .A2(G1986), .A3(G290), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT112), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT114), .ZN(new_n927));
  OAI221_X1 g502(.A(new_n927), .B1(new_n711), .B2(new_n920), .C1(new_n915), .C2(new_n917), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n765), .A2(new_n771), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n765), .A2(new_n771), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n914), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND4_X1   g506(.A1(new_n922), .A2(new_n926), .A3(new_n928), .A4(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT124), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n510), .A2(new_n905), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n907), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G1384), .B1(new_n505), .B2(new_n509), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT118), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT45), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n937), .B2(KEYINPUT45), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G2084), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  AOI211_X1 g520(.A(KEYINPUT50), .B(G1384), .C1(new_n505), .C2(new_n509), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n945), .A2(new_n946), .A3(new_n907), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n942), .A2(new_n689), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G8), .ZN(new_n949));
  NOR2_X1   g524(.A1(G168), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n933), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n908), .B1(new_n937), .B2(KEYINPUT45), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n510), .A2(KEYINPUT45), .A3(new_n905), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT118), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n955), .B2(new_n939), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n934), .A2(KEYINPUT50), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n937), .A2(new_n944), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n908), .A3(new_n958), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n956), .A2(G1966), .B1(new_n959), .B2(G2084), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(KEYINPUT124), .A3(new_n950), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n952), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT62), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n964), .B(G8), .C1(new_n960), .C2(G286), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT51), .B(new_n951), .C1(new_n948), .C2(new_n949), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n962), .A2(new_n963), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT45), .B(new_n905), .C1(new_n839), .C2(new_n840), .ZN(new_n968));
  INV_X1    g543(.A(G2078), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n936), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT125), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n947), .A2(G1961), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n970), .A2(KEYINPUT125), .A3(new_n971), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n956), .A2(KEYINPUT53), .A3(new_n969), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(G305), .A2(G1981), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n670), .B1(new_n579), .B2(new_n581), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT49), .ZN(new_n982));
  OR3_X1    g557(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n979), .B2(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n937), .A2(new_n908), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n981), .A2(KEYINPUT49), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n985), .A2(G8), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n750), .A2(G1976), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(G8), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT52), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n986), .A2(G8), .A3(new_n989), .A4(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n988), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT115), .B(G2090), .Z(new_n997));
  NOR2_X1   g572(.A1(new_n959), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(G1971), .B1(new_n968), .B2(new_n936), .ZN(new_n999));
  OAI21_X1  g574(.A(G8), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G166), .A2(new_n949), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT55), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(G8), .B(new_n1002), .C1(new_n998), .C2(new_n999), .ZN(new_n1005));
  AND4_X1   g580(.A1(new_n978), .A2(new_n996), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n967), .A2(new_n1006), .A3(G171), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT126), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n967), .A2(new_n1006), .A3(KEYINPUT126), .A4(G171), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n960), .A2(G8), .A3(G168), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n995), .A2(KEYINPUT117), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n988), .A2(new_n1017), .A3(new_n991), .A4(new_n994), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1004), .A2(KEYINPUT63), .A3(new_n1005), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT119), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(new_n1014), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT63), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1023), .A2(new_n1024), .A3(new_n1005), .A4(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1004), .A2(new_n996), .A3(new_n1005), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1028), .B2(new_n1014), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1021), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1022), .A2(new_n1005), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n986), .A2(G8), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n988), .A2(new_n992), .A3(new_n750), .ZN(new_n1033));
  INV_X1    g608(.A(new_n979), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1013), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n906), .A2(new_n907), .ZN(new_n1039));
  AND4_X1   g614(.A1(KEYINPUT53), .A2(new_n1039), .A3(new_n969), .A4(new_n968), .ZN(new_n1040));
  XOR2_X1   g615(.A(G171), .B(KEYINPUT54), .Z(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1042), .A2(new_n975), .A3(new_n976), .A4(new_n974), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1028), .B1(new_n1041), .B2(new_n978), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n1010), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n968), .A2(new_n936), .A3(new_n919), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n968), .A2(new_n936), .A3(KEYINPUT120), .A4(new_n919), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT58), .B(G1341), .Z(new_n1050));
  NAND2_X1  g625(.A1(new_n986), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(KEYINPUT59), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1052), .A2(new_n555), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1054), .B1(new_n1052), .B2(new_n555), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(KEYINPUT121), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n959), .A2(new_n703), .ZN(new_n1060));
  XNOR2_X1  g635(.A(G299), .B(KEYINPUT57), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n968), .A2(new_n936), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1062), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT61), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1061), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1065), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT122), .B1(new_n1059), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1056), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1058), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1052), .A2(new_n555), .A3(new_n1054), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n986), .A2(G2067), .ZN(new_n1082));
  INV_X1    g657(.A(G1348), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n959), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n604), .B1(new_n1084), .B2(KEYINPUT60), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT123), .B(new_n604), .C1(new_n1084), .C2(KEYINPUT60), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1084), .A2(KEYINPUT60), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1074), .A2(new_n1081), .A3(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1084), .A2(new_n596), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1065), .B1(new_n1093), .B2(new_n1067), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1045), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n932), .B1(new_n1038), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n922), .A2(new_n928), .A3(new_n930), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n736), .A2(G2067), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n915), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT127), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT46), .ZN(new_n1101));
  XOR2_X1   g676(.A(new_n920), .B(new_n1101), .Z(new_n1102));
  NOR2_X1   g677(.A1(new_n1100), .A2(KEYINPUT46), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n916), .A2(new_n711), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n914), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT47), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n924), .B(KEYINPUT48), .Z(new_n1109));
  AND4_X1   g684(.A1(new_n922), .A2(new_n928), .A3(new_n931), .A4(new_n1109), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1099), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1096), .A2(new_n1111), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g687(.A(new_n462), .B1(new_n898), .B2(new_n900), .ZN(new_n1114));
  AOI21_X1  g688(.A(G227), .B1(new_n636), .B2(new_n638), .ZN(new_n1115));
  INV_X1    g689(.A(G229), .ZN(new_n1116));
  NAND4_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n857), .ZN(G225));
  INV_X1    g691(.A(G225), .ZN(G308));
endmodule


