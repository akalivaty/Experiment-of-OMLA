

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765;

  INV_X1 U370 ( .A(n544), .ZN(n442) );
  INV_X2 U371 ( .A(G953), .ZN(n759) );
  NAND2_X1 U372 ( .A1(n514), .A2(n442), .ZN(n444) );
  NOR2_X1 U373 ( .A1(n712), .A2(n515), .ZN(n516) );
  XNOR2_X2 U374 ( .A(n428), .B(KEYINPUT77), .ZN(n514) );
  OR2_X2 U375 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U376 ( .A1(n739), .A2(n359), .ZN(n702) );
  NOR2_X1 U377 ( .A1(n355), .A2(n538), .ZN(n557) );
  AND2_X1 U378 ( .A1(n647), .A2(n549), .ZN(n551) );
  INV_X1 U379 ( .A(n465), .ZN(n585) );
  OR2_X1 U380 ( .A1(n654), .A2(G902), .ZN(n424) );
  XNOR2_X1 U381 ( .A(G146), .B(G125), .ZN(n452) );
  INV_X1 U382 ( .A(G143), .ZN(n390) );
  XNOR2_X1 U383 ( .A(G119), .B(G116), .ZN(n430) );
  XNOR2_X1 U384 ( .A(G146), .B(G113), .ZN(n435) );
  XNOR2_X1 U385 ( .A(n513), .B(n512), .ZN(n349) );
  XNOR2_X1 U386 ( .A(n513), .B(n512), .ZN(n387) );
  AND2_X1 U387 ( .A1(n576), .A2(n533), .ZN(n350) );
  INV_X1 U388 ( .A(n666), .ZN(n351) );
  INV_X1 U389 ( .A(n351), .ZN(n352) );
  INV_X1 U390 ( .A(n459), .ZN(n353) );
  OR2_X1 U391 ( .A1(n543), .A2(n705), .ZN(n647) );
  XNOR2_X2 U392 ( .A(n444), .B(n443), .ZN(n724) );
  XNOR2_X2 U393 ( .A(n429), .B(n409), .ZN(n751) );
  XNOR2_X2 U394 ( .A(n456), .B(n392), .ZN(n429) );
  XNOR2_X2 U395 ( .A(n505), .B(n391), .ZN(n456) );
  NOR2_X1 U396 ( .A1(n376), .A2(n699), .ZN(n375) );
  INV_X1 U397 ( .A(KEYINPUT97), .ZN(n473) );
  NAND2_X1 U398 ( .A1(n630), .A2(KEYINPUT65), .ZN(n384) );
  XNOR2_X1 U399 ( .A(n618), .B(KEYINPUT48), .ZN(n356) );
  INV_X1 U400 ( .A(n595), .ZN(n365) );
  XNOR2_X1 U401 ( .A(n361), .B(n429), .ZN(n648) );
  XNOR2_X1 U402 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n577) );
  NOR2_X1 U403 ( .A1(n719), .A2(n718), .ZN(n572) );
  INV_X1 U404 ( .A(KEYINPUT44), .ZN(n386) );
  INV_X1 U405 ( .A(KEYINPUT4), .ZN(n391) );
  NAND2_X1 U406 ( .A1(n716), .A2(n369), .ZN(n719) );
  INV_X1 U407 ( .A(KEYINPUT106), .ZN(n565) );
  NOR2_X1 U408 ( .A1(n383), .A2(n381), .ZN(n380) );
  OR2_X1 U409 ( .A1(n630), .A2(KEYINPUT65), .ZN(n382) );
  XNOR2_X1 U410 ( .A(n362), .B(KEYINPUT39), .ZN(n619) );
  OR2_X1 U411 ( .A1(n593), .A2(n363), .ZN(n362) );
  NAND2_X1 U412 ( .A1(n364), .A2(n716), .ZN(n363) );
  NOR2_X1 U413 ( .A1(n592), .A2(n365), .ZN(n364) );
  BUF_X1 U414 ( .A(n526), .Z(n515) );
  BUF_X1 U415 ( .A(n561), .Z(n626) );
  XNOR2_X1 U416 ( .A(n368), .B(KEYINPUT30), .ZN(n593) );
  NAND2_X1 U417 ( .A1(n370), .A2(n369), .ZN(n368) );
  NAND2_X1 U418 ( .A1(n367), .A2(n366), .ZN(n592) );
  INV_X1 U419 ( .A(n519), .ZN(n367) );
  NAND2_X1 U420 ( .A1(n648), .A2(n497), .ZN(n360) );
  XNOR2_X1 U421 ( .A(KEYINPUT42), .B(n580), .ZN(n764) );
  OR2_X1 U422 ( .A1(n764), .A2(n377), .ZN(n354) );
  NOR2_X1 U423 ( .A1(n349), .A2(n386), .ZN(n355) );
  INV_X1 U424 ( .A(n359), .ZN(n758) );
  NAND2_X1 U425 ( .A1(n356), .A2(n628), .ZN(n359) );
  INV_X1 U426 ( .A(n518), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n570), .B(n569), .ZN(n763) );
  INV_X1 U428 ( .A(n620), .ZN(n369) );
  INV_X1 U429 ( .A(n582), .ZN(n377) );
  XNOR2_X1 U430 ( .A(n581), .B(KEYINPUT64), .ZN(n582) );
  AND2_X1 U431 ( .A1(n374), .A2(n375), .ZN(n617) );
  NAND2_X1 U432 ( .A1(n373), .A2(n354), .ZN(n372) );
  NAND2_X1 U433 ( .A1(n357), .A2(n382), .ZN(n381) );
  NAND2_X1 U434 ( .A1(n359), .A2(n358), .ZN(n357) );
  INV_X1 U435 ( .A(n384), .ZN(n358) );
  XNOR2_X2 U436 ( .A(n360), .B(G472), .ZN(n540) );
  XNOR2_X1 U437 ( .A(n440), .B(n433), .ZN(n361) );
  INV_X1 U438 ( .A(n576), .ZN(n370) );
  NAND2_X1 U439 ( .A1(n372), .A2(n371), .ZN(n374) );
  NAND2_X1 U440 ( .A1(n763), .A2(n582), .ZN(n371) );
  INV_X1 U441 ( .A(n763), .ZN(n373) );
  AND2_X1 U442 ( .A1(n764), .A2(n377), .ZN(n376) );
  XNOR2_X2 U443 ( .A(n390), .B(G128), .ZN(n505) );
  NOR2_X2 U444 ( .A1(n385), .A2(n384), .ZN(n383) );
  XNOR2_X2 U445 ( .A(n560), .B(KEYINPUT87), .ZN(n385) );
  NAND2_X1 U446 ( .A1(n380), .A2(n378), .ZN(n635) );
  NAND2_X1 U447 ( .A1(n385), .A2(n379), .ZN(n378) );
  AND2_X1 U448 ( .A1(n758), .A2(n631), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n387), .B(KEYINPUT44), .ZN(n550) );
  XNOR2_X1 U450 ( .A(n349), .B(G122), .ZN(G24) );
  AND2_X1 U451 ( .A1(n529), .A2(n528), .ZN(n388) );
  OR2_X1 U452 ( .A1(G953), .A2(G237), .ZN(n389) );
  INV_X1 U453 ( .A(KEYINPUT85), .ZN(n605) );
  XNOR2_X1 U454 ( .A(n606), .B(n605), .ZN(n608) );
  INV_X1 U455 ( .A(KEYINPUT46), .ZN(n581) );
  XNOR2_X1 U456 ( .A(n474), .B(n473), .ZN(n563) );
  INV_X1 U457 ( .A(G137), .ZN(n434) );
  INV_X1 U458 ( .A(KEYINPUT65), .ZN(n631) );
  XNOR2_X1 U459 ( .A(n578), .B(n577), .ZN(n579) );
  INV_X1 U460 ( .A(KEYINPUT60), .ZN(n642) );
  XNOR2_X1 U461 ( .A(G131), .B(G134), .ZN(n392) );
  INV_X1 U462 ( .A(G140), .ZN(n393) );
  XNOR2_X1 U463 ( .A(n393), .B(G137), .ZN(n409) );
  XNOR2_X1 U464 ( .A(G101), .B(G107), .ZN(n395) );
  XNOR2_X1 U465 ( .A(G146), .B(KEYINPUT98), .ZN(n394) );
  XNOR2_X1 U466 ( .A(n395), .B(n394), .ZN(n399) );
  XNOR2_X1 U467 ( .A(G110), .B(G104), .ZN(n397) );
  NAND2_X1 U468 ( .A1(n759), .A2(G227), .ZN(n396) );
  XNOR2_X1 U469 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U470 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U471 ( .A(n751), .B(n400), .ZN(n660) );
  OR2_X2 U472 ( .A1(n660), .A2(G902), .ZN(n402) );
  INV_X1 U473 ( .A(G469), .ZN(n401) );
  XNOR2_X2 U474 ( .A(n402), .B(n401), .ZN(n517) );
  XNOR2_X1 U475 ( .A(n517), .B(KEYINPUT1), .ZN(n532) );
  NAND2_X1 U476 ( .A1(G234), .A2(n759), .ZN(n404) );
  INV_X1 U477 ( .A(KEYINPUT8), .ZN(n403) );
  XNOR2_X1 U478 ( .A(n404), .B(n403), .ZN(n500) );
  NAND2_X1 U479 ( .A1(n500), .A2(G221), .ZN(n408) );
  XNOR2_X1 U480 ( .A(KEYINPUT24), .B(KEYINPUT71), .ZN(n406) );
  XNOR2_X1 U481 ( .A(KEYINPUT86), .B(KEYINPUT99), .ZN(n405) );
  XNOR2_X1 U482 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U483 ( .A(n408), .B(n407), .ZN(n417) );
  INV_X1 U484 ( .A(n409), .ZN(n413) );
  XNOR2_X1 U485 ( .A(G119), .B(G110), .ZN(n411) );
  XNOR2_X1 U486 ( .A(G128), .B(KEYINPUT23), .ZN(n410) );
  XNOR2_X1 U487 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U488 ( .A(n413), .B(n412), .ZN(n415) );
  XNOR2_X1 U489 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n414) );
  XNOR2_X1 U490 ( .A(n452), .B(n414), .ZN(n752) );
  XNOR2_X1 U491 ( .A(n415), .B(n752), .ZN(n416) );
  XNOR2_X1 U492 ( .A(n417), .B(n416), .ZN(n654) );
  XNOR2_X1 U493 ( .A(G902), .B(KEYINPUT15), .ZN(n559) );
  NAND2_X1 U494 ( .A1(n559), .A2(G234), .ZN(n418) );
  XNOR2_X1 U495 ( .A(n418), .B(KEYINPUT20), .ZN(n425) );
  NAND2_X1 U496 ( .A1(n425), .A2(G217), .ZN(n422) );
  XOR2_X1 U497 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n420) );
  INV_X1 U498 ( .A(KEYINPUT25), .ZN(n419) );
  XNOR2_X1 U499 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U500 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X2 U501 ( .A(n424), .B(n423), .ZN(n705) );
  NAND2_X1 U502 ( .A1(G221), .A2(n425), .ZN(n427) );
  INV_X1 U503 ( .A(KEYINPUT21), .ZN(n426) );
  XNOR2_X1 U504 ( .A(n427), .B(n426), .ZN(n704) );
  XNOR2_X1 U505 ( .A(n704), .B(KEYINPUT100), .ZN(n528) );
  NAND2_X1 U506 ( .A1(n705), .A2(n528), .ZN(n519) );
  OR2_X2 U507 ( .A1(n532), .A2(n519), .ZN(n428) );
  XNOR2_X1 U508 ( .A(n430), .B(KEYINPUT3), .ZN(n432) );
  XOR2_X1 U509 ( .A(G101), .B(KEYINPUT70), .Z(n431) );
  XNOR2_X1 U510 ( .A(n432), .B(n431), .ZN(n450) );
  INV_X1 U511 ( .A(n450), .ZN(n433) );
  XNOR2_X1 U512 ( .A(KEYINPUT5), .B(KEYINPUT78), .ZN(n437) );
  XNOR2_X1 U513 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U514 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U515 ( .A(KEYINPUT79), .B(n389), .ZN(n492) );
  NAND2_X1 U516 ( .A1(n492), .A2(G210), .ZN(n438) );
  XNOR2_X1 U517 ( .A(n439), .B(n438), .ZN(n440) );
  INV_X1 U518 ( .A(G902), .ZN(n497) );
  XNOR2_X1 U519 ( .A(KEYINPUT104), .B(KEYINPUT6), .ZN(n441) );
  XNOR2_X1 U520 ( .A(n540), .B(n441), .ZN(n544) );
  XNOR2_X1 U521 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n443) );
  XNOR2_X2 U522 ( .A(G113), .B(G104), .ZN(n491) );
  XNOR2_X2 U523 ( .A(G122), .B(G107), .ZN(n502) );
  XNOR2_X1 U524 ( .A(n491), .B(n502), .ZN(n448) );
  XNOR2_X1 U525 ( .A(KEYINPUT16), .B(G110), .ZN(n446) );
  XNOR2_X1 U526 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n445) );
  XNOR2_X1 U527 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U528 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U529 ( .A(n450), .B(n449), .ZN(n745) );
  XNOR2_X1 U530 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n451) );
  XNOR2_X1 U531 ( .A(n452), .B(n451), .ZN(n455) );
  NAND2_X1 U532 ( .A1(n759), .A2(G224), .ZN(n453) );
  XNOR2_X1 U533 ( .A(n453), .B(KEYINPUT82), .ZN(n454) );
  XNOR2_X1 U534 ( .A(n455), .B(n454), .ZN(n457) );
  XNOR2_X1 U535 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U536 ( .A(n745), .B(n458), .ZN(n667) );
  INV_X1 U537 ( .A(n667), .ZN(n459) );
  NAND2_X1 U538 ( .A1(n459), .A2(n559), .ZN(n462) );
  INV_X1 U539 ( .A(G237), .ZN(n460) );
  NAND2_X1 U540 ( .A1(n497), .A2(n460), .ZN(n463) );
  NAND2_X1 U541 ( .A1(n463), .A2(G210), .ZN(n461) );
  XNOR2_X1 U542 ( .A(n462), .B(n461), .ZN(n561) );
  AND2_X1 U543 ( .A1(n463), .A2(G214), .ZN(n620) );
  OR2_X2 U544 ( .A1(n561), .A2(n620), .ZN(n465) );
  INV_X1 U545 ( .A(KEYINPUT19), .ZN(n464) );
  NAND2_X1 U546 ( .A1(n585), .A2(n464), .ZN(n467) );
  NAND2_X1 U547 ( .A1(n465), .A2(KEYINPUT19), .ZN(n466) );
  NAND2_X1 U548 ( .A1(n467), .A2(n466), .ZN(n603) );
  XOR2_X1 U549 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n469) );
  NAND2_X1 U550 ( .A1(G234), .A2(G237), .ZN(n468) );
  XNOR2_X1 U551 ( .A(n469), .B(n468), .ZN(n472) );
  NAND2_X1 U552 ( .A1(n472), .A2(G952), .ZN(n470) );
  XNOR2_X1 U553 ( .A(n470), .B(KEYINPUT94), .ZN(n730) );
  INV_X1 U554 ( .A(n730), .ZN(n471) );
  NAND2_X1 U555 ( .A1(n471), .A2(n759), .ZN(n567) );
  NAND2_X1 U556 ( .A1(n472), .A2(G902), .ZN(n474) );
  INV_X1 U557 ( .A(n563), .ZN(n477) );
  XNOR2_X1 U558 ( .A(G898), .B(KEYINPUT95), .ZN(n742) );
  NAND2_X1 U559 ( .A1(n742), .A2(G953), .ZN(n475) );
  XNOR2_X1 U560 ( .A(n475), .B(KEYINPUT96), .ZN(n746) );
  INV_X1 U561 ( .A(n746), .ZN(n476) );
  NAND2_X1 U562 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U563 ( .A1(n567), .A2(n478), .ZN(n479) );
  NAND2_X1 U564 ( .A1(n603), .A2(n479), .ZN(n480) );
  XNOR2_X1 U565 ( .A(n480), .B(KEYINPUT0), .ZN(n526) );
  INV_X1 U566 ( .A(n515), .ZN(n521) );
  NAND2_X1 U567 ( .A1(n724), .A2(n521), .ZN(n483) );
  XOR2_X1 U568 ( .A(KEYINPUT83), .B(KEYINPUT34), .Z(n481) );
  XNOR2_X1 U569 ( .A(n481), .B(KEYINPUT73), .ZN(n482) );
  XNOR2_X1 U570 ( .A(n483), .B(n482), .ZN(n511) );
  XOR2_X1 U571 ( .A(KEYINPUT12), .B(G140), .Z(n485) );
  XNOR2_X1 U572 ( .A(G143), .B(G122), .ZN(n484) );
  XNOR2_X1 U573 ( .A(n485), .B(n484), .ZN(n489) );
  XOR2_X1 U574 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n487) );
  XNOR2_X1 U575 ( .A(G131), .B(KEYINPUT101), .ZN(n486) );
  XNOR2_X1 U576 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U577 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U578 ( .A(n490), .B(n752), .ZN(n496) );
  XNOR2_X1 U579 ( .A(n491), .B(KEYINPUT103), .ZN(n494) );
  NAND2_X1 U580 ( .A1(n492), .A2(G214), .ZN(n493) );
  XNOR2_X1 U581 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U582 ( .A(n496), .B(n495), .ZN(n637) );
  NAND2_X1 U583 ( .A1(n637), .A2(n497), .ZN(n499) );
  XOR2_X1 U584 ( .A(KEYINPUT13), .B(G475), .Z(n498) );
  XNOR2_X1 U585 ( .A(n499), .B(n498), .ZN(n527) );
  INV_X1 U586 ( .A(n527), .ZN(n597) );
  NAND2_X1 U587 ( .A1(n500), .A2(G217), .ZN(n504) );
  XNOR2_X1 U588 ( .A(G134), .B(KEYINPUT7), .ZN(n501) );
  XNOR2_X1 U589 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U590 ( .A(n504), .B(n503), .ZN(n508) );
  XOR2_X1 U591 ( .A(G116), .B(KEYINPUT9), .Z(n506) );
  XNOR2_X1 U592 ( .A(n505), .B(n506), .ZN(n507) );
  XNOR2_X1 U593 ( .A(n508), .B(n507), .ZN(n657) );
  OR2_X1 U594 ( .A1(n657), .A2(G902), .ZN(n509) );
  XNOR2_X1 U595 ( .A(n509), .B(G478), .ZN(n594) );
  INV_X1 U596 ( .A(n594), .ZN(n522) );
  NOR2_X1 U597 ( .A1(n597), .A2(n522), .ZN(n510) );
  NAND2_X1 U598 ( .A1(n511), .A2(n510), .ZN(n513) );
  XOR2_X1 U599 ( .A(KEYINPUT88), .B(KEYINPUT35), .Z(n512) );
  NAND2_X1 U600 ( .A1(n514), .A2(n540), .ZN(n712) );
  XNOR2_X1 U601 ( .A(n516), .B(KEYINPUT31), .ZN(n695) );
  BUF_X1 U602 ( .A(n517), .Z(n518) );
  NOR2_X1 U603 ( .A1(n592), .A2(n540), .ZN(n520) );
  NAND2_X1 U604 ( .A1(n521), .A2(n520), .ZN(n678) );
  AND2_X1 U605 ( .A1(n695), .A2(n678), .ZN(n523) );
  NAND2_X1 U606 ( .A1(n527), .A2(n522), .ZN(n692) );
  OR2_X1 U607 ( .A1(n527), .A2(n522), .ZN(n696) );
  AND2_X1 U608 ( .A1(n692), .A2(n696), .ZN(n720) );
  NOR2_X1 U609 ( .A1(n523), .A2(n720), .ZN(n525) );
  NOR2_X1 U610 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n524) );
  NOR2_X1 U611 ( .A1(n525), .A2(n524), .ZN(n537) );
  INV_X1 U612 ( .A(n526), .ZN(n530) );
  OR2_X1 U613 ( .A1(n527), .A2(n594), .ZN(n718) );
  INV_X1 U614 ( .A(n718), .ZN(n529) );
  NAND2_X1 U615 ( .A1(n530), .A2(n388), .ZN(n531) );
  XNOR2_X1 U616 ( .A(n531), .B(KEYINPUT22), .ZN(n547) );
  INV_X1 U617 ( .A(n547), .ZN(n534) );
  BUF_X1 U618 ( .A(n532), .Z(n533) );
  INV_X1 U619 ( .A(n533), .ZN(n590) );
  NAND2_X1 U620 ( .A1(n534), .A2(n533), .ZN(n539) );
  NOR2_X1 U621 ( .A1(n539), .A2(n442), .ZN(n535) );
  XOR2_X1 U622 ( .A(KEYINPUT89), .B(n535), .Z(n536) );
  NAND2_X1 U623 ( .A1(n536), .A2(n705), .ZN(n646) );
  NAND2_X1 U624 ( .A1(n537), .A2(n646), .ZN(n538) );
  XNOR2_X1 U625 ( .A(n540), .B(KEYINPUT105), .ZN(n576) );
  NAND2_X1 U626 ( .A1(n350), .A2(n534), .ZN(n542) );
  INV_X1 U627 ( .A(KEYINPUT67), .ZN(n541) );
  XNOR2_X1 U628 ( .A(n542), .B(n541), .ZN(n543) );
  INV_X1 U629 ( .A(n705), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n544), .A2(n573), .ZN(n545) );
  OR2_X1 U631 ( .A1(n545), .A2(n533), .ZN(n546) );
  XNOR2_X1 U632 ( .A(n548), .B(KEYINPUT32), .ZN(n645) );
  AND2_X1 U633 ( .A1(KEYINPUT66), .A2(n645), .ZN(n549) );
  NAND2_X1 U634 ( .A1(n550), .A2(n551), .ZN(n555) );
  NAND2_X1 U635 ( .A1(n647), .A2(n645), .ZN(n553) );
  NAND2_X1 U636 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n552) );
  NAND2_X1 U637 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U638 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U639 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U640 ( .A(n558), .B(KEYINPUT45), .ZN(n632) );
  INV_X1 U641 ( .A(n559), .ZN(n629) );
  NAND2_X1 U642 ( .A1(n632), .A2(n629), .ZN(n560) );
  XNOR2_X1 U643 ( .A(KEYINPUT76), .B(KEYINPUT38), .ZN(n562) );
  XNOR2_X1 U644 ( .A(n626), .B(n562), .ZN(n716) );
  OR2_X1 U645 ( .A1(n759), .A2(n563), .ZN(n564) );
  NOR2_X1 U646 ( .A1(G900), .A2(n564), .ZN(n566) );
  XNOR2_X1 U647 ( .A(n566), .B(n565), .ZN(n568) );
  NAND2_X1 U648 ( .A1(n568), .A2(n567), .ZN(n595) );
  INV_X1 U649 ( .A(n692), .ZN(n687) );
  NAND2_X1 U650 ( .A1(n619), .A2(n687), .ZN(n570) );
  INV_X1 U651 ( .A(KEYINPUT40), .ZN(n569) );
  XNOR2_X1 U652 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n571) );
  XNOR2_X1 U653 ( .A(n572), .B(n571), .ZN(n732) );
  AND2_X1 U654 ( .A1(n595), .A2(n704), .ZN(n574) );
  NAND2_X1 U655 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U656 ( .A(n575), .B(KEYINPUT69), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n583), .A2(n370), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n579), .A2(n366), .ZN(n602) );
  NOR2_X1 U659 ( .A1(n732), .A2(n602), .ZN(n580) );
  AND2_X1 U660 ( .A1(n583), .A2(n687), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n584), .A2(n442), .ZN(n621) );
  XNOR2_X1 U662 ( .A(n621), .B(KEYINPUT111), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n586), .A2(n585), .ZN(n589) );
  INV_X1 U664 ( .A(KEYINPUT90), .ZN(n587) );
  XNOR2_X1 U665 ( .A(n587), .B(KEYINPUT36), .ZN(n588) );
  XNOR2_X1 U666 ( .A(n589), .B(n588), .ZN(n591) );
  AND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n699) );
  OR2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n599) );
  INV_X1 U671 ( .A(n626), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n686) );
  INV_X1 U674 ( .A(n602), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n611) );
  NAND2_X1 U676 ( .A1(n611), .A2(KEYINPUT47), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n720), .A2(KEYINPUT47), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U679 ( .A1(n686), .A2(n609), .ZN(n610) );
  XOR2_X1 U680 ( .A(n610), .B(KEYINPUT84), .Z(n615) );
  INV_X1 U681 ( .A(n611), .ZN(n688) );
  INV_X1 U682 ( .A(n720), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n688), .A2(n612), .ZN(n613) );
  NOR2_X1 U684 ( .A1(KEYINPUT47), .A2(n613), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n616) );
  AND2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n618) );
  INV_X1 U687 ( .A(n696), .ZN(n683) );
  NAND2_X1 U688 ( .A1(n683), .A2(n619), .ZN(n701) );
  NOR2_X1 U689 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n622), .A2(n533), .ZN(n625) );
  XNOR2_X1 U691 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n623) );
  XOR2_X1 U692 ( .A(n623), .B(KEYINPUT107), .Z(n624) );
  XNOR2_X1 U693 ( .A(n625), .B(n624), .ZN(n627) );
  NAND2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n644) );
  AND2_X1 U695 ( .A1(n701), .A2(n644), .ZN(n628) );
  NAND2_X1 U696 ( .A1(n629), .A2(KEYINPUT2), .ZN(n630) );
  BUF_X1 U697 ( .A(n632), .Z(n633) );
  INV_X1 U698 ( .A(n633), .ZN(n739) );
  NAND2_X1 U699 ( .A1(n702), .A2(KEYINPUT2), .ZN(n634) );
  AND2_X2 U700 ( .A1(n635), .A2(n634), .ZN(n666) );
  NAND2_X1 U701 ( .A1(n666), .A2(G475), .ZN(n639) );
  XOR2_X1 U702 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n636) );
  XNOR2_X1 U703 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U704 ( .A(n639), .B(n638), .ZN(n641) );
  INV_X1 U705 ( .A(G952), .ZN(n640) );
  NAND2_X1 U706 ( .A1(n640), .A2(G953), .ZN(n672) );
  NAND2_X1 U707 ( .A1(n641), .A2(n672), .ZN(n643) );
  XNOR2_X1 U708 ( .A(n643), .B(n642), .ZN(G60) );
  XNOR2_X1 U709 ( .A(n644), .B(G140), .ZN(G42) );
  XNOR2_X1 U710 ( .A(n645), .B(G119), .ZN(G21) );
  XNOR2_X1 U711 ( .A(n646), .B(G101), .ZN(G3) );
  XNOR2_X1 U712 ( .A(n647), .B(G110), .ZN(G12) );
  NAND2_X1 U713 ( .A1(n666), .A2(G472), .ZN(n650) );
  XNOR2_X1 U714 ( .A(n648), .B(KEYINPUT62), .ZN(n649) );
  XNOR2_X1 U715 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U716 ( .A1(n651), .A2(n672), .ZN(n653) );
  XOR2_X1 U717 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n652) );
  XNOR2_X1 U718 ( .A(n653), .B(n652), .ZN(G57) );
  NAND2_X1 U719 ( .A1(n352), .A2(G217), .ZN(n655) );
  XNOR2_X1 U720 ( .A(n655), .B(n654), .ZN(n656) );
  INV_X1 U721 ( .A(n672), .ZN(n664) );
  NOR2_X1 U722 ( .A1(n656), .A2(n664), .ZN(G66) );
  NAND2_X1 U723 ( .A1(n352), .A2(G478), .ZN(n658) );
  XNOR2_X1 U724 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X1 U725 ( .A1(n659), .A2(n664), .ZN(G63) );
  NAND2_X1 U726 ( .A1(n352), .A2(G469), .ZN(n663) );
  XOR2_X1 U727 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n661) );
  XNOR2_X1 U728 ( .A(n660), .B(n661), .ZN(n662) );
  XNOR2_X1 U729 ( .A(n663), .B(n662), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n665), .A2(n664), .ZN(G54) );
  NAND2_X1 U731 ( .A1(n666), .A2(G210), .ZN(n671) );
  XNOR2_X1 U732 ( .A(KEYINPUT92), .B(KEYINPUT54), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n668), .B(KEYINPUT55), .ZN(n669) );
  XNOR2_X1 U734 ( .A(n353), .B(n669), .ZN(n670) );
  XNOR2_X1 U735 ( .A(n671), .B(n670), .ZN(n673) );
  NAND2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n675) );
  XNOR2_X1 U737 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n674) );
  XNOR2_X1 U738 ( .A(n675), .B(n674), .ZN(G51) );
  NOR2_X1 U739 ( .A1(n692), .A2(n678), .ZN(n676) );
  XOR2_X1 U740 ( .A(KEYINPUT112), .B(n676), .Z(n677) );
  XNOR2_X1 U741 ( .A(G104), .B(n677), .ZN(G6) );
  NOR2_X1 U742 ( .A1(n678), .A2(n696), .ZN(n682) );
  XOR2_X1 U743 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n680) );
  XNOR2_X1 U744 ( .A(G107), .B(KEYINPUT27), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n682), .B(n681), .ZN(G9) );
  XOR2_X1 U747 ( .A(G128), .B(KEYINPUT29), .Z(n685) );
  NAND2_X1 U748 ( .A1(n688), .A2(n683), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n685), .B(n684), .ZN(G30) );
  XOR2_X1 U750 ( .A(G143), .B(n686), .Z(G45) );
  XOR2_X1 U751 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n690) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U753 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U754 ( .A(G146), .B(n691), .ZN(G48) );
  NOR2_X1 U755 ( .A1(n692), .A2(n695), .ZN(n693) );
  XOR2_X1 U756 ( .A(KEYINPUT116), .B(n693), .Z(n694) );
  XNOR2_X1 U757 ( .A(G113), .B(n694), .ZN(G15) );
  NOR2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U759 ( .A(G116), .B(KEYINPUT117), .ZN(n697) );
  XNOR2_X1 U760 ( .A(n698), .B(n697), .ZN(G18) );
  XNOR2_X1 U761 ( .A(n699), .B(G125), .ZN(n700) );
  XNOR2_X1 U762 ( .A(n700), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U763 ( .A(G134), .B(n701), .ZN(G36) );
  XOR2_X1 U764 ( .A(KEYINPUT2), .B(n702), .Z(n736) );
  NAND2_X1 U765 ( .A1(n533), .A2(n519), .ZN(n703) );
  XNOR2_X1 U766 ( .A(n703), .B(KEYINPUT50), .ZN(n710) );
  XNOR2_X1 U767 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n707) );
  NOR2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U769 ( .A(n707), .B(n706), .Z(n708) );
  NOR2_X1 U770 ( .A1(n708), .A2(n540), .ZN(n709) );
  NAND2_X1 U771 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U772 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U773 ( .A(n713), .B(KEYINPUT119), .ZN(n714) );
  XOR2_X1 U774 ( .A(KEYINPUT51), .B(n714), .Z(n715) );
  NOR2_X1 U775 ( .A1(n732), .A2(n715), .ZN(n727) );
  NOR2_X1 U776 ( .A1(n716), .A2(n369), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U780 ( .A(n723), .B(KEYINPUT120), .ZN(n725) );
  INV_X1 U781 ( .A(n724), .ZN(n731) );
  NOR2_X1 U782 ( .A1(n725), .A2(n731), .ZN(n726) );
  NOR2_X1 U783 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n728), .B(KEYINPUT52), .ZN(n729) );
  NOR2_X1 U785 ( .A1(n730), .A2(n729), .ZN(n734) );
  NOR2_X1 U786 ( .A1(n732), .A2(n731), .ZN(n733) );
  OR2_X1 U787 ( .A1(n734), .A2(n733), .ZN(n735) );
  OR2_X1 U788 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U789 ( .A1(n737), .A2(G953), .ZN(n738) );
  XNOR2_X1 U790 ( .A(n738), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U791 ( .A1(n739), .A2(G953), .ZN(n744) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n740) );
  XOR2_X1 U793 ( .A(KEYINPUT61), .B(n740), .Z(n741) );
  NOR2_X1 U794 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U795 ( .A1(n744), .A2(n743), .ZN(n750) );
  XNOR2_X1 U796 ( .A(n745), .B(KEYINPUT123), .ZN(n747) );
  NAND2_X1 U797 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U798 ( .A(n748), .B(KEYINPUT124), .ZN(n749) );
  XNOR2_X1 U799 ( .A(n750), .B(n749), .ZN(G69) );
  XNOR2_X1 U800 ( .A(n752), .B(KEYINPUT125), .ZN(n753) );
  XNOR2_X1 U801 ( .A(n751), .B(n753), .ZN(n757) );
  XOR2_X1 U802 ( .A(KEYINPUT126), .B(n757), .Z(n754) );
  XNOR2_X1 U803 ( .A(G227), .B(n754), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n756), .A2(G953), .ZN(n762) );
  XNOR2_X1 U806 ( .A(n758), .B(n757), .ZN(n760) );
  NAND2_X1 U807 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U808 ( .A1(n762), .A2(n761), .ZN(G72) );
  XOR2_X1 U809 ( .A(G131), .B(n763), .Z(G33) );
  XNOR2_X1 U810 ( .A(G137), .B(KEYINPUT127), .ZN(n765) );
  XNOR2_X1 U811 ( .A(n765), .B(n764), .ZN(G39) );
endmodule

