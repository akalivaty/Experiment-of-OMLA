//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032;
  NAND2_X1  g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT103), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT103), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT104), .B(G92gat), .ZN(new_n209));
  INV_X1    g008(.A(G85gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n209), .A2(new_n210), .B1(KEYINPUT8), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n207), .A2(new_n208), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G99gat), .B(G106gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n207), .A2(new_n212), .A3(new_n214), .A4(new_n208), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT9), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(G57gat), .A2(G64gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G57gat), .A2(G64gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G71gat), .A2(G78gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT98), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n219), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT98), .A2(G71gat), .A3(G78gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n225), .A2(KEYINPUT9), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n219), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n222), .A2(KEYINPUT99), .A3(new_n223), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT99), .B1(new_n222), .B2(new_n223), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT100), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G57gat), .B(G64gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT99), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n233), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT100), .A3(new_n232), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n230), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT101), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI211_X1 g045(.A(KEYINPUT101), .B(new_n230), .C1(new_n238), .C2(new_n243), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n218), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n218), .A2(new_n244), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT10), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n236), .A2(new_n237), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT100), .B1(new_n242), .B2(new_n232), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n229), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT101), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n244), .A2(new_n245), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT10), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n218), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT105), .B1(new_n251), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT105), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n249), .B1(new_n257), .B2(new_n218), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n263), .B(new_n260), .C1(new_n264), .C2(KEYINPUT10), .ZN(new_n265));
  NAND2_X1  g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G120gat), .B(G148gat), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT107), .ZN(new_n270));
  XNOR2_X1  g069(.A(G176gat), .B(G204gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n274), .B2(KEYINPUT106), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n274), .A2(KEYINPUT106), .ZN(new_n276));
  OR3_X1    g075(.A1(new_n268), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n272), .B(KEYINPUT108), .Z(new_n278));
  NAND2_X1  g077(.A1(new_n248), .A2(new_n250), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n258), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n273), .B1(new_n280), .B2(new_n260), .ZN(new_n281));
  INV_X1    g080(.A(new_n274), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n218), .ZN(new_n286));
  XNOR2_X1  g085(.A(G43gat), .B(G50gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT15), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n288), .A2(new_n289), .B1(G29gat), .B2(G36gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(KEYINPUT15), .ZN(new_n291));
  OR3_X1    g090(.A1(KEYINPUT93), .A2(G29gat), .A3(G36gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT93), .B1(G29gat), .B2(G36gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(KEYINPUT14), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT14), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n295), .B(KEYINPUT93), .C1(G29gat), .C2(G36gat), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n290), .A2(new_n291), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n291), .ZN(new_n298));
  INV_X1    g097(.A(G29gat), .ZN(new_n299));
  INV_X1    g098(.A(G36gat), .ZN(new_n300));
  OAI221_X1 g099(.A(new_n296), .B1(new_n299), .B2(new_n300), .C1(new_n287), .C2(KEYINPUT15), .ZN(new_n301));
  INV_X1    g100(.A(new_n294), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(G232gat), .A2(G233gat), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n286), .A2(new_n304), .B1(KEYINPUT41), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT17), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n297), .A2(new_n303), .A3(KEYINPUT17), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n218), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G190gat), .B(G218gat), .Z(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n305), .A2(KEYINPUT41), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n314), .B(KEYINPUT102), .Z(new_n315));
  XNOR2_X1  g114(.A(G134gat), .B(G162gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n311), .A2(new_n312), .ZN(new_n319));
  OR3_X1    g118(.A1(new_n313), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n313), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n257), .A2(KEYINPUT21), .ZN(new_n324));
  NAND2_X1  g123(.A1(G231gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n324), .B(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G127gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n324), .B(new_n325), .ZN(new_n329));
  INV_X1    g128(.A(G127gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G15gat), .B(G22gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT16), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(G1gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(G1gat), .B2(new_n333), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G8gat), .ZN(new_n337));
  INV_X1    g136(.A(G8gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n335), .B(new_n338), .C1(G1gat), .C2(new_n333), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n257), .B2(KEYINPUT21), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n331), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n345));
  INV_X1    g144(.A(G155gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G183gat), .B(G211gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  AND3_X1   g148(.A1(new_n342), .A2(new_n344), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n342), .B2(new_n344), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n285), .B(new_n323), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n308), .A2(new_n337), .A3(new_n339), .A4(new_n309), .ZN(new_n353));
  NAND2_X1  g152(.A1(G229gat), .A2(G233gat), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n303), .A2(new_n297), .B1(new_n337), .B2(new_n339), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT18), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G113gat), .B(G141gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G197gat), .ZN(new_n361));
  XOR2_X1   g160(.A(KEYINPUT11), .B(G169gat), .Z(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT12), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n353), .A2(KEYINPUT18), .A3(new_n354), .A4(new_n356), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n354), .B(KEYINPUT13), .Z(new_n367));
  NOR2_X1   g166(.A1(new_n304), .A2(new_n340), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(new_n355), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT95), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(KEYINPUT95), .B(new_n367), .C1(new_n368), .C2(new_n355), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n366), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT96), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n366), .A2(new_n371), .A3(KEYINPUT96), .A4(new_n372), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT94), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n357), .A2(KEYINPUT94), .A3(new_n358), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n376), .A2(new_n377), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n364), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n374), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT35), .ZN(new_n386));
  INV_X1    g185(.A(G141gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G148gat), .ZN(new_n388));
  INV_X1    g187(.A(G148gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G141gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n393));
  INV_X1    g192(.A(G162gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n346), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT2), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT80), .B(G162gat), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(G155gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(G141gat), .B(G148gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT2), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n346), .A2(new_n394), .A3(KEYINPUT78), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(G155gat), .B2(G162gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n406), .A3(new_n396), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n398), .A2(new_n401), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT3), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n410));
  OAI221_X1 g209(.A(new_n410), .B1(new_n403), .B2(new_n407), .C1(new_n398), .C2(new_n401), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n330), .A2(G134gat), .ZN(new_n412));
  INV_X1    g211(.A(G134gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(G127gat), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT69), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(G127gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n330), .A2(G134gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT69), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT1), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(G113gat), .B2(G120gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(G113gat), .A2(G120gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n415), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(G113gat), .A2(G120gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(new_n420), .A3(new_n422), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n427), .A2(new_n418), .A3(new_n416), .A4(new_n417), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n411), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n429), .B2(new_n408), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n392), .A2(new_n397), .A3(new_n393), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n400), .A2(G155gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT2), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n402), .A2(KEYINPUT2), .ZN(new_n437));
  INV_X1    g236(.A(new_n407), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n434), .A2(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n425), .A2(new_n428), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT4), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n430), .A2(new_n431), .A3(new_n433), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT5), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n440), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n408), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n431), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n429), .A2(new_n408), .A3(new_n432), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT4), .B1(new_n439), .B2(new_n440), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n450), .A2(KEYINPUT5), .A3(new_n431), .A4(new_n430), .ZN(new_n451));
  XNOR2_X1  g250(.A(G1gat), .B(G29gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT0), .ZN(new_n453));
  XNOR2_X1  g252(.A(G57gat), .B(G85gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n447), .A2(new_n451), .A3(KEYINPUT6), .A4(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT82), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n447), .A2(new_n451), .ZN(new_n459));
  INV_X1    g258(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n451), .A3(new_n455), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(G169gat), .A2(G176gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT26), .ZN(new_n467));
  NAND2_X1  g266(.A1(G183gat), .A2(G190gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G169gat), .A2(G176gat), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT26), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(new_n466), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n476));
  INV_X1    g275(.A(G183gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT27), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT27), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G183gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n476), .A2(new_n478), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT67), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(KEYINPUT67), .A3(new_n483), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n478), .A2(new_n480), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n481), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT68), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT28), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n475), .B1(new_n488), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n466), .A2(KEYINPUT23), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(G169gat), .B2(G176gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n470), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n476), .A2(new_n477), .A3(new_n481), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT24), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n468), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT64), .ZN(new_n506));
  NAND3_X1  g305(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT64), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n468), .A2(new_n508), .A3(new_n504), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n503), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(G183gat), .A2(G190gat), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n505), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n501), .B1(new_n513), .B2(new_n500), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n440), .B1(new_n496), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n482), .A2(KEYINPUT67), .A3(new_n483), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT67), .B1(new_n482), .B2(new_n483), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n495), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n474), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(new_n429), .A3(new_n515), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n517), .A2(G227gat), .A3(new_n522), .A4(G233gat), .ZN(new_n523));
  XOR2_X1   g322(.A(G71gat), .B(G99gat), .Z(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G43gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT33), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(KEYINPUT32), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n523), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n527), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n523), .A2(KEYINPUT32), .ZN(new_n533));
  INV_X1    g332(.A(new_n523), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n533), .B(new_n526), .C1(new_n534), .C2(KEYINPUT33), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n517), .A2(new_n522), .B1(G227gat), .B2(G233gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT34), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n535), .A3(new_n538), .ZN(new_n541));
  AND4_X1   g340(.A1(new_n386), .A2(new_n465), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(G8gat), .B(G36gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT75), .ZN(new_n544));
  XNOR2_X1  g343(.A(G64gat), .B(G92gat), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n544), .B(new_n545), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G226gat), .A2(G233gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n496), .B2(new_n516), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n521), .A2(KEYINPUT74), .A3(new_n515), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G211gat), .B(G218gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G211gat), .A2(G218gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT22), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(G197gat), .A2(G204gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(G197gat), .A2(G204gat), .ZN(new_n559));
  OAI22_X1  g358(.A1(new_n557), .A2(KEYINPUT71), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n554), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT72), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n557), .A2(KEYINPUT71), .ZN(new_n566));
  XNOR2_X1  g365(.A(G197gat), .B(G204gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n562), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n566), .A2(new_n553), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(KEYINPUT72), .B(new_n554), .C1(new_n560), .C2(new_n563), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n570), .A2(KEYINPUT73), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT73), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n521), .A2(new_n515), .ZN(new_n576));
  INV_X1    g375(.A(new_n548), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT29), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n552), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n550), .A2(new_n578), .A3(new_n551), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n521), .A2(new_n577), .A3(new_n515), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n574), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(KEYINPUT30), .B(new_n547), .C1(new_n580), .C2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(new_n582), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n575), .ZN(new_n588));
  INV_X1    g387(.A(new_n551), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT74), .B1(new_n521), .B2(new_n515), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n577), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n579), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n574), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n594), .A2(KEYINPUT76), .A3(KEYINPUT30), .A4(new_n547), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n593), .A3(new_n546), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT77), .B(KEYINPUT30), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n547), .B1(new_n580), .B2(new_n583), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n596), .A2(KEYINPUT89), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT89), .B1(new_n596), .B2(new_n601), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n542), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n570), .A2(new_n605), .A3(new_n408), .A4(new_n571), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n409), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT85), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n411), .A2(new_n605), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n572), .B2(new_n573), .ZN(new_n611));
  NAND2_X1  g410(.A1(G228gat), .A2(G233gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n606), .A2(KEYINPUT85), .A3(new_n409), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n609), .A2(new_n611), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n612), .B(KEYINPUT83), .Z(new_n616));
  AOI21_X1  g415(.A(KEYINPUT29), .B1(new_n439), .B2(new_n410), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT73), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n569), .A2(new_n565), .ZN(new_n619));
  INV_X1    g418(.A(new_n559), .ZN(new_n620));
  NAND2_X1  g419(.A1(G197gat), .A2(G204gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n620), .A2(new_n621), .B1(new_n561), .B2(new_n562), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n553), .B1(new_n622), .B2(new_n566), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n571), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n618), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n570), .A2(KEYINPUT73), .A3(new_n571), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n617), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n564), .A2(KEYINPUT84), .A3(new_n569), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT84), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n631), .A3(new_n605), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n439), .B1(new_n632), .B2(new_n410), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n616), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n615), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(G22gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G78gat), .B(G106gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT31), .B(G50gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G22gat), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n615), .A2(new_n634), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n636), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT86), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n636), .A2(new_n643), .A3(new_n641), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n640), .B1(new_n615), .B2(new_n634), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n639), .B1(new_n645), .B2(KEYINPUT86), .ZN(new_n646));
  AOI22_X1  g445(.A1(KEYINPUT87), .A2(new_n642), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT87), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n636), .A2(new_n648), .A3(new_n639), .A4(new_n641), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT88), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n642), .A2(KEYINPUT87), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT88), .A4(new_n649), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n385), .B1(new_n604), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n465), .A2(new_n540), .A3(new_n386), .A4(new_n541), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n546), .B1(new_n588), .B2(new_n593), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT76), .B1(new_n658), .B2(KEYINPUT30), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n584), .A2(new_n585), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n601), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT89), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n586), .A2(new_n595), .B1(new_n599), .B2(new_n600), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT89), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n657), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n652), .A3(new_n649), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT88), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n653), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(KEYINPUT92), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n463), .A2(new_n462), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n455), .B1(new_n447), .B2(new_n451), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT81), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT81), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n461), .A2(new_n675), .A3(new_n462), .A4(new_n463), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n458), .ZN(new_n678));
  INV_X1    g477(.A(new_n540), .ZN(new_n679));
  INV_X1    g478(.A(new_n541), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n670), .A2(new_n678), .A3(new_n664), .A4(new_n681), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n656), .A2(new_n671), .B1(KEYINPUT35), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT37), .B1(new_n588), .B2(new_n593), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(new_n547), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT37), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n594), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT38), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT38), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n581), .A2(new_n574), .A3(new_n582), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT37), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n574), .B1(new_n591), .B2(new_n592), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n693), .A2(new_n684), .A3(new_n547), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n456), .A2(KEYINPUT82), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n456), .A2(KEYINPUT82), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n464), .A2(new_n695), .A3(new_n696), .A4(new_n600), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n669), .A2(new_n653), .B1(new_n688), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT39), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n430), .A2(new_n433), .A3(new_n441), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT90), .ZN(new_n702));
  INV_X1    g501(.A(new_n431), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n701), .B2(new_n703), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n700), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n706), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n444), .A2(new_n445), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n700), .B1(new_n709), .B2(new_n431), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n704), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n707), .A2(new_n711), .A3(new_n460), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT40), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(KEYINPUT91), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n463), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n712), .B2(KEYINPUT91), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n663), .A2(new_n665), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n699), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n664), .A2(new_n678), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n669), .A2(new_n720), .A3(new_n653), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n681), .A2(KEYINPUT36), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT36), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n679), .B2(new_n680), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n719), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n384), .B1(new_n683), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT97), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT97), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n730), .B(new_n384), .C1(new_n683), .C2(new_n727), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n352), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n678), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g534(.A1(new_n663), .A2(new_n665), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT16), .B(G8gat), .Z(new_n738));
  AND3_X1   g537(.A1(new_n732), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n338), .B1(new_n732), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT42), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT42), .B2(new_n739), .ZN(G1325gat));
  NAND2_X1  g541(.A1(new_n729), .A2(new_n731), .ZN(new_n743));
  INV_X1    g542(.A(new_n352), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n681), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n745), .A2(G15gat), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G15gat), .B1(new_n745), .B2(new_n725), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1326gat));
  XNOR2_X1  g548(.A(KEYINPUT43), .B(G22gat), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n752), .A3(new_n655), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n732), .B2(new_n655), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n755), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(new_n753), .A3(new_n750), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1327gat));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n350), .A2(new_n351), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n284), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n322), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n743), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n733), .A2(new_n299), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n764), .B1(new_n729), .B2(new_n731), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n769), .A2(KEYINPUT45), .A3(new_n299), .A4(new_n733), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n721), .A2(KEYINPUT110), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n669), .A2(new_n720), .A3(new_n772), .A4(new_n653), .ZN(new_n773));
  AND4_X1   g572(.A1(new_n719), .A2(new_n725), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n322), .B1(new_n683), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n323), .A2(new_n776), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n683), .B2(new_n727), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n777), .A2(new_n384), .A3(new_n763), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G29gat), .B1(new_n780), .B2(new_n678), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n768), .A2(new_n770), .A3(new_n781), .ZN(G1328gat));
  NAND2_X1  g581(.A1(new_n737), .A2(new_n300), .ZN(new_n783));
  OR3_X1    g582(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G36gat), .B1(new_n780), .B2(new_n736), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT46), .B1(new_n766), .B2(new_n783), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(G1329gat));
  INV_X1    g586(.A(G43gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n788), .A3(new_n681), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT47), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G43gat), .B1(new_n780), .B2(new_n725), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n792), .B(new_n789), .C1(new_n790), .C2(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1330gat));
  AOI21_X1  g595(.A(G50gat), .B1(new_n769), .B2(new_n655), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n655), .A2(G50gat), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n780), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT48), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT48), .B1(new_n797), .B2(new_n799), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1331gat));
  NAND2_X1  g603(.A1(new_n682), .A2(KEYINPUT35), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n604), .A2(new_n655), .A3(new_n385), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT92), .B1(new_n666), .B2(new_n670), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n719), .A2(new_n771), .A3(new_n725), .A4(new_n773), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR4_X1   g609(.A1(new_n761), .A2(new_n384), .A3(new_n322), .A4(new_n285), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n733), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g614(.A1(new_n812), .A2(new_n736), .ZN(new_n816));
  NOR2_X1   g615(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n817));
  AND2_X1   g616(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n816), .B2(new_n817), .ZN(G1333gat));
  INV_X1    g619(.A(G71gat), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n812), .B2(new_n746), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n725), .A2(new_n821), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n813), .A2(KEYINPUT112), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT112), .B1(new_n813), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g626(.A1(new_n813), .A2(new_n655), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g628(.A1(new_n762), .A2(new_n384), .A3(new_n285), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n323), .B1(new_n808), .B2(new_n809), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n779), .B(new_n830), .C1(new_n831), .C2(KEYINPUT44), .ZN(new_n832));
  OAI21_X1  g631(.A(G85gat), .B1(new_n832), .B2(new_n678), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n762), .A2(new_n384), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n322), .B(new_n834), .C1(new_n683), .C2(new_n774), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n810), .A2(KEYINPUT51), .A3(new_n322), .A4(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n284), .A2(new_n210), .A3(new_n733), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n833), .B1(new_n840), .B2(new_n841), .ZN(G1336gat));
  NOR3_X1   g641(.A1(new_n285), .A2(new_n736), .A3(G92gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n832), .A2(new_n736), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n209), .ZN(new_n846));
  XNOR2_X1  g645(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(G1337gat));
  INV_X1    g647(.A(G99gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n285), .A2(new_n746), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n839), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G99gat), .B1(new_n832), .B2(new_n725), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1338gat));
  NAND4_X1  g652(.A1(new_n777), .A2(new_n655), .A3(new_n779), .A4(new_n830), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n285), .A2(new_n670), .A3(G106gat), .ZN(new_n855));
  AOI22_X1  g654(.A1(G106gat), .A2(new_n854), .B1(new_n839), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT114), .B1(new_n854), .B2(G106gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT53), .ZN(new_n858));
  OAI21_X1  g657(.A(G106gat), .B1(new_n832), .B2(new_n670), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n855), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(KEYINPUT53), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n858), .A2(new_n863), .ZN(G1339gat));
  NOR2_X1   g663(.A1(new_n352), .A2(new_n384), .ZN(new_n865));
  INV_X1    g664(.A(new_n374), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n353), .A2(new_n356), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n368), .A2(new_n355), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n867), .A2(new_n354), .B1(new_n868), .B2(new_n367), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n363), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n322), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n251), .A2(new_n261), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n273), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n267), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n272), .B1(new_n281), .B2(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n871), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n268), .A2(new_n275), .A3(new_n276), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n876), .A2(KEYINPUT55), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT115), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n876), .A2(new_n877), .A3(new_n883), .A4(KEYINPUT55), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n880), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n870), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n277), .B2(new_n283), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n383), .B1(new_n878), .B2(new_n872), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n890), .B2(new_n322), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n865), .B1(new_n891), .B2(new_n761), .ZN(new_n892));
  NOR4_X1   g691(.A1(new_n892), .A2(new_n678), .A3(new_n655), .A4(new_n746), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(new_n736), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n384), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n284), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g697(.A1(new_n894), .A2(new_n762), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g699(.A1(new_n737), .A2(new_n323), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n413), .B1(new_n893), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n901), .B(KEYINPUT116), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n893), .A2(new_n413), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n904), .A2(new_n907), .A3(new_n908), .ZN(G1343gat));
  INV_X1    g708(.A(new_n272), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n266), .B1(new_n251), .B2(new_n261), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(KEYINPUT54), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n267), .B2(new_n875), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n883), .B1(new_n913), .B2(KEYINPUT55), .ZN(new_n914));
  INV_X1    g713(.A(new_n884), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n889), .B(new_n277), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n888), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n322), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n886), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n761), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n744), .A2(new_n383), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n725), .A2(new_n733), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n737), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n922), .A2(new_n655), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n387), .A3(new_n384), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT58), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT57), .B1(new_n892), .B2(new_n670), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT57), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n922), .A2(new_n930), .A3(new_n655), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n929), .A2(new_n931), .A3(new_n384), .A4(new_n924), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT118), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G141gat), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n932), .A2(KEYINPUT118), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n928), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n932), .A2(G141gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n926), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT58), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(G1344gat));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n389), .A3(new_n284), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n930), .B1(new_n922), .B2(new_n655), .ZN(new_n942));
  AOI211_X1 g741(.A(KEYINPUT57), .B(new_n670), .C1(new_n920), .C2(new_n921), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n284), .A3(new_n924), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT119), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT59), .B1(new_n946), .B2(new_n389), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n945), .A2(G148gat), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n945), .B2(G148gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n941), .B1(new_n948), .B2(new_n949), .ZN(G1345gat));
  NAND3_X1  g749(.A1(new_n925), .A2(new_n346), .A3(new_n762), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n944), .A2(new_n762), .A3(new_n924), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n346), .ZN(G1346gat));
  NAND3_X1  g752(.A1(new_n944), .A2(new_n322), .A3(new_n924), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n400), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n892), .A2(new_n670), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n923), .A2(new_n400), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n905), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n955), .A2(new_n958), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n736), .A2(new_n733), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n922), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n670), .A2(new_n681), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(G169gat), .A3(new_n384), .ZN(new_n965));
  INV_X1    g764(.A(G169gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n961), .A2(new_n963), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n383), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT120), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n965), .A2(KEYINPUT120), .A3(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1348gat));
  NAND3_X1  g772(.A1(new_n961), .A2(new_n670), .A3(new_n850), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g774(.A(new_n477), .B1(new_n967), .B2(new_n761), .ZN(new_n976));
  XNOR2_X1  g775(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n491), .A2(new_n494), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n961), .A2(new_n978), .A3(new_n963), .A4(new_n762), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n977), .B1(new_n976), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n980), .A2(new_n981), .ZN(G1350gat));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n322), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G190gat), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n983), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n964), .A2(new_n493), .A3(new_n322), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(G1351gat));
  INV_X1    g788(.A(G197gat), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n960), .A2(new_n725), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(KEYINPUT122), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n993), .A2(KEYINPUT123), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT123), .B1(new_n993), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g797(.A1(new_n998), .A2(new_n929), .A3(new_n384), .A4(new_n931), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n990), .B1(new_n999), .B2(KEYINPUT124), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n1000), .B1(KEYINPUT124), .B2(new_n999), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n892), .A2(new_n670), .A3(new_n991), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1002), .A2(new_n990), .A3(new_n384), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n1003), .ZN(G1352gat));
  AND2_X1   g803(.A1(new_n944), .A2(new_n998), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(new_n284), .ZN(new_n1006));
  XNOR2_X1  g805(.A(KEYINPUT125), .B(G204gat), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n285), .A2(new_n1007), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g809(.A(new_n1010), .B(KEYINPUT62), .Z(new_n1011));
  NAND2_X1  g810(.A1(new_n1008), .A2(new_n1011), .ZN(G1353gat));
  AOI21_X1  g811(.A(new_n761), .B1(new_n993), .B2(new_n995), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n929), .A2(new_n931), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT63), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1014), .A2(new_n1015), .A3(G211gat), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n761), .A2(G211gat), .ZN(new_n1017));
  NAND4_X1  g816(.A1(new_n956), .A2(KEYINPUT126), .A3(new_n992), .A4(new_n1017), .ZN(new_n1018));
  NAND4_X1  g817(.A1(new_n922), .A2(new_n655), .A3(new_n992), .A4(new_n1017), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g822(.A(new_n1015), .B1(new_n1014), .B2(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(KEYINPUT127), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1014), .A2(G211gat), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1026), .A2(KEYINPUT63), .ZN(new_n1027));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1028));
  NAND4_X1  g827(.A1(new_n1027), .A2(new_n1028), .A3(new_n1016), .A4(new_n1022), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1025), .A2(new_n1029), .ZN(G1354gat));
  AOI21_X1  g829(.A(G218gat), .B1(new_n1002), .B2(new_n322), .ZN(new_n1031));
  AND2_X1   g830(.A1(new_n322), .A2(G218gat), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1031), .B1(new_n1005), .B2(new_n1032), .ZN(G1355gat));
endmodule


