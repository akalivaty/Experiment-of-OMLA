//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G116), .A2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n214), .B(new_n220), .C1(G97), .C2(G257), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G1), .B2(G20), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n209), .B(new_n223), .C1(new_n225), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  OR2_X1    g0043(.A1(KEYINPUT8), .A2(G58), .ZN(new_n244));
  NAND2_X1  g0044(.A1(KEYINPUT8), .A2(G58), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n206), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G150), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  OAI22_X1  g0050(.A1(new_n246), .A2(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT65), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(new_n206), .B2(new_n201), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n224), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G50), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n255), .B1(new_n205), .B2(G20), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n260), .A2(G50), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n256), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT9), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G223), .A2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G222), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n267), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n274), .B(new_n277), .C1(G77), .C2(new_n270), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n276), .A2(new_n279), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n278), .B(new_n282), .C1(new_n217), .C2(new_n283), .ZN(new_n284));
  XOR2_X1   g0084(.A(new_n284), .B(KEYINPUT64), .Z(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G200), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n256), .A2(KEYINPUT9), .A3(new_n259), .A4(new_n262), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n284), .B(KEYINPUT64), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G190), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n265), .A2(new_n286), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT10), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n289), .A2(new_n287), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT10), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n292), .A2(new_n293), .A3(new_n286), .A4(new_n265), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT15), .B(G87), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n246), .A2(new_n250), .B1(new_n296), .B2(new_n247), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n206), .A2(new_n202), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n255), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n257), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n202), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n260), .A2(G77), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n303), .A2(new_n304), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n272), .A2(G232), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n270), .B(new_n309), .C1(new_n219), .C2(new_n272), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n277), .C1(G107), .C2(new_n270), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n311), .B(new_n282), .C1(new_n211), .C2(new_n283), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G200), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n308), .B(new_n313), .C1(new_n314), .C2(new_n312), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n317), .B1(G179), .B2(new_n312), .C1(new_n306), .C2(new_n307), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  INV_X1    g0120(.A(new_n263), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT66), .B1(new_n285), .B2(G179), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT66), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n288), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n285), .A2(new_n316), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n295), .A2(new_n320), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT69), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n291), .A2(new_n294), .B1(new_n327), .B2(new_n326), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n333), .A2(KEYINPUT69), .A3(new_n320), .A4(new_n329), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n276), .A2(G232), .A3(new_n279), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT76), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n217), .A2(G1698), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n338), .B1(G223), .B2(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n267), .B2(new_n212), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n277), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n282), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G169), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n337), .A2(new_n343), .A3(G179), .A4(new_n282), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n339), .A2(new_n340), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT7), .B1(new_n350), .B2(new_n206), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n269), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n349), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n268), .A2(new_n206), .A3(new_n269), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n349), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n218), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G58), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n218), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G58), .A2(G68), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n249), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n348), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n351), .B2(new_n353), .ZN(new_n367));
  INV_X1    g0167(.A(new_n365), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n369), .A2(new_n255), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n205), .A2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n244), .A2(new_n372), .A3(new_n245), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n300), .A2(new_n255), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n244), .A2(new_n372), .A3(KEYINPUT73), .A4(new_n245), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n246), .A2(new_n300), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n378), .A2(KEYINPUT74), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT74), .B1(new_n378), .B2(new_n379), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT75), .B1(new_n371), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n355), .A2(new_n356), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT72), .B1(new_n384), .B2(new_n352), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n385), .B2(new_n357), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT16), .B1(new_n386), .B2(new_n368), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n369), .A2(new_n255), .ZN(new_n388));
  OAI211_X1 g0188(.A(KEYINPUT75), .B(new_n382), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n347), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT77), .A3(KEYINPUT18), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n344), .A2(new_n314), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n344), .A2(G200), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n371), .A2(new_n393), .A3(new_n382), .A4(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT17), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n382), .B1(new_n387), .B2(new_n388), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n389), .ZN(new_n400));
  OR2_X1    g0200(.A1(KEYINPUT77), .A2(KEYINPUT18), .ZN(new_n401));
  NAND2_X1  g0201(.A1(KEYINPUT77), .A2(KEYINPUT18), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n400), .A2(new_n347), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n392), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n218), .A2(G20), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n405), .B1(new_n247), .B2(new_n202), .C1(new_n250), .C2(new_n216), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n255), .ZN(new_n407));
  XOR2_X1   g0207(.A(KEYINPUT71), .B(KEYINPUT11), .Z(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G13), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n405), .A2(G1), .A3(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n260), .A2(G68), .B1(KEYINPUT12), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n407), .A2(new_n409), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n415), .B(new_n416), .C1(KEYINPUT12), .C2(new_n412), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n217), .A2(new_n272), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n270), .B(new_n418), .C1(G232), .C2(new_n272), .ZN(new_n419));
  INV_X1    g0219(.A(G97), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n267), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n276), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n283), .A2(new_n219), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n423), .A2(new_n281), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR4_X1   g0228(.A1(new_n423), .A2(new_n281), .A3(new_n426), .A4(new_n424), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n417), .B1(new_n430), .B2(G200), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(new_n429), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G190), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n404), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(G169), .B1(new_n428), .B2(new_n429), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT14), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(G179), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(G169), .C1(new_n428), .C2(new_n429), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n417), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n335), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT80), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n275), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n205), .B(G45), .C1(new_n275), .C2(KEYINPUT5), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n277), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT81), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n449), .A2(new_n456), .A3(new_n450), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n457), .A2(G274), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n453), .B1(new_n451), .B2(KEYINPUT81), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n455), .A2(G270), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G264), .A2(G1698), .ZN(new_n461));
  INV_X1    g0261(.A(G257), .ZN(new_n462));
  OAI221_X1 g0262(.A(new_n461), .B1(new_n462), .B2(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(new_n277), .C1(G303), .C2(new_n270), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G200), .ZN(new_n466));
  INV_X1    g0266(.A(G116), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n300), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n376), .B1(G1), .B2(new_n267), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(new_n206), .C1(G33), .C2(new_n420), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(new_n255), .C1(new_n206), .C2(G116), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT20), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n472), .A2(new_n473), .ZN(new_n475));
  OAI221_X1 g0275(.A(new_n468), .B1(new_n469), .B2(new_n467), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n466), .A2(new_n477), .A3(KEYINPUT86), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT86), .B1(new_n466), .B2(new_n477), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n465), .A2(new_n314), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n296), .A2(new_n300), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n270), .A2(new_n206), .A3(G68), .ZN(new_n483));
  XOR2_X1   g0283(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n484));
  NOR2_X1   g0284(.A1(new_n247), .A2(new_n420), .ZN(new_n485));
  AOI21_X1  g0285(.A(G20), .B1(new_n484), .B2(new_n421), .ZN(new_n486));
  NOR3_X1   g0286(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n487));
  OAI221_X1 g0287(.A(new_n483), .B1(new_n484), .B2(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n482), .B1(new_n488), .B2(new_n255), .ZN(new_n489));
  INV_X1    g0289(.A(new_n469), .ZN(new_n490));
  XOR2_X1   g0290(.A(new_n296), .B(KEYINPUT85), .Z(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n211), .B1(new_n268), .B2(new_n269), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G1698), .ZN(new_n494));
  OAI211_X1 g0294(.A(G238), .B(new_n272), .C1(new_n339), .C2(new_n340), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT83), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n270), .A2(KEYINPUT83), .A3(G238), .A4(new_n272), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G116), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n494), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n277), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n205), .A2(G45), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n213), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n276), .B(new_n503), .C1(G274), .C2(new_n502), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n489), .A2(new_n492), .B1(new_n505), .B2(new_n316), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G179), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n469), .A2(new_n212), .ZN(new_n508));
  AOI211_X1 g0308(.A(new_n482), .B(new_n508), .C1(new_n488), .C2(new_n255), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(G200), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n509), .B(new_n510), .C1(new_n314), .C2(new_n505), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(G274), .A3(new_n454), .A4(new_n457), .ZN(new_n514));
  OAI211_X1 g0314(.A(G270), .B(new_n276), .C1(new_n451), .C2(new_n453), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n514), .A2(new_n464), .A3(G179), .A4(new_n515), .ZN(new_n516));
  OR2_X1    g0316(.A1(new_n477), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n476), .A2(new_n465), .A3(G169), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n476), .A2(new_n465), .A3(KEYINPUT21), .A4(G169), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n481), .A2(new_n512), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT82), .ZN(new_n524));
  INV_X1    g0324(.A(G200), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n270), .A2(G250), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n272), .B1(new_n526), .B2(KEYINPUT4), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G1698), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n529), .B(G244), .C1(new_n340), .C2(new_n339), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(new_n470), .C1(new_n493), .C2(KEYINPUT4), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n277), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT79), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(KEYINPUT79), .B(new_n277), .C1(new_n527), .C2(new_n531), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(G257), .B(new_n276), .C1(new_n451), .C2(new_n453), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n514), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n525), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G107), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n354), .B2(new_n358), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT78), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n250), .A2(new_n202), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT6), .ZN(new_n547));
  XNOR2_X1  g0347(.A(G97), .B(G107), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n542), .B(new_n544), .C1(new_n549), .C2(new_n206), .ZN(new_n550));
  AND2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n206), .B1(new_n553), .B2(new_n545), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT78), .B1(new_n554), .B2(new_n543), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n255), .B1(new_n541), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n300), .A2(new_n420), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n490), .A2(G97), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n538), .A2(new_n532), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n561), .A2(new_n314), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n539), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n536), .A2(new_n324), .A3(new_n538), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n316), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n564), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n524), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n536), .A2(new_n538), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n557), .A2(new_n558), .ZN(new_n570));
  INV_X1    g0370(.A(new_n562), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n559), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n564), .A2(new_n560), .A3(new_n565), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(KEYINPUT82), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n462), .A2(G1698), .ZN(new_n576));
  OAI221_X1 g0376(.A(new_n576), .B1(G250), .B2(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n577));
  INV_X1    g0377(.A(G294), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n267), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n455), .A2(G264), .B1(new_n579), .B2(new_n277), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(G190), .A3(new_n514), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT25), .ZN(new_n582));
  AOI211_X1 g0382(.A(G107), .B(new_n257), .C1(KEYINPUT87), .C2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(KEYINPUT87), .B2(new_n582), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT87), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(KEYINPUT25), .C1(new_n257), .C2(G107), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n584), .B(new_n586), .C1(new_n540), .C2(new_n469), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT88), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n580), .A2(new_n514), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G200), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n270), .A2(new_n206), .A3(G87), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n591), .B(KEYINPUT22), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n206), .A2(G107), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n594), .B(KEYINPUT23), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT24), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n592), .A2(KEYINPUT24), .A3(new_n593), .A4(new_n595), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n255), .A3(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n588), .A2(new_n590), .A3(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n588), .A2(new_n600), .B1(new_n316), .B2(new_n589), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n580), .A2(new_n324), .A3(new_n514), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n581), .A2(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n446), .A2(new_n523), .A3(new_n575), .A4(new_n604), .ZN(G372));
  NAND2_X1  g0405(.A1(new_n397), .A2(new_n347), .ZN(new_n606));
  XOR2_X1   g0406(.A(new_n606), .B(KEYINPUT18), .Z(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n445), .B1(new_n437), .B2(new_n318), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(new_n396), .ZN(new_n610));
  INV_X1    g0410(.A(new_n295), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n328), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n446), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n566), .A2(new_n511), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT26), .ZN(new_n616));
  INV_X1    g0416(.A(new_n522), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n588), .A2(new_n600), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n589), .A2(new_n316), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(new_n603), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n617), .A2(new_n620), .B1(new_n581), .B2(new_n601), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n566), .B1(new_n621), .B2(new_n572), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n511), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n507), .B(new_n616), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n613), .B1(new_n614), .B2(new_n626), .ZN(G369));
  NOR2_X1   g0427(.A1(new_n411), .A2(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n205), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G213), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n617), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n601), .A2(new_n581), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n618), .A2(new_n634), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n620), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n602), .A2(new_n603), .A3(new_n634), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(KEYINPUT89), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(KEYINPUT89), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n635), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n634), .B(KEYINPUT90), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n602), .A2(new_n603), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n641), .A2(new_n642), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n481), .A2(new_n522), .ZN(new_n648));
  INV_X1    g0448(.A(new_n634), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n477), .A2(new_n649), .ZN(new_n650));
  MUX2_X1   g0450(.A(new_n648), .B(new_n522), .S(new_n650), .Z(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT91), .Z(G399));
  INV_X1    g0455(.A(new_n207), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G41), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n487), .A2(new_n467), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n657), .A2(new_n658), .A3(new_n205), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n227), .B2(new_n657), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n660), .B(KEYINPUT28), .Z(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT29), .B1(new_n625), .B2(new_n644), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n617), .A2(new_n620), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n572), .A3(new_n636), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n624), .B1(new_n664), .B2(new_n573), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n616), .A2(new_n507), .ZN(new_n666));
  OAI211_X1 g0466(.A(KEYINPUT29), .B(new_n649), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n505), .A2(new_n465), .A3(new_n324), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n568), .A3(new_n589), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n460), .A2(KEYINPUT92), .A3(G179), .A4(new_n464), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT92), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n516), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n561), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n580), .A2(new_n504), .A3(new_n501), .ZN(new_n679));
  AND4_X1   g0479(.A1(new_n673), .A2(new_n677), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n561), .B1(new_n674), .B2(new_n676), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n673), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n672), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT93), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(KEYINPUT93), .B(new_n672), .C1(new_n680), .C2(new_n682), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n634), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT31), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n575), .A2(new_n523), .A3(new_n604), .A4(new_n644), .ZN(new_n690));
  INV_X1    g0490(.A(new_n644), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n670), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n661), .B1(new_n696), .B2(G1), .ZN(G364));
  XOR2_X1   g0497(.A(new_n652), .B(KEYINPUT94), .Z(new_n698));
  INV_X1    g0498(.A(new_n657), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n628), .A2(G45), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G1), .A3(new_n700), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n698), .B(new_n701), .C1(G330), .C2(new_n651), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT95), .Z(new_n703));
  NOR2_X1   g0503(.A1(G13), .A2(G33), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n224), .B1(G20), .B2(new_n316), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n350), .A2(new_n207), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT96), .Z(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G45), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n227), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n239), .A2(G45), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n714), .A2(new_n715), .B1(new_n467), .B2(new_n656), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n270), .A2(new_n207), .A3(G355), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n709), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n206), .A2(new_n324), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n720), .A2(G190), .A3(G200), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G311), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n720), .A2(new_n314), .A3(G200), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n270), .B1(new_n725), .B2(G322), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n720), .A2(new_n525), .A3(G190), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT33), .B(G317), .Z(new_n729));
  OAI21_X1  g0529(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G179), .A2(G200), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n206), .B1(new_n731), .B2(G190), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n724), .B(new_n730), .C1(G294), .C2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n314), .A2(new_n525), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n719), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G326), .ZN(new_n738));
  NOR4_X1   g0538(.A1(new_n206), .A2(new_n525), .A3(G179), .A4(G190), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT97), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT97), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G283), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n735), .A2(G20), .A3(new_n324), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n731), .A2(G20), .A3(new_n314), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n746), .A2(G303), .B1(G329), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n734), .A2(new_n738), .A3(new_n744), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n743), .A2(G107), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n751), .B(new_n270), .C1(new_n212), .C2(new_n745), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT98), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n218), .A2(new_n728), .B1(new_n722), .B2(new_n202), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n737), .A2(G50), .B1(new_n733), .B2(G97), .ZN(new_n755));
  INV_X1    g0555(.A(new_n725), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(new_n360), .ZN(new_n757));
  OR3_X1    g0557(.A1(new_n753), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n748), .A2(G159), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT32), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n750), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n718), .B1(new_n761), .B2(new_n707), .ZN(new_n762));
  INV_X1    g0562(.A(new_n706), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n651), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n703), .B1(new_n701), .B2(new_n764), .ZN(G396));
  OAI21_X1  g0565(.A(new_n315), .B1(new_n308), .B2(new_n649), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n318), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n318), .A2(new_n634), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n626), .B2(new_n691), .ZN(new_n770));
  INV_X1    g0570(.A(new_n769), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n644), .B(new_n771), .C1(new_n665), .C2(new_n666), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(new_n694), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n694), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n701), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n743), .A2(G87), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n723), .B2(new_n747), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT100), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n728), .A2(new_n780), .B1(new_n732), .B2(new_n420), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n350), .B1(new_n782), .B2(new_n736), .C1(new_n756), .C2(new_n578), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n781), .B(new_n783), .C1(G107), .C2(new_n746), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n779), .B(new_n784), .C1(new_n467), .C2(new_n722), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G143), .A2(new_n725), .B1(new_n727), .B2(G150), .ZN(new_n786));
  INV_X1    g0586(.A(G137), .ZN(new_n787));
  INV_X1    g0587(.A(G159), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(new_n787), .B2(new_n736), .C1(new_n788), .C2(new_n722), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT34), .ZN(new_n790));
  INV_X1    g0590(.A(G132), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n270), .B1(new_n747), .B2(new_n791), .C1(new_n360), .C2(new_n732), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n743), .B2(G68), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n790), .B(new_n793), .C1(new_n216), .C2(new_n745), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n785), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n707), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n707), .A2(new_n704), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT99), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n796), .B1(G77), .B2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n701), .B(new_n800), .C1(new_n704), .C2(new_n769), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT101), .Z(new_n802));
  NAND2_X1  g0602(.A1(new_n776), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT102), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G384));
  XOR2_X1   g0605(.A(new_n549), .B(KEYINPUT103), .Z(new_n806));
  AOI21_X1  g0606(.A(new_n467), .B1(new_n806), .B2(KEYINPUT35), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n807), .B(new_n225), .C1(KEYINPUT35), .C2(new_n806), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT104), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT36), .ZN(new_n810));
  OAI21_X1  g0610(.A(G77), .B1(new_n360), .B2(new_n218), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n811), .A2(new_n226), .B1(G50), .B2(new_n218), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(G1), .A3(new_n411), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n384), .A2(new_n352), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n365), .B1(new_n814), .B2(G68), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(KEYINPUT16), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n388), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n632), .B1(new_n818), .B2(new_n382), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n404), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n632), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n383), .A2(new_n390), .B1(new_n347), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT37), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n395), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n382), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n347), .A2(new_n821), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n395), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n822), .A2(new_n824), .B1(KEYINPUT37), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT38), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT38), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n831), .B(new_n828), .C1(new_n404), .C2(new_n819), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT39), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT106), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n820), .A2(KEYINPUT38), .A3(new_n829), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n400), .A2(new_n821), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n837), .A2(new_n395), .A3(new_n606), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(KEYINPUT37), .B1(new_n824), .B2(new_n822), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n837), .B1(new_n607), .B2(new_n396), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n831), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT39), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n836), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n833), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n835), .B1(new_n844), .B2(new_n834), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n445), .A2(KEYINPUT105), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT105), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n444), .B2(new_n417), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n846), .A2(new_n634), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n608), .A2(new_n632), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n417), .A2(new_n634), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n436), .B(new_n852), .C1(new_n846), .C2(new_n848), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n444), .A2(new_n417), .A3(new_n634), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n772), .B2(new_n768), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n820), .A2(new_n829), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n831), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n836), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n850), .A2(new_n851), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n669), .A2(new_n446), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n613), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n861), .B(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(KEYINPUT107), .A2(KEYINPUT31), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n687), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n865), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n685), .A2(new_n634), .A3(new_n686), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n690), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT108), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n866), .A2(new_n690), .A3(KEYINPUT108), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n853), .A2(new_n854), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n771), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n859), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n875), .B1(new_n871), .B2(new_n872), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n836), .A2(new_n841), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n878), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n877), .A2(new_n878), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n446), .A2(new_n873), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n882), .B(new_n883), .Z(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(G330), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n864), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n886), .A2(KEYINPUT109), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(KEYINPUT109), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n887), .B(new_n888), .C1(new_n864), .C2(new_n885), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n628), .A2(new_n205), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n810), .B(new_n813), .C1(new_n889), .C2(new_n890), .ZN(G367));
  INV_X1    g0691(.A(new_n653), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n573), .A2(new_n644), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT110), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n691), .A2(new_n560), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n572), .A2(new_n573), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n509), .A2(new_n649), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n507), .A2(new_n902), .A3(new_n511), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n507), .B2(new_n902), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n905));
  OR3_X1    g0705(.A1(new_n643), .A2(KEYINPUT42), .A3(new_n898), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n573), .B1(new_n898), .B2(new_n620), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n644), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT42), .B1(new_n643), .B2(new_n898), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n900), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n900), .B1(new_n910), .B2(new_n905), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OR3_X1    g0715(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n915), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n657), .B(KEYINPUT41), .Z(new_n918));
  NAND3_X1  g0718(.A1(new_n643), .A2(new_n645), .A3(new_n897), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT45), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n646), .A2(new_n898), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT111), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT44), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(KEYINPUT44), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n923), .A2(KEYINPUT44), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n646), .A2(new_n898), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n921), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(KEYINPUT112), .A3(new_n653), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n647), .B1(new_n617), .B2(new_n634), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n643), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n698), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n892), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(new_n695), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n653), .A2(KEYINPUT112), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n921), .A2(new_n935), .A3(new_n924), .A4(new_n927), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n918), .B1(new_n937), .B2(new_n696), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n700), .A2(G1), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n916), .B(new_n917), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n746), .A2(G58), .B1(G137), .B2(new_n748), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n737), .A2(G143), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n941), .B(new_n942), .C1(new_n248), .C2(new_n756), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G68), .B2(new_n733), .ZN(new_n944));
  AOI22_X1  g0744(.A1(G50), .A2(new_n721), .B1(new_n727), .B2(G159), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT113), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n743), .A2(G77), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n944), .A2(new_n946), .A3(new_n270), .A4(new_n947), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n350), .B1(new_n723), .B2(new_n736), .C1(new_n756), .C2(new_n782), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n742), .A2(new_n420), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n745), .A2(new_n467), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT46), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n721), .A2(G283), .B1(G107), .B2(new_n733), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n953), .B(new_n954), .C1(new_n578), .C2(new_n728), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n748), .A2(G317), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n948), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT47), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n701), .B1(new_n958), .B2(new_n707), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n708), .B1(new_n207), .B2(new_n296), .C1(new_n712), .C2(new_n235), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n763), .C2(new_n904), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n940), .A2(new_n961), .ZN(G387));
  INV_X1    g0762(.A(KEYINPUT116), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n934), .B2(new_n699), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n933), .A2(new_n695), .ZN(new_n965));
  OAI211_X1 g0765(.A(KEYINPUT116), .B(new_n657), .C1(new_n933), .C2(new_n695), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n932), .A2(new_n892), .A3(new_n939), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n711), .B1(new_n232), .B2(new_n713), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n658), .A2(new_n207), .A3(new_n270), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n218), .A2(new_n202), .ZN(new_n972));
  INV_X1    g0772(.A(new_n246), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n216), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n658), .B1(new_n974), .B2(KEYINPUT50), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n975), .B(new_n713), .C1(KEYINPUT50), .C2(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n971), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n656), .A2(new_n540), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n709), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n721), .A2(G303), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n727), .A2(G311), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n725), .A2(G317), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n737), .A2(G322), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n986));
  AOI22_X1  g0786(.A1(new_n985), .A2(new_n986), .B1(G283), .B2(new_n733), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n578), .B2(new_n745), .C1(new_n986), .C2(new_n985), .ZN(new_n988));
  XNOR2_X1  g0788(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n748), .A2(G326), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n270), .B1(new_n743), .B2(G116), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n728), .A2(new_n246), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n270), .B1(new_n722), .B2(new_n218), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(G50), .C2(new_n725), .ZN(new_n997));
  INV_X1    g0797(.A(new_n950), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n491), .A2(new_n733), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n736), .A2(new_n788), .B1(new_n248), .B2(new_n747), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G77), .B2(new_n746), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n994), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n979), .B1(new_n1003), .B2(new_n707), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n647), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n1005), .B2(new_n763), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n967), .B(new_n968), .C1(new_n701), .C2(new_n1006), .ZN(G393));
  NAND2_X1  g0807(.A1(new_n928), .A2(new_n653), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n921), .A2(new_n892), .A3(new_n924), .A4(new_n927), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n939), .A3(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n725), .A2(G311), .B1(new_n737), .B2(G317), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT52), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n727), .A2(G303), .B1(G116), .B2(new_n733), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n270), .B1(new_n748), .B2(G322), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n746), .A2(G283), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n751), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1012), .B(new_n1016), .C1(G294), .C2(new_n721), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n350), .B1(new_n748), .B2(G143), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n777), .B(new_n1018), .C1(new_n218), .C2(new_n745), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n727), .A2(G50), .B1(G77), .B2(new_n733), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n246), .B2(new_n722), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n725), .A2(G159), .B1(new_n737), .B2(G150), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT51), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT117), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n701), .B1(new_n1026), .B2(new_n707), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n708), .B1(new_n420), .B2(new_n207), .C1(new_n712), .C2(new_n242), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n763), .C2(new_n897), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1010), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n934), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n929), .A2(new_n936), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n934), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1030), .B1(new_n1033), .B2(new_n657), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(G390));
  OAI211_X1 g0835(.A(new_n649), .B(new_n767), .C1(new_n665), .C2(new_n666), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n855), .B1(new_n1036), .B2(new_n768), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1037), .A2(new_n849), .A3(new_n880), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n834), .B1(new_n833), .B2(new_n843), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT106), .B1(new_n859), .B2(KEYINPUT39), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n856), .A2(new_n849), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1038), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n771), .A2(G330), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1045), .B(new_n855), .C1(new_n871), .C2(new_n872), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(KEYINPUT118), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1045), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n693), .A3(new_n874), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT118), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1042), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n1046), .C1(new_n1053), .C2(new_n1038), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1048), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n446), .A2(G330), .A3(new_n873), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1056), .A2(new_n862), .A3(new_n613), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n873), .A2(new_n1049), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(KEYINPUT119), .A3(new_n855), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1050), .A2(KEYINPUT119), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1045), .B1(new_n871), .B2(new_n872), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n874), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1036), .A2(new_n768), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1059), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n772), .A2(new_n768), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n874), .B1(new_n1049), .B2(new_n693), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1046), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1057), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1055), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1048), .A2(new_n1051), .A3(new_n1054), .A4(new_n1068), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n657), .A3(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1048), .A2(new_n1051), .A3(new_n939), .A4(new_n1054), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(KEYINPUT54), .B(G143), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n787), .A2(new_n728), .B1(new_n722), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G159), .B2(new_n733), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n745), .A2(new_n248), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT53), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n743), .A2(G50), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n270), .B1(new_n756), .B2(new_n791), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G128), .B2(new_n737), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G125), .B2(new_n748), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT120), .Z(new_n1084));
  OAI221_X1 g0884(.A(new_n350), .B1(new_n212), .B2(new_n745), .C1(new_n756), .C2(new_n467), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G283), .B2(new_n737), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n742), .A2(new_n218), .B1(new_n578), .B2(new_n747), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT121), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n727), .A2(G107), .B1(G77), .B2(new_n733), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(KEYINPUT121), .B2(new_n1087), .C1(new_n420), .C2(new_n722), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n701), .B1(new_n1092), .B2(new_n707), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n973), .B2(new_n799), .C1(new_n845), .C2(new_n705), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1073), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1072), .A2(new_n1095), .ZN(G378));
  INV_X1    g0896(.A(new_n1057), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1071), .A2(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n850), .A2(new_n851), .A3(new_n860), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n333), .B(KEYINPUT55), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n263), .A2(new_n821), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT56), .Z(new_n1102));
  OR2_X1    g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT124), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1103), .A2(KEYINPUT124), .A3(new_n1104), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n882), .C2(G330), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n882), .A2(G330), .A3(new_n1106), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1099), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n882), .A2(G330), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1106), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n861), .B(new_n1108), .C1(new_n1113), .C2(new_n1105), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1098), .A2(new_n1115), .A3(KEYINPUT57), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n657), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT57), .B1(new_n1098), .B2(new_n1115), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1103), .A2(new_n704), .A3(new_n1104), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n270), .B1(new_n746), .B2(G77), .ZN(new_n1121));
  AOI21_X1  g0921(.A(G41), .B1(new_n733), .B2(G68), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n728), .C2(new_n420), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n743), .A2(G58), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n491), .A2(new_n721), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n725), .A2(G107), .B1(new_n737), .B2(G116), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1123), .B(new_n1127), .C1(G283), .C2(new_n748), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT58), .Z(new_n1129));
  OAI21_X1  g0929(.A(new_n216), .B1(new_n339), .B2(G41), .ZN(new_n1130));
  AOI21_X1  g0930(.A(G33), .B1(new_n748), .B2(G124), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n275), .B(new_n1131), .C1(new_n742), .C2(new_n788), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT123), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(G125), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n745), .A2(new_n1074), .B1(new_n736), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G128), .B2(new_n725), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G132), .A2(new_n727), .B1(new_n721), .B2(G137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(new_n248), .C2(new_n732), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT122), .Z(new_n1140));
  OR2_X1    g0940(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1129), .B(new_n1130), .C1(new_n1134), .C2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n701), .B1(new_n1145), .B2(new_n707), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1120), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n216), .B2(new_n797), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1115), .B2(new_n939), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1119), .A2(new_n1149), .ZN(G375));
  OAI221_X1 g0950(.A(new_n350), .B1(new_n722), .B2(new_n540), .C1(new_n467), .C2(new_n728), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G294), .B2(new_n737), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n756), .A2(new_n780), .B1(new_n782), .B2(new_n747), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G97), .B2(new_n746), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1152), .A2(new_n947), .A3(new_n999), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n270), .B1(new_n722), .B2(new_n248), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n728), .A2(new_n1074), .B1(new_n732), .B2(new_n216), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(G137), .C2(new_n725), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n737), .A2(G132), .B1(G128), .B2(new_n748), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1124), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n745), .A2(new_n788), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1155), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n707), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(G68), .B2(new_n799), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n701), .B(new_n1164), .C1(new_n855), .C2(new_n704), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n939), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1064), .A2(new_n1067), .A3(new_n1057), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(new_n918), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1167), .B1(new_n1170), .B2(new_n1068), .ZN(G381));
  INV_X1    g0971(.A(KEYINPUT125), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1072), .A2(new_n1172), .A3(new_n1095), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n1072), .B2(new_n1095), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n1149), .A3(new_n1119), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1176), .A2(G384), .A3(G381), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1034), .A2(new_n940), .A3(new_n961), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1178), .A2(G396), .A3(G393), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(G407));
  OAI211_X1 g0980(.A(G407), .B(G213), .C1(G343), .C2(new_n1176), .ZN(G409));
  NAND2_X1  g0981(.A1(new_n1098), .A2(new_n1115), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1149), .B1(new_n1182), .B2(new_n918), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G378), .B(new_n1149), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT60), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1168), .B1(new_n1068), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT126), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1169), .A2(KEYINPUT60), .ZN(new_n1191));
  OAI211_X1 g0991(.A(KEYINPUT126), .B(new_n1168), .C1(new_n1068), .C2(new_n1187), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1190), .A2(new_n657), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1193), .A2(G384), .A3(new_n1167), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G384), .B1(new_n1193), .B2(new_n1167), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(G213), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(G343), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1186), .A2(KEYINPUT63), .A3(new_n1196), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(G387), .A2(G390), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(G393), .B(G396), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1201), .A2(new_n1178), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(new_n1201), .B2(new_n1178), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1200), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1198), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1198), .A2(G2897), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1193), .A2(new_n1167), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n804), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1193), .A2(G384), .A3(new_n1167), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1208), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT63), .B1(new_n1207), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1207), .A2(new_n1196), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT61), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1206), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT62), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1186), .A2(new_n1221), .A3(new_n1196), .A4(new_n1199), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1219), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1207), .B2(new_n1215), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1217), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1220), .B1(new_n1225), .B2(new_n1205), .ZN(G405));
  NAND2_X1  g1026(.A1(G375), .A2(new_n1175), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1185), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1196), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1227), .B(new_n1185), .C1(new_n1195), .C2(new_n1194), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1205), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1229), .A2(new_n1205), .A3(new_n1230), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(G402));
endmodule


