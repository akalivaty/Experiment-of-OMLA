//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1112,
    new_n1113, new_n1114;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n461), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n463), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n470), .B(new_n472), .C1(new_n461), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n462), .B1(new_n463), .B2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n473), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(G2105), .A3(new_n464), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI221_X1 g061(.A(new_n481), .B1(new_n468), .B2(new_n482), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI21_X1  g063(.A(G2104), .B1(new_n461), .B2(G114), .ZN(new_n489));
  INV_X1    g064(.A(G102), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(new_n461), .ZN(new_n491));
  INV_X1    g066(.A(new_n485), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G126), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n468), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n461), .A3(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n475), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n511), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  XNOR2_X1  g094(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n513), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n522), .B1(G89), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT68), .B(G51), .Z(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n515), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT69), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n526), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n510), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n513), .A2(new_n534), .B1(new_n515), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n507), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(KEYINPUT72), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(KEYINPUT72), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(G651), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n515), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n523), .A2(G81), .B1(G43), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT73), .Z(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  NOR3_X1   g130(.A1(new_n515), .A2(KEYINPUT74), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT76), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n557), .B1(G651), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n523), .A2(G91), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT75), .Z(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n544), .A2(G49), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT77), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n523), .A2(G87), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(new_n544), .A2(G48), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n507), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n571), .B(new_n575), .C1(new_n576), .C2(new_n513), .ZN(G305));
  AOI22_X1  g152(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n510), .ZN(new_n579));
  INV_X1    g154(.A(G85), .ZN(new_n580));
  INV_X1    g155(.A(G47), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n513), .A2(new_n580), .B1(new_n515), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n523), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n587));
  XOR2_X1   g162(.A(new_n586), .B(new_n587), .Z(new_n588));
  AOI22_X1  g163(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G54), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n589), .A2(new_n510), .B1(new_n590), .B2(new_n515), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n585), .B1(new_n592), .B2(G868), .ZN(G321));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G299), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(new_n595), .B2(G168), .ZN(G297));
  OAI21_X1  g172(.A(new_n596), .B1(new_n595), .B2(G168), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n546), .A2(new_n595), .ZN(new_n601));
  INV_X1    g176(.A(new_n592), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n603), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(KEYINPUT80), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(KEYINPUT80), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n607), .B(new_n608), .C1(G111), .C2(new_n461), .ZN(new_n609));
  INV_X1    g184(.A(G135), .ZN(new_n610));
  INV_X1    g185(.A(G123), .ZN(new_n611));
  OAI221_X1 g186(.A(new_n609), .B1(new_n468), .B2(new_n610), .C1(new_n485), .C2(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(KEYINPUT81), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(KEYINPUT81), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G2096), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n476), .A2(new_n471), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT79), .B(KEYINPUT13), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n619), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n617), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2438), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2430), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n637), .A2(G14), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2072), .B(G2078), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(KEYINPUT17), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n645), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT85), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n643), .A3(new_n639), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT18), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n647), .A2(new_n639), .A3(new_n641), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n616), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n657), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n658), .A2(new_n659), .ZN(new_n663));
  AOI22_X1  g238(.A1(new_n661), .A2(KEYINPUT20), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n657), .A3(new_n660), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n664), .B(new_n666), .C1(KEYINPUT20), .C2(new_n661), .ZN(new_n667));
  XOR2_X1   g242(.A(G1991), .B(G1996), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  NAND2_X1  g248(.A1(new_n469), .A2(G131), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT86), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n492), .A2(G119), .ZN(new_n676));
  NOR2_X1   g251(.A1(G95), .A2(G2105), .ZN(new_n677));
  OAI21_X1  g252(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n676), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT87), .Z(new_n680));
  MUX2_X1   g255(.A(G25), .B(new_n680), .S(G29), .Z(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT35), .B(G1991), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G24), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n583), .B2(new_n684), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(G1986), .Z(new_n687));
  OAI21_X1  g262(.A(KEYINPUT88), .B1(G16), .B2(G23), .ZN(new_n688));
  OR3_X1    g263(.A1(KEYINPUT88), .A2(G16), .A3(G23), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n688), .B(new_n689), .C1(G288), .C2(new_n684), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n691));
  INV_X1    g266(.A(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n684), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n684), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G6), .B(G305), .S(G16), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n694), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT34), .Z(new_n703));
  NAND3_X1  g278(.A1(new_n683), .A2(new_n687), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT36), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G26), .ZN(new_n707));
  OR2_X1    g282(.A1(G104), .A2(G2105), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n465), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI221_X1 g285(.A(new_n710), .B1(new_n709), .B2(new_n708), .C1(G116), .C2(new_n461), .ZN(new_n711));
  INV_X1    g286(.A(G140), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n468), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G128), .B2(new_n492), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n707), .B1(new_n714), .B2(new_n706), .ZN(new_n715));
  MUX2_X1   g290(.A(new_n707), .B(new_n715), .S(KEYINPUT28), .Z(new_n716));
  INV_X1    g291(.A(G2078), .ZN(new_n717));
  NOR2_X1   g292(.A1(G164), .A2(new_n706), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G27), .B2(new_n706), .ZN(new_n719));
  OAI22_X1  g294(.A1(new_n716), .A2(G2067), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n684), .A2(G4), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n592), .B2(new_n684), .ZN(new_n722));
  INV_X1    g297(.A(G1348), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT30), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n706), .B1(new_n725), .B2(G28), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT95), .Z(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n725), .B2(G28), .ZN(new_n728));
  NAND2_X1  g303(.A1(G171), .A2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G5), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n724), .B(new_n732), .C1(new_n731), .C2(new_n730), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n720), .B(new_n733), .C1(new_n717), .C2(new_n719), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G21), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G168), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(G1966), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT31), .B(G11), .ZN(new_n739));
  OR2_X1    g314(.A1(G29), .A2(G33), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n469), .A2(G139), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n471), .A2(G103), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT25), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n741), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n745), .B1(new_n741), .B2(new_n744), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n747), .A2(new_n748), .B1(new_n461), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n740), .B1(new_n750), .B2(new_n706), .ZN(new_n751));
  INV_X1    g326(.A(G2072), .ZN(new_n752));
  INV_X1    g327(.A(new_n615), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n751), .A2(new_n752), .B1(new_n753), .B2(G29), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n734), .A2(new_n738), .A3(new_n739), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n684), .A2(G19), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n547), .B2(new_n684), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(G1341), .ZN(new_n758));
  NOR2_X1   g333(.A1(G29), .A2(G32), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n471), .A2(G105), .ZN(new_n760));
  INV_X1    g335(.A(G141), .ZN(new_n761));
  INV_X1    g336(.A(G129), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n760), .B1(new_n468), .B2(new_n761), .C1(new_n485), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT93), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n768));
  OR3_X1    g343(.A1(new_n763), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n763), .B2(new_n767), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n759), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  NOR2_X1   g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n775), .A2(new_n776), .A3(G29), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n478), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT92), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G2084), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n716), .A2(G2067), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n779), .A2(G2084), .B1(new_n757), .B2(G1341), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n774), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G35), .ZN(new_n785));
  OAI21_X1  g360(.A(KEYINPUT96), .B1(new_n785), .B2(G29), .ZN(new_n786));
  OR3_X1    g361(.A1(new_n785), .A2(KEYINPUT96), .A3(G29), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n786), .B(new_n787), .C1(G162), .C2(new_n706), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G2090), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT97), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n791), .B1(new_n752), .B2(new_n751), .C1(G2090), .C2(new_n789), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n755), .A2(new_n758), .A3(new_n784), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n684), .A2(G20), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n560), .A2(new_n562), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n684), .ZN(new_n796));
  MUX2_X1   g371(.A(new_n794), .B(new_n796), .S(KEYINPUT23), .Z(new_n797));
  XOR2_X1   g372(.A(KEYINPUT98), .B(G1956), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n705), .A2(new_n793), .A3(new_n799), .ZN(G150));
  INV_X1    g375(.A(G150), .ZN(G311));
  AOI22_X1  g376(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(new_n510), .ZN(new_n803));
  INV_X1    g378(.A(G93), .ZN(new_n804));
  INV_X1    g379(.A(G55), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n513), .A2(new_n804), .B1(new_n515), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(G860), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT37), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n592), .A2(G559), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n803), .A2(new_n806), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n546), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT39), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n810), .B(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(G860), .ZN(G145));
  XNOR2_X1  g390(.A(new_n679), .B(new_n619), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n492), .A2(G130), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n469), .A2(G142), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT101), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(KEYINPUT101), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n821), .B(new_n822), .C1(G118), .C2(new_n461), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n818), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n484), .A2(G138), .A3(new_n461), .A4(new_n464), .ZN(new_n827));
  AOI211_X1 g402(.A(new_n826), .B(new_n498), .C1(new_n827), .C2(KEYINPUT4), .ZN(new_n828));
  AOI21_X1  g403(.A(KEYINPUT99), .B1(new_n495), .B2(new_n499), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n493), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n714), .ZN(new_n833));
  OAI211_X1 g408(.A(KEYINPUT100), .B(new_n493), .C1(new_n828), .C2(new_n829), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n833), .B1(new_n832), .B2(new_n834), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n825), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n750), .A2(new_n770), .A3(new_n769), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n750), .B1(new_n770), .B2(new_n769), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n500), .A2(new_n826), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n495), .A2(KEYINPUT99), .A3(new_n499), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT100), .B1(new_n843), .B2(new_n493), .ZN(new_n844));
  INV_X1    g419(.A(new_n834), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n714), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n824), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n837), .A2(new_n840), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n840), .B1(new_n837), .B2(new_n848), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n817), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n835), .A2(new_n836), .A3(new_n825), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n824), .B1(new_n846), .B2(new_n847), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n853), .A2(new_n854), .B1(new_n839), .B2(new_n838), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n837), .A2(new_n840), .A3(new_n848), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n816), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n851), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n615), .B(new_n487), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n851), .A2(new_n857), .A3(new_n852), .A4(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G160), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n478), .A3(new_n862), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT103), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n864), .A2(new_n869), .A3(new_n865), .A4(new_n866), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n868), .A2(KEYINPUT40), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT40), .B1(new_n868), .B2(new_n870), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(G395));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n592), .B1(G299), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n874), .B2(G299), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n795), .A2(KEYINPUT104), .A3(new_n592), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n876), .A2(KEYINPUT41), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT41), .B1(new_n876), .B2(new_n877), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n603), .B(new_n812), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n882), .A2(KEYINPUT42), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(G303), .B(KEYINPUT105), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G305), .ZN(new_n887));
  XNOR2_X1  g462(.A(G288), .B(new_n583), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n890), .A3(new_n887), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(KEYINPUT107), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT42), .B1(new_n882), .B2(new_n884), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n885), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n885), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(G868), .B2(new_n811), .ZN(G295));
  OAI21_X1  g476(.A(new_n900), .B1(G868), .B2(new_n811), .ZN(G331));
  XNOR2_X1  g477(.A(new_n812), .B(G301), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G168), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(G168), .ZN(new_n906));
  OAI22_X1  g481(.A1(new_n878), .A2(new_n879), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n883), .A3(new_n904), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(KEYINPUT108), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n895), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n907), .A2(KEYINPUT108), .A3(new_n894), .A4(new_n909), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n865), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n911), .A2(new_n915), .A3(new_n865), .A4(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(new_n913), .B2(KEYINPUT43), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n917), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n914), .A2(new_n919), .A3(KEYINPUT44), .A4(new_n916), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(G397));
  AOI21_X1  g498(.A(G1384), .B1(new_n832), .B2(new_n834), .ZN(new_n924));
  XNOR2_X1  g499(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G40), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n478), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT111), .ZN(new_n930));
  INV_X1    g505(.A(new_n771), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(G1996), .A3(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n714), .B(G2067), .Z(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n679), .B(new_n682), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n929), .A2(G1996), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n937), .A2(new_n931), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n932), .A2(new_n934), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n929), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n583), .B(G1986), .Z(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT126), .ZN(new_n943));
  INV_X1    g518(.A(G8), .ZN(new_n944));
  INV_X1    g519(.A(new_n928), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT116), .ZN(new_n946));
  AOI21_X1  g521(.A(G1384), .B1(new_n493), .B2(new_n500), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n925), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(KEYINPUT116), .A3(new_n925), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1384), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n830), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n737), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n948), .A2(KEYINPUT112), .A3(KEYINPUT50), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n947), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n830), .A2(new_n961), .A3(new_n953), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n781), .A3(new_n928), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n944), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(G168), .A2(new_n944), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT125), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n943), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n965), .ZN(new_n970));
  AOI21_X1  g545(.A(G1966), .B1(new_n952), .B2(new_n956), .ZN(new_n971));
  OAI21_X1  g546(.A(G8), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT125), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n967), .B(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n974), .A3(KEYINPUT126), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(new_n975), .A3(KEYINPUT51), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n968), .B1(new_n971), .B2(new_n970), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n943), .B(new_n978), .C1(new_n966), .C2(new_n968), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n830), .A2(new_n928), .A3(new_n953), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n982), .B(G8), .C1(new_n692), .C2(G288), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(KEYINPUT113), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(G288), .A2(new_n984), .A3(new_n692), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n985), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(G305), .B(KEYINPUT49), .ZN(new_n990));
  INV_X1    g565(.A(G1981), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n575), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n990), .B(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n982), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n944), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n989), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(G303), .A2(G8), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT55), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n963), .A2(new_n928), .A3(new_n964), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(G2090), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n924), .A2(KEYINPUT45), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1971), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(G8), .B(new_n1001), .C1(new_n1003), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1006), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n945), .B1(new_n954), .B2(KEYINPUT50), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(KEYINPUT50), .B2(new_n948), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(G2090), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n944), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n998), .B(new_n1007), .C1(new_n1012), .C2(new_n1001), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1002), .A2(KEYINPUT120), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n963), .A2(new_n1016), .A3(new_n928), .A4(new_n964), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1004), .A2(new_n717), .A3(new_n1005), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1018), .A2(new_n731), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n952), .A2(KEYINPUT53), .A3(new_n717), .A4(new_n956), .ZN(new_n1022));
  AOI21_X1  g597(.A(G301), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT62), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n976), .A2(new_n1024), .A3(new_n977), .A4(new_n979), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n981), .A2(new_n1014), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  OAI211_X1 g602(.A(G8), .B(G168), .C1(new_n970), .C2(new_n971), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT117), .Z(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1029), .B2(new_n1013), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1028), .B(KEYINPUT117), .ZN(new_n1031));
  OAI21_X1  g606(.A(G8), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1027), .B1(new_n1032), .B2(new_n1000), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1031), .A2(new_n1007), .A3(new_n998), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n997), .A2(new_n692), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1035), .A2(G288), .B1(G1981), .B2(G305), .ZN(new_n1036));
  XOR2_X1   g611(.A(new_n1036), .B(KEYINPUT115), .Z(new_n1037));
  AOI22_X1  g612(.A1(new_n1030), .A2(new_n1034), .B1(new_n996), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1007), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n998), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1026), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1021), .A2(G301), .A3(new_n1022), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n926), .A2(new_n1019), .A3(G2078), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n928), .A3(new_n1004), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1021), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT54), .B(new_n1042), .C1(new_n1045), .C2(G301), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1021), .A2(G301), .A3(new_n1044), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1023), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1046), .A2(new_n980), .A3(new_n1049), .A4(new_n1014), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT123), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n795), .B1(new_n1053), .B2(KEYINPUT57), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(KEYINPUT57), .ZN(new_n1055));
  XOR2_X1   g630(.A(new_n1054), .B(new_n1055), .Z(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT56), .B(G2072), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1004), .A2(new_n1005), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT119), .ZN(new_n1059));
  INV_X1    g634(.A(G1956), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1010), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1004), .A2(new_n1062), .A3(new_n1005), .A4(new_n1057), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1056), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1054), .B(new_n1055), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1066), .A2(new_n1061), .A3(new_n1059), .A4(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1052), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT124), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1051), .A2(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT124), .B(KEYINPUT61), .C1(new_n1072), .C2(new_n1052), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1348), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n982), .A2(G2067), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n602), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n592), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1074), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT121), .B(G1341), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT58), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1082), .A2(G1996), .B1(new_n995), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1086));
  NAND2_X1  g661(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1085), .A2(new_n547), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1085), .A2(new_n547), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(new_n1086), .ZN(new_n1090));
  NOR4_X1   g665(.A1(new_n1075), .A2(KEYINPUT60), .A3(new_n602), .A4(new_n1077), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1081), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1071), .A2(new_n1073), .A3(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1067), .B(new_n592), .C1(new_n1077), .C2(new_n1075), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1094), .A2(new_n1065), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1050), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n942), .B1(new_n1041), .B2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n929), .A2(G1986), .A3(G290), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT48), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n939), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n937), .B(KEYINPUT46), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n930), .B1(new_n931), .B2(new_n933), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1104));
  XNOR2_X1  g679(.A(new_n1103), .B(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n680), .A2(new_n682), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n932), .A2(new_n934), .A3(new_n938), .A4(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(G2067), .B2(new_n833), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1100), .B(new_n1105), .C1(new_n930), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1097), .A2(new_n1109), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g685(.A(G319), .ZN(new_n1112));
  NOR2_X1   g686(.A1(G229), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g687(.A1(G227), .A2(G401), .ZN(new_n1114));
  NAND4_X1  g688(.A1(new_n917), .A2(new_n867), .A3(new_n1113), .A4(new_n1114), .ZN(G225));
  INV_X1    g689(.A(G225), .ZN(G308));
endmodule


