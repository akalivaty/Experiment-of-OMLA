//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n643, new_n644,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(G319));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(KEYINPUT69), .B(G125), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n462), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT69), .B1(new_n471), .B2(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(G137), .ZN(new_n475));
  INV_X1    g050(.A(G101), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(new_n469), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n473), .A2(KEYINPUT70), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2105), .C1(new_n467), .C2(new_n472), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n471), .A2(KEYINPUT71), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n470), .B2(new_n462), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(new_n474), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  INV_X1    g063(.A(G100), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n489), .A2(new_n474), .A3(KEYINPUT72), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT72), .B1(new_n489), .B2(new_n474), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G112), .B2(new_n474), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n486), .A2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(G136), .B2(new_n494), .ZN(G162));
  NAND2_X1  g070(.A1(KEYINPUT4), .A2(G138), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n470), .B2(new_n462), .ZN(new_n497));
  AND2_X1   g072(.A1(G102), .A2(G2104), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n474), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n500), .B1(new_n470), .B2(new_n462), .ZN(new_n501));
  AND2_X1   g076(.A1(G114), .A2(G2104), .ZN(new_n502));
  OAI21_X1  g077(.A(G2105), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n474), .C1(new_n463), .C2(new_n464), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n499), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT73), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT73), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT74), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(new_n519), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT73), .A2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(KEYINPUT6), .A3(new_n527), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n524), .A2(new_n528), .A3(G50), .A4(G543), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT75), .B(G88), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n524), .A2(new_n528), .A3(new_n513), .A4(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(new_n529), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n518), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  OAI211_X1 g113(.A(KEYINPUT77), .B(new_n518), .C1(new_n533), .C2(new_n534), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  AND3_X1   g117(.A1(new_n524), .A2(new_n528), .A3(new_n513), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G89), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n517), .A2(KEYINPUT6), .B1(new_n520), .B2(new_n523), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n545), .A2(G51), .A3(G543), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n549));
  AND2_X1   g124(.A1(G63), .A2(G651), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n548), .A2(new_n549), .B1(new_n513), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n544), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n544), .A2(KEYINPUT78), .A3(new_n546), .A4(new_n551), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(G168));
  NAND2_X1  g131(.A1(new_n524), .A2(new_n528), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n510), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G52), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n543), .A2(G90), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n517), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(G301));
  INV_X1    g138(.A(G301), .ZN(G171));
  XOR2_X1   g139(.A(KEYINPUT79), .B(G43), .Z(new_n565));
  NAND2_X1  g140(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n543), .A2(G81), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n567), .B1(new_n566), .B2(new_n568), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n569), .A2(new_n570), .B1(new_n517), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  AND3_X1   g149(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G36), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G188));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n581));
  AND2_X1   g156(.A1(KEYINPUT5), .A2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(KEYINPUT5), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n511), .A2(KEYINPUT82), .A3(new_n512), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n580), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n543), .A2(G91), .ZN(new_n590));
  INV_X1    g165(.A(G53), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(KEYINPUT9), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(KEYINPUT9), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n545), .A2(G543), .A3(new_n593), .A4(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n524), .A2(new_n528), .A3(G543), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(new_n594), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n589), .A2(new_n590), .A3(new_n596), .A4(new_n598), .ZN(G299));
  INV_X1    g174(.A(G168), .ZN(G286));
  NAND2_X1  g175(.A1(new_n558), .A2(G49), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n543), .A2(G87), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(G288));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n511), .B2(new_n512), .ZN(new_n606));
  AND2_X1   g181(.A1(G48), .A2(G543), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n528), .B(new_n524), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n526), .A2(new_n527), .ZN(new_n609));
  INV_X1    g184(.A(G61), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n511), .B2(new_n512), .ZN(new_n611));
  AND2_X1   g186(.A1(G73), .A2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(G305));
  NAND2_X1  g189(.A1(new_n558), .A2(G47), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n543), .A2(G85), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n615), .B(new_n616), .C1(new_n517), .C2(new_n617), .ZN(G290));
  NAND2_X1  g193(.A1(G301), .A2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n543), .A2(G92), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT10), .Z(new_n621));
  NOR3_X1   g196(.A1(new_n582), .A2(new_n583), .A3(new_n581), .ZN(new_n622));
  AOI21_X1  g197(.A(KEYINPUT82), .B1(new_n511), .B2(new_n512), .ZN(new_n623));
  OAI21_X1  g198(.A(G66), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g200(.A1(G79), .A2(G543), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G66), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n584), .B2(new_n585), .ZN(new_n629));
  INV_X1    g204(.A(new_n626), .ZN(new_n630));
  OAI21_X1  g205(.A(KEYINPUT83), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n627), .A2(new_n631), .A3(G651), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n558), .A2(G54), .ZN(new_n633));
  AND3_X1   g208(.A1(new_n632), .A2(KEYINPUT84), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(KEYINPUT84), .B1(new_n632), .B2(new_n633), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n621), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT85), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n621), .B(new_n638), .C1(new_n634), .C2(new_n635), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n619), .B1(new_n640), .B2(G868), .ZN(G284));
  OAI21_X1  g216(.A(new_n619), .B1(new_n640), .B2(G868), .ZN(G321));
  NAND2_X1  g217(.A1(G286), .A2(G868), .ZN(new_n643));
  XNOR2_X1  g218(.A(G299), .B(KEYINPUT86), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(G868), .B2(new_n644), .ZN(G297));
  OAI21_X1  g220(.A(new_n643), .B1(G868), .B2(new_n644), .ZN(G280));
  INV_X1    g221(.A(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n640), .B1(new_n647), .B2(G860), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT87), .ZN(G148));
  OAI21_X1  g224(.A(KEYINPUT88), .B1(new_n573), .B2(G868), .ZN(new_n650));
  AOI21_X1  g225(.A(G559), .B1(new_n637), .B2(new_n639), .ZN(new_n651));
  INV_X1    g226(.A(G868), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  MUX2_X1   g228(.A(new_n650), .B(KEYINPUT88), .S(new_n653), .Z(G323));
  XNOR2_X1  g229(.A(G323), .B(KEYINPUT11), .ZN(G282));
  MUX2_X1   g230(.A(G99), .B(G111), .S(G2105), .Z(new_n656));
  AOI22_X1  g231(.A1(new_n487), .A2(G123), .B1(G2104), .B2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G135), .ZN(new_n658));
  INV_X1    g233(.A(new_n494), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(G2096), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT12), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT13), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT89), .ZN(new_n666));
  INV_X1    g241(.A(G2100), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(KEYINPUT13), .ZN(new_n669));
  OR4_X1    g244(.A1(KEYINPUT89), .A2(new_n668), .A3(G2100), .A4(new_n669), .ZN(new_n670));
  OAI22_X1  g245(.A1(new_n668), .A2(new_n669), .B1(KEYINPUT89), .B2(G2100), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n662), .A2(new_n670), .A3(new_n671), .ZN(G156));
  XOR2_X1   g247(.A(KEYINPUT15), .B(G2435), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2438), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2427), .ZN(new_n675));
  INV_X1    g250(.A(G2430), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(KEYINPUT14), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2451), .B(G2454), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2443), .B(G2446), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1341), .B(G1348), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  OAI21_X1  g262(.A(G14), .B1(new_n684), .B2(new_n685), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(G401));
  XNOR2_X1  g264(.A(G2072), .B(G2078), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT17), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2084), .B(G2090), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT91), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2067), .B(G2678), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT92), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n694), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(new_n693), .C1(new_n690), .C2(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n690), .A2(new_n694), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT18), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n696), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(new_n661), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G2100), .ZN(G227));
  XOR2_X1   g279(.A(G1971), .B(G1976), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT19), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1956), .B(G2474), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1961), .B(G1966), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT20), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n707), .A2(new_n708), .ZN(new_n714));
  INV_X1    g289(.A(new_n709), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n706), .B2(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n711), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1991), .B(G1996), .ZN(new_n722));
  XNOR2_X1  g297(.A(G1981), .B(G1986), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n721), .B(new_n724), .Z(G229));
  XOR2_X1   g300(.A(KEYINPUT31), .B(G11), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT101), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT30), .B(G28), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n660), .B2(new_n728), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n494), .A2(G139), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT25), .Z(new_n734));
  AOI22_X1  g309(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n734), .C1(new_n474), .C2(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G33), .B(new_n736), .S(G29), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G2072), .ZN(new_n738));
  NOR2_X1   g313(.A1(G27), .A2(G29), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G164), .B2(G29), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n738), .B1(G2078), .B2(new_n740), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n731), .B(new_n741), .C1(G2078), .C2(new_n740), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT95), .B(G16), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G19), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n573), .B2(new_n744), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G1341), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n728), .A2(G26), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  MUX2_X1   g324(.A(G104), .B(G116), .S(G2105), .Z(new_n750));
  AOI22_X1  g325(.A1(new_n487), .A2(G128), .B1(G2104), .B2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G140), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n659), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n749), .B1(new_n753), .B2(G29), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2067), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n737), .A2(G2072), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT98), .Z(new_n757));
  NAND4_X1  g332(.A1(new_n742), .A2(new_n747), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G16), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G5), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G171), .B2(new_n759), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(G1961), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n728), .A2(G32), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n487), .A2(G129), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT26), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  AND2_X1   g343(.A1(G105), .A2(G2104), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n767), .A2(new_n768), .B1(new_n474), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n494), .A2(G141), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n763), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n774), .A2(new_n775), .B1(G1961), .B2(new_n761), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n762), .B(new_n776), .C1(new_n774), .C2(new_n775), .ZN(new_n777));
  NOR2_X1   g352(.A1(G29), .A2(G35), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G162), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT29), .ZN(new_n780));
  INV_X1    g355(.A(G2084), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G34), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(G29), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n481), .B2(G29), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n780), .A2(G2090), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n743), .A2(G20), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT23), .ZN(new_n788));
  INV_X1    g363(.A(G299), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n759), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n777), .A2(new_n786), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n785), .A2(new_n781), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT100), .ZN(new_n795));
  NOR2_X1   g370(.A1(G16), .A2(G21), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G168), .B2(G16), .ZN(new_n797));
  INV_X1    g372(.A(G1966), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n795), .B(new_n799), .C1(new_n780), .C2(G2090), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n758), .A2(new_n793), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G4), .A2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n640), .B2(G16), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G1348), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(G1348), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n801), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(G25), .A2(G29), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n494), .A2(G131), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT94), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n474), .A2(G95), .ZN(new_n810));
  NAND2_X1  g385(.A1(G107), .A2(G2105), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n469), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n487), .B2(G119), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n807), .B1(new_n814), .B2(new_n728), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  MUX2_X1   g392(.A(G24), .B(G290), .S(new_n744), .Z(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(G1986), .Z(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G23), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT96), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G288), .B2(new_n759), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT33), .B(G1976), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(G6), .A2(G16), .ZN(new_n825));
  INV_X1    g400(.A(G305), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G16), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT32), .B(G1981), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n537), .A2(new_n539), .A3(new_n744), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n743), .A2(G22), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n830), .A2(G1971), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(G1971), .B1(new_n830), .B2(new_n831), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n824), .B(new_n829), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n817), .B(new_n819), .C1(KEYINPUT34), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT97), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n806), .B1(new_n839), .B2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(new_n806), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(G150));
  NAND2_X1  g420(.A1(new_n640), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(new_n517), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT102), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n558), .A2(G55), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n543), .A2(G93), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n572), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n850), .A2(KEYINPUT103), .A3(new_n853), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n849), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n853), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n855), .B1(new_n862), .B2(new_n572), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n847), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  AOI21_X1  g440(.A(G860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  INV_X1    g442(.A(new_n862), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G860), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(new_n753), .B(G164), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  MUX2_X1   g448(.A(G106), .B(G118), .S(G2105), .Z(new_n874));
  AOI22_X1  g449(.A1(new_n487), .A2(G130), .B1(G2104), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G142), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n659), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n664), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n814), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n878), .A2(new_n814), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n873), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n879), .A3(new_n872), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n773), .B(new_n736), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n882), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(G162), .B(new_n660), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n481), .B(KEYINPUT104), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(new_n893), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g473(.A1(G303), .A2(new_n826), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n901));
  XNOR2_X1  g476(.A(G288), .B(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G290), .ZN(new_n903));
  NAND2_X1  g478(.A1(G303), .A2(new_n826), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n900), .B2(new_n904), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g483(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n905), .ZN(new_n912));
  INV_X1    g487(.A(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n862), .A2(new_n572), .ZN(new_n915));
  INV_X1    g490(.A(new_n855), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n917), .A2(new_n651), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n651), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n636), .B(new_n789), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n918), .B2(new_n919), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n910), .B(new_n914), .C1(new_n927), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n910), .A2(new_n914), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n925), .A2(new_n926), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n928), .A4(new_n924), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(G868), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n930), .A2(KEYINPUT108), .A3(G868), .A4(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n868), .A2(new_n652), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(G295));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n941));
  NAND3_X1  g516(.A1(G168), .A2(new_n941), .A3(G171), .ZN(new_n942));
  NOR2_X1   g517(.A1(G286), .A2(KEYINPUT109), .ZN(new_n943));
  OAI21_X1  g518(.A(G301), .B1(G168), .B2(new_n941), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n863), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n863), .A2(new_n945), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n923), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n921), .A3(new_n947), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n912), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n895), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n912), .B1(new_n949), .B2(new_n950), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n949), .A2(new_n950), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n908), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n895), .A4(new_n951), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n954), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n955), .B1(new_n954), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT126), .ZN(new_n963));
  INV_X1    g538(.A(new_n773), .ZN(new_n964));
  INV_X1    g539(.A(G1996), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n753), .A2(G2067), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n753), .A2(G2067), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n773), .A2(G1996), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n966), .A2(new_n968), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n473), .A2(KEYINPUT70), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n477), .A2(new_n474), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT110), .B(G40), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n972), .A2(new_n480), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n507), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n971), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n814), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n816), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n984), .A2(new_n816), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n971), .A2(KEYINPUT111), .A3(new_n980), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n983), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  NOR2_X1   g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n980), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n507), .A2(KEYINPUT50), .A3(new_n976), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT50), .B1(new_n507), .B2(new_n976), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n997), .A2(G2084), .A3(new_n975), .ZN(new_n998));
  INV_X1    g573(.A(new_n975), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT45), .B1(new_n507), .B2(new_n976), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1966), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(G8), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT122), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(G168), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n554), .A2(KEYINPUT122), .A3(G8), .A4(new_n555), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(new_n1010), .A3(KEYINPUT51), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n979), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n798), .B1(new_n1014), .B2(new_n975), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n977), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n507), .A2(KEYINPUT50), .A3(new_n976), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n999), .A2(new_n1019), .A3(new_n781), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1006), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1012), .B1(new_n1021), .B2(new_n1009), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1009), .B1(new_n1003), .B2(new_n998), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1011), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1006), .B1(KEYINPUT113), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n537), .A2(new_n539), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1026), .A2(KEYINPUT113), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1029), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n537), .A2(new_n539), .A3(new_n1027), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT112), .B(G1971), .Z(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n1014), .B2(new_n975), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n999), .A2(new_n1019), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1006), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1033), .B(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n975), .A2(new_n977), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n1006), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT114), .B1(G305), .B2(G1981), .ZN(new_n1043));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n608), .A2(new_n1044), .A3(new_n613), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1047), .B(new_n1044), .C1(new_n608), .C2(new_n613), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT49), .B1(new_n1052), .B2(KEYINPUT116), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT115), .B1(KEYINPUT116), .B2(KEYINPUT49), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n1054), .B(new_n1048), .C1(new_n1045), .C2(new_n1043), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1042), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  INV_X1    g632(.A(new_n977), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(new_n478), .A3(new_n480), .A4(new_n974), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  OR2_X1    g635(.A1(G288), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1061), .A3(G8), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1042), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1056), .A2(new_n1057), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1048), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT116), .B1(new_n1067), .B2(KEYINPUT115), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1055), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1042), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1065), .B(new_n1063), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT117), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1040), .A2(new_n1066), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G2078), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n999), .A2(new_n1002), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n999), .A2(new_n1019), .ZN(new_n1078));
  INV_X1    g653(.A(G1961), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1076), .A2(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR4_X1   g655(.A1(new_n975), .A2(new_n1000), .A3(new_n1001), .A4(G2078), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT53), .ZN(new_n1082));
  AOI21_X1  g657(.A(G301), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1025), .A2(new_n1074), .A3(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1024), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT124), .B1(new_n1024), .B2(KEYINPUT62), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1089));
  AND3_X1   g664(.A1(G299), .A2(KEYINPUT119), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G299), .A2(new_n1089), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT119), .B1(G299), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1090), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1956), .B1(new_n999), .B2(new_n1019), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT120), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1014), .A2(new_n975), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1094), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n791), .B1(new_n997), .B2(new_n975), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1097), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n999), .A2(new_n1002), .A3(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1093), .A2(new_n1091), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1100), .B(new_n1102), .C1(new_n1103), .C2(new_n1090), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1099), .A2(new_n1104), .A3(KEYINPUT61), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1348), .B1(new_n999), .B2(new_n1019), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n975), .A2(G2067), .A3(new_n977), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1106), .A2(KEYINPUT60), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n635), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n632), .A2(KEYINPUT84), .A3(new_n633), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n638), .B1(new_n1111), .B2(new_n621), .ZN(new_n1112));
  INV_X1    g687(.A(new_n639), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1108), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1105), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G1348), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1107), .B1(new_n1078), .B2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1117), .A2(new_n637), .A3(new_n639), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1107), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1078), .A2(new_n1116), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n637), .A2(new_n639), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT60), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n999), .A2(new_n1002), .A3(new_n965), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT121), .B(new_n1124), .C1(new_n975), .C2(new_n977), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT121), .B1(new_n1059), .B2(new_n1124), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n573), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT59), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n573), .B(new_n1130), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1115), .A2(new_n1122), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1121), .A2(new_n1104), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1137), .A2(new_n1099), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1079), .B1(new_n997), .B2(new_n975), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n467), .A2(new_n472), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1142), .A2(KEYINPUT123), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(KEYINPUT123), .ZN(new_n1144));
  OAI21_X1  g719(.A(G2105), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AND4_X1   g720(.A1(KEYINPUT53), .A2(new_n973), .A3(G40), .A4(new_n1075), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1002), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1141), .B(new_n1147), .C1(new_n1081), .C2(KEYINPUT53), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(G171), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1140), .B1(new_n1083), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1080), .A2(G301), .A3(new_n1082), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1148), .A2(G171), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(KEYINPUT54), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(new_n1024), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(new_n1074), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1085), .A2(new_n1088), .B1(new_n1139), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1039), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G288), .A2(G1976), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1070), .A2(new_n1158), .B1(new_n1044), .B2(new_n826), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1072), .A2(new_n1157), .B1(new_n1159), .B2(new_n1071), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1021), .A2(G168), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1074), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1072), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1162), .A2(new_n1161), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1040), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1160), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n994), .B1(new_n1156), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n983), .A2(new_n989), .A3(new_n986), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n968), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n980), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT125), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(new_n1173), .A3(new_n980), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n968), .A2(new_n964), .A3(new_n969), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n980), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n980), .A2(new_n965), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT46), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT47), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1179), .B(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n980), .A2(new_n992), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT48), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n990), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1172), .A2(new_n1174), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n963), .B1(new_n1168), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1139), .A2(new_n1155), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1074), .A2(new_n1084), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1025), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1024), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1167), .A2(new_n1187), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n994), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n1172), .A2(new_n1174), .A3(new_n1184), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1197), .A2(new_n1198), .A3(KEYINPUT126), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1186), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g775(.A(G229), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n954), .A2(new_n959), .ZN(new_n1203));
  NOR2_X1   g777(.A1(G227), .A2(new_n460), .ZN(new_n1204));
  OAI21_X1  g778(.A(new_n1204), .B1(new_n687), .B2(new_n688), .ZN(new_n1205));
  XNOR2_X1  g779(.A(new_n1205), .B(KEYINPUT127), .ZN(new_n1206));
  AND4_X1   g780(.A1(new_n1202), .A2(new_n1203), .A3(new_n897), .A4(new_n1206), .ZN(G308));
  NAND4_X1  g781(.A1(new_n1203), .A2(new_n1206), .A3(new_n1202), .A4(new_n897), .ZN(G225));
endmodule


