//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n591, new_n592, new_n593, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n628, new_n629, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n472), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n466), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n469), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n476), .A2(new_n483), .ZN(G160));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  AND4_X1   g062(.A1(G2105), .A2(new_n473), .A3(new_n469), .A4(new_n468), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  OAI221_X1 g065(.A(new_n486), .B1(new_n474), .B2(new_n487), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n471), .B1(KEYINPUT68), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT69), .ZN(new_n499));
  INV_X1    g074(.A(new_n493), .ZN(new_n500));
  OAI21_X1  g075(.A(G2105), .B1(new_n496), .B2(G114), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n494), .A2(KEYINPUT68), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n499), .A2(new_n505), .B1(new_n488), .B2(G126), .ZN(new_n506));
  INV_X1    g081(.A(G138), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(G2105), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n473), .A2(new_n468), .A3(new_n508), .A4(new_n469), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n469), .A2(new_n478), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(new_n508), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n520), .A2(new_n521), .B1(G50), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(new_n524), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(new_n517), .A3(KEYINPUT70), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G88), .ZN(new_n537));
  OAI21_X1  g112(.A(KEYINPUT71), .B1(new_n518), .B2(new_n519), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n526), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(G166));
  NAND3_X1  g115(.A1(new_n533), .A2(G89), .A3(new_n535), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n534), .A2(G51), .A3(G543), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n528), .A2(new_n527), .ZN(new_n547));
  NAND2_X1  g122(.A1(G63), .A2(G651), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n517), .A2(KEYINPUT72), .A3(G63), .A4(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n541), .A2(new_n545), .A3(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n547), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G651), .B1(G52), .B2(new_n525), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT73), .B(G90), .Z(new_n558));
  NAND3_X1  g133(.A1(new_n533), .A2(new_n535), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n547), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n564), .A2(G651), .B1(G43), .B2(new_n525), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n533), .A2(G81), .A3(new_n535), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n547), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n533), .A2(new_n535), .ZN(new_n578));
  INV_X1    g153(.A(G91), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n534), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G53), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n582), .A2(new_n583), .B1(KEYINPUT74), .B2(KEYINPUT9), .ZN(new_n584));
  AND2_X1   g159(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n585));
  NOR2_X1   g160(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n525), .B(G53), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT75), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n584), .A2(KEYINPUT75), .A3(new_n587), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n581), .B1(new_n588), .B2(new_n589), .ZN(G299));
  NAND2_X1  g165(.A1(new_n539), .A2(KEYINPUT76), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n526), .A2(new_n537), .A3(new_n592), .A4(new_n538), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(G303));
  NAND2_X1  g169(.A1(new_n536), .A2(G87), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n517), .A2(G74), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n525), .B2(G49), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(new_n536), .A2(G86), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n547), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G48), .B2(new_n525), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  NOR3_X1   g182(.A1(new_n607), .A2(KEYINPUT78), .A3(new_n519), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G47), .B2(new_n525), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n536), .A2(G85), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT78), .B1(new_n607), .B2(new_n519), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n547), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n525), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n536), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n578), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n618), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n613), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n613), .B1(new_n623), .B2(G868), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(new_n588), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n584), .A2(KEYINPUT75), .A3(new_n587), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n580), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n626), .B1(new_n629), .B2(G868), .ZN(G297));
  OAI21_X1  g205(.A(new_n626), .B1(new_n629), .B2(G868), .ZN(G280));
  NAND2_X1  g206(.A1(new_n619), .A2(new_n622), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n617), .ZN(new_n633));
  INV_X1    g208(.A(G860), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT79), .B(G559), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT80), .ZN(G148));
  INV_X1    g212(.A(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n567), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n633), .A2(new_n635), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n638), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g217(.A1(new_n511), .A2(new_n465), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  OR2_X1    g221(.A1(G99), .A2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n647), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n648));
  INV_X1    g223(.A(G123), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n489), .B2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n474), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(G135), .B2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(G2096), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n652), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G2096), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n646), .A2(new_n654), .A3(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1341), .B(G1348), .Z(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT82), .ZN(new_n669));
  XOR2_X1   g244(.A(G2451), .B(G2454), .Z(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(new_n671));
  OR2_X1    g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n671), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n672), .A2(G14), .A3(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(G2067), .B(G2678), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT83), .ZN(new_n676));
  NOR2_X1   g251(.A1(G2072), .A2(G2078), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n444), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2084), .B(G2090), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n678), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT85), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(KEYINPUT85), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(new_n676), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n678), .B(KEYINPUT17), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n686), .B(new_n679), .C1(new_n676), .C2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n679), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n687), .A2(new_n676), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n682), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(new_n653), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT86), .B(G2100), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G227));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1956), .B(G2474), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1961), .B(G1966), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT20), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n698), .B(new_n699), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n702), .B(new_n703), .C1(new_n697), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(G1981), .B(G1986), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(G229));
  NOR2_X1   g286(.A1(G6), .A2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n604), .B(KEYINPUT77), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(G16), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT32), .B(G1981), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G22), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G166), .B2(new_n717), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1971), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(G23), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n595), .A2(new_n597), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n717), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT33), .B(G1976), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR3_X1   g300(.A1(new_n716), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G25), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n651), .A2(G131), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n488), .A2(G119), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n471), .A2(G107), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n731), .B1(new_n737), .B2(new_n730), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT35), .B(G1991), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n738), .B(new_n739), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n717), .A2(G24), .ZN(new_n741));
  INV_X1    g316(.A(G290), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n717), .ZN(new_n743));
  INV_X1    g318(.A(G1986), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n728), .A2(new_n729), .A3(new_n740), .A4(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n747));
  OR3_X1    g322(.A1(new_n746), .A2(KEYINPUT88), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT88), .B(KEYINPUT36), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G140), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n474), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n755));
  INV_X1    g330(.A(G116), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(G2105), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n488), .B2(G128), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G29), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT90), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n730), .A2(G26), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT28), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT91), .B(G2067), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT26), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n769), .A2(new_n770), .B1(G105), .B2(new_n465), .ZN(new_n771));
  INV_X1    g346(.A(G141), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n488), .A2(KEYINPUT95), .A3(G129), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(KEYINPUT95), .B1(new_n488), .B2(G129), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n771), .B1(new_n772), .B2(new_n474), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(new_n730), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n730), .B2(G32), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  NOR2_X1   g357(.A1(G4), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n623), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n781), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G27), .A2(G29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G164), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT96), .B(G2078), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT97), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G1348), .B2(new_n784), .ZN(new_n792));
  NAND2_X1  g367(.A1(G160), .A2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT24), .B(G34), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(new_n730), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT92), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G2084), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n730), .A2(G33), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n651), .A2(G139), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT25), .ZN(new_n804));
  NAND2_X1  g379(.A1(G115), .A2(G2104), .ZN(new_n805));
  INV_X1    g380(.A(G127), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n479), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n804), .B1(G2105), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n801), .B1(new_n809), .B2(G29), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n442), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT94), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n779), .B2(new_n780), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n786), .A2(new_n792), .A3(new_n800), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT31), .B(G11), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT30), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(G28), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n730), .B1(new_n816), .B2(G28), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n815), .B1(new_n817), .B2(new_n818), .C1(new_n655), .C2(new_n730), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n717), .A2(G21), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G168), .B2(new_n717), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1966), .ZN(new_n822));
  INV_X1    g397(.A(G1961), .ZN(new_n823));
  NOR2_X1   g398(.A1(G171), .A2(new_n717), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G5), .B2(new_n717), .ZN(new_n825));
  AOI211_X1 g400(.A(new_n819), .B(new_n822), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n717), .A2(G20), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT23), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n629), .B2(new_n717), .ZN(new_n829));
  INV_X1    g404(.A(G1956), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n730), .A2(G35), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G162), .B2(new_n730), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT29), .B(G2090), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n798), .B2(new_n797), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n825), .A2(new_n823), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n568), .A2(G16), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G16), .B2(G19), .ZN(new_n839));
  INV_X1    g414(.A(G1341), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n810), .A2(new_n442), .ZN(new_n843));
  NOR4_X1   g418(.A1(new_n837), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n826), .A2(new_n831), .A3(new_n836), .A4(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n766), .A2(new_n814), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n748), .A2(new_n750), .A3(new_n846), .ZN(G150));
  INV_X1    g422(.A(G150), .ZN(G311));
  NAND2_X1  g423(.A1(new_n623), .A2(G559), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT38), .Z(new_n850));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n547), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n519), .B1(new_n853), .B2(KEYINPUT98), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(KEYINPUT98), .B2(new_n853), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n533), .A2(G93), .A3(new_n535), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n525), .A2(G55), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n856), .A2(KEYINPUT99), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT99), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n567), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n568), .B(new_n855), .C1(new_n858), .C2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n850), .B(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n634), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n860), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  NAND2_X1  g445(.A1(new_n488), .A2(G130), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  INV_X1    g447(.A(G118), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n872), .A2(KEYINPUT102), .B1(new_n873), .B2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(KEYINPUT102), .B2(new_n872), .ZN(new_n875));
  INV_X1    g450(.A(G142), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n871), .B(new_n875), .C1(new_n876), .C2(new_n474), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(new_n644), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n737), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n759), .B(new_n515), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n776), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n809), .A2(KEYINPUT101), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n809), .B(KEYINPUT101), .Z(new_n884));
  AND2_X1   g459(.A1(new_n880), .A2(new_n777), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n880), .A2(new_n777), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n879), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(new_n879), .A3(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n890), .A2(new_n889), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G160), .B(KEYINPUT100), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n491), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(new_n652), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n652), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n898), .B(KEYINPUT105), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n890), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n888), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n883), .A2(new_n887), .A3(KEYINPUT104), .A4(new_n879), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n901), .A2(new_n903), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n900), .A4(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n900), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n891), .A2(new_n892), .B1(new_n897), .B2(new_n896), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n907), .A2(new_n911), .ZN(G395));
  NAND2_X1  g487(.A1(new_n860), .A2(new_n638), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n863), .B(new_n640), .Z(new_n914));
  NAND2_X1  g489(.A1(G299), .A2(new_n623), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n633), .A2(new_n629), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n633), .A2(new_n629), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT106), .B1(G299), .B2(new_n623), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n919), .A2(new_n920), .A3(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n915), .ZN(new_n922));
  XOR2_X1   g497(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n923));
  OAI22_X1  g498(.A1(new_n921), .A2(KEYINPUT41), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n917), .B1(new_n914), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT42), .ZN(new_n926));
  NAND2_X1  g501(.A1(G305), .A2(G290), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n713), .A2(new_n742), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n722), .A2(KEYINPUT108), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n930));
  NAND2_X1  g505(.A1(G288), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(G166), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n539), .A3(new_n931), .ZN(new_n934));
  AND4_X1   g509(.A1(new_n927), .A2(new_n928), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n927), .A2(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n926), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n913), .B1(new_n939), .B2(new_n638), .ZN(G295));
  OAI21_X1  g515(.A(new_n913), .B1(new_n939), .B2(new_n638), .ZN(G331));
  NAND2_X1  g516(.A1(new_n542), .A2(new_n544), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n549), .B2(new_n550), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n943), .A2(new_n541), .B1(new_n559), .B2(new_n557), .ZN(new_n944));
  NOR2_X1   g519(.A1(G286), .A2(G301), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n861), .A2(new_n862), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT109), .ZN(new_n948));
  INV_X1    g523(.A(new_n946), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n863), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n861), .A2(new_n946), .A3(new_n951), .A4(new_n862), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n922), .A2(new_n923), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT41), .A4(new_n915), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n950), .A2(new_n922), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n957), .A2(KEYINPUT110), .B1(new_n947), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n953), .A2(new_n956), .A3(new_n961), .ZN(new_n962));
  AOI211_X1 g537(.A(KEYINPUT111), .B(new_n937), .C1(new_n960), .C2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(KEYINPUT110), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(new_n947), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n967), .B2(new_n938), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n950), .A2(new_n947), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n924), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n948), .A2(new_n952), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n937), .B(new_n971), .C1(new_n972), .C2(new_n958), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n900), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n973), .A2(new_n977), .A3(new_n900), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n972), .B2(new_n958), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n938), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n978), .B1(new_n963), .B2(new_n968), .ZN(new_n984));
  INV_X1    g559(.A(new_n980), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n985), .B2(new_n974), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n983), .B1(new_n987), .B2(new_n976), .ZN(new_n988));
  AOI211_X1 g563(.A(KEYINPUT112), .B(KEYINPUT44), .C1(new_n984), .C2(new_n986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(G397));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n488), .A2(G126), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n498), .A2(KEYINPUT69), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n503), .A2(new_n504), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n514), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n991), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT113), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n506), .B2(new_n514), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n651), .A2(G137), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT114), .B(G40), .Z(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1004), .A2(new_n482), .A3(new_n466), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1996), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(new_n776), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1008), .B(KEYINPUT116), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n759), .B(G2067), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n777), .A2(new_n1009), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1011), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n737), .B(new_n739), .Z(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1008), .A2(new_n744), .A3(new_n742), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1008), .A2(G1986), .A3(G290), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT115), .Z(new_n1023));
  AND2_X1   g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n591), .A2(G8), .A3(new_n593), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n591), .A2(KEYINPUT55), .A3(G8), .A4(new_n593), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1971), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1007), .B1(new_n997), .B2(new_n1002), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT45), .B(new_n991), .C1(new_n995), .C2(new_n996), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT117), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n999), .A2(new_n1034), .A3(KEYINPUT45), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n476), .A2(new_n483), .A3(new_n1005), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n999), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G2090), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1030), .A2(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1029), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1036), .A2(new_n1030), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(G8), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  INV_X1    g626(.A(G1981), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n599), .A2(new_n1052), .A3(new_n603), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n599), .B2(new_n603), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1055), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(KEYINPUT49), .A3(new_n1053), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1044), .B1(new_n1037), .B2(new_n999), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n722), .A2(G1976), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1060), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1045), .A2(new_n1050), .A3(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT125), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1033), .A2(new_n1035), .A3(KEYINPUT53), .A4(new_n443), .ZN(new_n1071));
  INV_X1    g646(.A(G40), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n481), .A2(KEYINPUT123), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n471), .B1(new_n481), .B2(KEYINPUT123), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1072), .B(new_n476), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1003), .A2(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1076), .A2(KEYINPUT124), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(KEYINPUT124), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1071), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1036), .B2(G2078), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n999), .A2(new_n1038), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n1037), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n823), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(G171), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1088), .A2(new_n1080), .A3(G2078), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1081), .A2(G301), .A3(new_n1085), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1087), .B(KEYINPUT54), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G171), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1079), .B2(new_n1090), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G168), .A2(new_n1044), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1041), .A2(new_n798), .ZN(new_n1096));
  INV_X1    g671(.A(G1966), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1088), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1095), .B1(new_n1099), .B2(G8), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1095), .B2(KEYINPUT122), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1100), .A2(new_n1102), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1102), .ZN(new_n1104));
  OAI211_X1 g679(.A(G8), .B(new_n1104), .C1(new_n1099), .C2(G286), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1093), .A2(new_n1094), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1070), .A2(new_n1091), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n584), .A2(new_n587), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n581), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n629), .A2(KEYINPUT57), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1084), .A2(new_n830), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1084), .A2(KEYINPUT119), .A3(new_n830), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  AND4_X1   g694(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1113), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1112), .B(new_n1120), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1108), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1117), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT119), .B1(new_n1084), .B2(new_n830), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1121), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1112), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1118), .A2(new_n1113), .A3(new_n1121), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(KEYINPUT61), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1037), .A2(new_n999), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT58), .B(G1341), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1036), .B2(G1996), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n568), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT59), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1124), .A2(new_n1130), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT121), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1124), .A2(new_n1130), .A3(new_n1139), .A4(new_n1136), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1131), .A2(G2067), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n782), .B2(new_n1084), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT60), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(new_n623), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(KEYINPUT60), .B2(new_n1142), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1138), .A2(new_n1140), .A3(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1142), .A2(new_n633), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1129), .B1(new_n1122), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1107), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1099), .A2(new_n1095), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1105), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1103), .A2(KEYINPUT62), .A3(new_n1105), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1092), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1070), .A3(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1060), .A2(new_n1064), .A3(new_n722), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1059), .B1(new_n1159), .B2(new_n1054), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1050), .B2(new_n1067), .ZN(new_n1161));
  AOI211_X1 g736(.A(new_n1044), .B(G286), .C1(new_n1096), .C2(new_n1098), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1045), .A2(new_n1068), .A3(new_n1162), .A4(new_n1050), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1048), .A2(G8), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1067), .B1(new_n1166), .B2(new_n1029), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1167), .A2(KEYINPUT63), .A3(new_n1050), .A4(new_n1162), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1161), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1169), .A2(KEYINPUT118), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n1171));
  AOI211_X1 g746(.A(new_n1171), .B(new_n1161), .C1(new_n1165), .C2(new_n1168), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1158), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1024), .B1(new_n1149), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1012), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n732), .A2(new_n736), .A3(new_n739), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1016), .A2(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n759), .A2(G2067), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1175), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1012), .B1(new_n776), .B2(new_n1013), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1010), .B(KEYINPUT46), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT47), .Z(new_n1183));
  XNOR2_X1  g758(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1184));
  AOI211_X1 g759(.A(new_n1179), .B(new_n1183), .C1(new_n1019), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1174), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g761(.A1(new_n899), .A2(new_n900), .A3(new_n906), .ZN(new_n1188));
  NOR2_X1   g762(.A1(G227), .A2(new_n462), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n1190));
  XNOR2_X1  g764(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  NOR2_X1   g765(.A1(G229), .A2(G401), .ZN(new_n1192));
  AND2_X1   g766(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n1188), .A2(new_n987), .A3(new_n1193), .ZN(G308));
  OAI211_X1 g768(.A(new_n1193), .B(new_n987), .C1(new_n910), .C2(new_n909), .ZN(G225));
endmodule


