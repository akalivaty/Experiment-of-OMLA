//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  OAI21_X1  g001(.A(G214), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n189), .A2(new_n191), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT82), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n190), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(G143), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n196), .A2(new_n197), .A3(new_n198), .A4(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n193), .A2(new_n195), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n191), .A2(new_n189), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT82), .B1(new_n206), .B2(G125), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n200), .A2(new_n201), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT64), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n198), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n203), .B1(new_n207), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G224), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G953), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G110), .B(G122), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT65), .B1(new_n223), .B2(G116), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  INV_X1    g039(.A(G116), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G119), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n226), .A2(G119), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(KEYINPUT5), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G113), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT5), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(G107), .ZN(new_n238));
  INV_X1    g052(.A(G107), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT3), .A3(G104), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G101), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT77), .B1(new_n239), .B2(G104), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT77), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n237), .A3(G107), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n241), .A2(new_n242), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n237), .A2(G107), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n239), .A2(G104), .ZN(new_n248));
  OAI21_X1  g062(.A(G101), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n232), .A2(KEYINPUT2), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT2), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G113), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n228), .A2(new_n230), .A3(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n235), .A2(new_n246), .A3(new_n249), .A4(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n238), .A2(new_n240), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n243), .A2(new_n245), .ZN(new_n257));
  OAI21_X1  g071(.A(G101), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n246), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n260), .B(G101), .C1(new_n256), .C2(new_n257), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n253), .B1(new_n228), .B2(new_n230), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n228), .A2(new_n230), .A3(new_n253), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n222), .B(new_n255), .C1(new_n259), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n220), .A2(KEYINPUT7), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n203), .B(new_n266), .C1(new_n207), .C2(new_n216), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n221), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n234), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT83), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n269), .B1(new_n231), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n270), .B2(new_n231), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n246), .A2(new_n249), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n274), .A3(new_n254), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n235), .A2(new_n254), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n222), .B(KEYINPUT8), .Z(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n268), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n255), .B1(new_n259), .B2(new_n264), .ZN(new_n283));
  INV_X1    g097(.A(new_n222), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT6), .A3(new_n265), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n217), .B(new_n220), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n283), .A2(new_n288), .A3(new_n284), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n282), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n291), .B1(new_n282), .B2(new_n290), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n188), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n291), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n221), .A2(new_n265), .A3(new_n267), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n279), .B1(new_n275), .B2(new_n277), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n297), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n282), .A2(new_n290), .A3(new_n291), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT84), .A3(new_n188), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT9), .B(G234), .ZN(new_n307));
  INV_X1    g121(.A(G217), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n307), .A2(new_n308), .A3(G953), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n190), .A2(G128), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT86), .B1(new_n189), .B2(G143), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT86), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n190), .A3(G128), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G134), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G116), .B(G122), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT14), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n226), .A2(KEYINPUT14), .A3(G122), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(KEYINPUT87), .A3(G107), .A4(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n323));
  INV_X1    g137(.A(G122), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G116), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n226), .A2(G122), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n325), .A2(new_n326), .A3(new_n319), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(G107), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n318), .A2(new_n239), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n317), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n318), .A2(new_n239), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n333), .A2(new_n331), .B1(new_n315), .B2(new_n316), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT13), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT13), .B1(new_n312), .B2(new_n314), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n335), .A2(new_n336), .A3(new_n311), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n334), .B1(new_n337), .B2(new_n316), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT88), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n332), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n332), .B2(new_n338), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n310), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n342), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n309), .A3(new_n340), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n345), .A3(new_n299), .ZN(new_n346));
  INV_X1    g160(.A(G478), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(KEYINPUT15), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n343), .A2(new_n345), .A3(new_n299), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n353));
  XNOR2_X1  g167(.A(G113), .B(G122), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(new_n237), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n198), .A2(KEYINPUT16), .A3(G140), .ZN(new_n356));
  XNOR2_X1  g170(.A(G125), .B(G140), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(KEYINPUT16), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G146), .ZN(new_n359));
  INV_X1    g173(.A(G140), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G125), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n198), .A2(G140), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT19), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT19), .B1(new_n361), .B2(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n192), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G131), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  AOI21_X1  g181(.A(G143), .B1(new_n367), .B2(G214), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(G143), .A3(G214), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n370), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n372), .A2(new_n368), .A3(G131), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n359), .B(new_n365), .C1(new_n371), .C2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n357), .B(new_n192), .ZN(new_n375));
  OAI211_X1 g189(.A(KEYINPUT18), .B(G131), .C1(new_n372), .C2(new_n368), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT18), .A2(G131), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n369), .A2(new_n370), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n355), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n381));
  INV_X1    g195(.A(new_n356), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n361), .A2(new_n362), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT16), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n192), .ZN(new_n386));
  OAI211_X1 g200(.A(KEYINPUT17), .B(G131), .C1(new_n372), .C2(new_n368), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n386), .A2(new_n359), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G131), .B1(new_n372), .B2(new_n368), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n369), .A2(new_n366), .A3(new_n370), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT17), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n381), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n380), .B1(new_n393), .B2(new_n355), .ZN(new_n394));
  OR2_X1    g208(.A1(G475), .A2(G902), .ZN(new_n395));
  OAI211_X1 g209(.A(KEYINPUT85), .B(new_n353), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n392), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n386), .A2(new_n359), .A3(new_n387), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n355), .B(new_n379), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n392), .A2(new_n386), .A3(new_n359), .A4(new_n387), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n355), .B1(new_n401), .B2(new_n379), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n299), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G475), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n374), .A2(new_n379), .ZN(new_n405));
  INV_X1    g219(.A(new_n355), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n395), .B1(new_n407), .B2(new_n399), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT20), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI211_X1 g224(.A(KEYINPUT85), .B(new_n395), .C1(new_n407), .C2(new_n399), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n396), .B(new_n404), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(G234), .A2(G237), .ZN(new_n413));
  INV_X1    g227(.A(G953), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(G952), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(G902), .A3(G953), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT21), .B(G898), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n352), .A2(new_n412), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n296), .A2(new_n306), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G221), .B1(new_n307), .B2(G902), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT75), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT80), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT11), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n316), .B2(G137), .ZN(new_n429));
  INV_X1    g243(.A(G137), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(KEYINPUT11), .A3(G134), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n316), .A2(G137), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G131), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n429), .A2(new_n431), .A3(new_n366), .A4(new_n432), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT79), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n202), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n209), .A2(KEYINPUT79), .A3(new_n199), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n196), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n246), .A3(new_n249), .ZN(new_n441));
  INV_X1    g255(.A(new_n206), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n273), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n436), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n426), .A2(KEYINPUT80), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n427), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n206), .B1(new_n246), .B2(new_n249), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n274), .B2(new_n440), .ZN(new_n448));
  OAI211_X1 g262(.A(KEYINPUT80), .B(new_n426), .C1(new_n448), .C2(new_n436), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT10), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n442), .A2(new_n451), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n441), .A2(new_n451), .B1(new_n274), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n261), .A2(new_n211), .A3(new_n215), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n259), .A2(new_n454), .A3(KEYINPUT78), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT78), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n211), .A2(new_n215), .ZN(new_n457));
  INV_X1    g271(.A(new_n257), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n242), .B1(new_n458), .B2(new_n241), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n459), .B2(new_n260), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n246), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n436), .B(new_n453), .C1(new_n455), .C2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G140), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n414), .A2(G227), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n464), .B(new_n465), .Z(new_n466));
  NAND3_X1  g280(.A1(new_n450), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT81), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n466), .ZN(new_n470));
  INV_X1    g284(.A(new_n463), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT78), .B1(new_n259), .B2(new_n454), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n460), .A2(new_n456), .A3(new_n461), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n436), .B1(new_n474), .B2(new_n453), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n470), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n450), .A2(new_n463), .A3(KEYINPUT81), .A4(new_n466), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n469), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G469), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n478), .A2(new_n479), .A3(new_n299), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n453), .B1(new_n455), .B2(new_n462), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n434), .A2(new_n435), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n466), .A3(new_n463), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n450), .A2(new_n463), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n466), .B(KEYINPUT76), .Z(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n479), .B1(new_n487), .B2(new_n299), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n425), .B1(new_n480), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n187), .B1(new_n422), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT84), .B1(new_n305), .B2(new_n188), .ZN(new_n491));
  INV_X1    g305(.A(new_n188), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n295), .B(new_n492), .C1(new_n303), .C2(new_n304), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n478), .A2(new_n479), .A3(new_n299), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n486), .B1(new_n450), .B2(new_n463), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n471), .A2(new_n475), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(new_n466), .ZN(new_n498));
  OAI21_X1  g312(.A(G469), .B1(new_n498), .B2(G902), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n424), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n494), .A2(KEYINPUT89), .A3(new_n500), .A4(new_n421), .ZN(new_n501));
  NOR2_X1   g315(.A1(G472), .A2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT32), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n482), .A2(new_n211), .A3(new_n215), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n263), .A2(new_n262), .ZN(new_n507));
  INV_X1    g321(.A(new_n432), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n316), .A2(G137), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n206), .A2(new_n435), .A3(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n507), .B1(new_n506), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT28), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT66), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(KEYINPUT66), .B(KEYINPUT28), .C1(new_n512), .C2(new_n513), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT28), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n367), .A2(G210), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT27), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(G101), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n507), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n506), .A2(new_n529), .A3(new_n511), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n529), .B1(new_n506), .B2(new_n511), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n525), .A3(new_n518), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT31), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n511), .B1(new_n436), .B2(new_n457), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT30), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n530), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n512), .B1(new_n538), .B2(new_n528), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT31), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n540), .A3(new_n525), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n505), .B1(new_n527), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n536), .A2(new_n528), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(new_n518), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n513), .A2(KEYINPUT67), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT28), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n520), .A2(KEYINPUT29), .A3(new_n525), .ZN(new_n549));
  AOI21_X1  g363(.A(G902), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n526), .B1(new_n519), .B2(new_n518), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n516), .A2(new_n517), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT29), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n539), .B2(new_n525), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G472), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n540), .B1(new_n539), .B2(new_n525), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n507), .B1(new_n537), .B2(new_n530), .ZN(new_n558));
  NOR4_X1   g372(.A1(new_n558), .A2(KEYINPUT31), .A3(new_n526), .A4(new_n512), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n521), .A2(new_n526), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n503), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n543), .B(new_n556), .C1(new_n562), .C2(KEYINPUT32), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n308), .B1(G234), .B2(new_n299), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT23), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(KEYINPUT69), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n189), .A2(G119), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n223), .A2(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n223), .A2(G128), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT69), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT23), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n565), .A2(KEYINPUT69), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G110), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT68), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n223), .B2(G128), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n189), .A2(KEYINPUT68), .A3(G119), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n567), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(KEYINPUT24), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT24), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G110), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n577), .A2(new_n587), .A3(KEYINPUT70), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT70), .ZN(new_n589));
  AOI21_X1  g403(.A(G110), .B1(new_n569), .B2(new_n574), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT68), .B1(new_n189), .B2(G119), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n578), .A2(new_n223), .A3(G128), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n585), .B1(new_n593), .B2(new_n567), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n589), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n383), .A2(G146), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n358), .B2(G146), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n588), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n386), .A2(new_n359), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n593), .A2(new_n567), .A3(new_n585), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n569), .A2(new_n574), .A3(G110), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n414), .A2(G221), .A3(G234), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT71), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT22), .B(G137), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n598), .A2(new_n602), .A3(new_n607), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT25), .B1(new_n611), .B2(new_n299), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n598), .A2(new_n602), .A3(new_n607), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n607), .B1(new_n598), .B2(new_n602), .ZN(new_n614));
  OAI211_X1 g428(.A(KEYINPUT25), .B(new_n299), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n564), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT73), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n564), .A2(G902), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT72), .Z(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n611), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n564), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n299), .B1(new_n613), .B2(new_n614), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT25), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n624), .B1(new_n627), .B2(new_n615), .ZN(new_n628));
  INV_X1    g442(.A(new_n622), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT73), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n563), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n632), .A2(KEYINPUT74), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(KEYINPUT74), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n490), .B(new_n501), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  NAND3_X1  g450(.A1(new_n561), .A2(new_n541), .A3(new_n535), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n299), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n562), .B1(new_n638), .B2(G472), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n500), .A2(new_n639), .A3(new_n631), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n420), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n305), .A2(new_n642), .A3(new_n188), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n347), .A2(G902), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT33), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n309), .B1(new_n344), .B2(new_n340), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n341), .A2(new_n310), .A3(new_n342), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT33), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT90), .B(G478), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n346), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n412), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n643), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n641), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT91), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT34), .B(G104), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  AOI21_X1  g474(.A(new_n412), .B1(new_n349), .B2(new_n351), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n643), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n641), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  OAI21_X1  g480(.A(KEYINPUT92), .B1(new_n607), .B2(KEYINPUT36), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n607), .A2(KEYINPUT92), .A3(KEYINPUT36), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT93), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n669), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT93), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n672), .A3(new_n667), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n603), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n670), .A2(new_n673), .A3(new_n602), .A4(new_n598), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n676), .A3(new_n621), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n617), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n639), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n501), .A2(new_n490), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(new_n294), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n500), .A2(new_n563), .A3(new_n683), .A4(new_n678), .ZN(new_n684));
  INV_X1    g498(.A(new_n412), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n414), .A2(G900), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(G902), .A3(new_n413), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n687), .A2(KEYINPUT94), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(KEYINPUT94), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n688), .A2(new_n415), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n352), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  INV_X1    g508(.A(new_n539), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n525), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT67), .B1(new_n512), .B2(new_n513), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n545), .A2(new_n544), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n299), .B1(new_n700), .B2(new_n525), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n543), .B(new_n702), .C1(new_n562), .C2(KEYINPUT32), .ZN(new_n703));
  INV_X1    g517(.A(new_n678), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n305), .B(KEYINPUT38), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n352), .A2(new_n412), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n705), .A2(new_n706), .A3(new_n492), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n690), .B(KEYINPUT39), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n500), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n190), .ZN(G45));
  OAI211_X1 g528(.A(new_n412), .B(new_n691), .C1(new_n651), .C2(new_n654), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n684), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT95), .B(G146), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G48));
  NAND2_X1  g532(.A1(new_n623), .A2(new_n630), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n637), .A2(new_n502), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n504), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n637), .A2(new_n505), .B1(new_n555), .B2(G472), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n479), .B1(new_n478), .B2(new_n299), .ZN(new_n724));
  INV_X1    g538(.A(new_n423), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n480), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(new_n726), .A3(new_n656), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT96), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n723), .A2(new_n726), .A3(KEYINPUT96), .A4(new_n656), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NAND3_X1  g547(.A1(new_n723), .A2(new_n726), .A3(new_n663), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT97), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT97), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n723), .A2(new_n726), .A3(new_n663), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  NAND2_X1  g553(.A1(new_n726), .A2(new_n683), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n563), .A2(new_n421), .A3(new_n678), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n223), .ZN(G21));
  INV_X1    g557(.A(KEYINPUT98), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n525), .B1(new_n548), .B2(new_n520), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n744), .B1(new_n745), .B2(new_n557), .ZN(new_n746));
  INV_X1    g560(.A(new_n520), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n700), .B2(KEYINPUT28), .ZN(new_n748));
  OAI211_X1 g562(.A(KEYINPUT98), .B(new_n535), .C1(new_n748), .C2(new_n525), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n541), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n502), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n628), .A2(new_n629), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n638), .A2(G472), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT99), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n502), .A2(new_n750), .B1(new_n638), .B2(G472), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT99), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n752), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n643), .A2(new_n707), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n726), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  INV_X1    g577(.A(new_n715), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n756), .A2(new_n678), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n740), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n198), .ZN(G27));
  NAND4_X1  g581(.A1(new_n303), .A2(new_n423), .A3(new_n188), .A4(new_n304), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT100), .Z(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n498), .B2(G469), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n768), .B1(new_n495), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(new_n563), .A3(new_n764), .A4(new_n631), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT42), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n715), .A2(new_n775), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n773), .A3(new_n563), .A4(new_n752), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  INV_X1    g594(.A(KEYINPUT102), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n495), .A2(new_n772), .ZN(new_n782));
  INV_X1    g596(.A(new_n768), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n563), .A2(new_n631), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT101), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n692), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n661), .A2(KEYINPUT101), .A3(new_n691), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n781), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT101), .B1(new_n661), .B2(new_n691), .ZN(new_n790));
  AND4_X1   g604(.A1(KEYINPUT101), .A2(new_n352), .A3(new_n685), .A4(new_n691), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n723), .A3(KEYINPUT102), .A4(new_n773), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  NOR2_X1   g609(.A1(new_n639), .A2(new_n704), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT106), .ZN(new_n797));
  INV_X1    g611(.A(new_n651), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n412), .B1(new_n798), .B2(new_n653), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT105), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT44), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT107), .Z(new_n808));
  NAND3_X1  g622(.A1(new_n303), .A2(new_n188), .A3(new_n304), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT104), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT45), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n479), .B1(new_n487), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n498), .A2(KEYINPUT45), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n771), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n811), .B1(new_n815), .B2(KEYINPUT46), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n816), .A2(new_n495), .ZN(new_n817));
  INV_X1    g631(.A(new_n815), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT46), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(KEYINPUT104), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT103), .B1(new_n815), .B2(KEYINPUT46), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n813), .A2(new_n814), .ZN(new_n822));
  AND4_X1   g636(.A1(KEYINPUT103), .A2(new_n822), .A3(KEYINPUT46), .A4(new_n770), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n817), .B(new_n820), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n423), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n709), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n806), .A2(KEYINPUT44), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n808), .A2(new_n810), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G137), .ZN(G39));
  INV_X1    g645(.A(KEYINPUT47), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n824), .A2(KEYINPUT47), .A3(new_n423), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n563), .A2(new_n631), .A3(new_n715), .A4(new_n809), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G140), .ZN(G42));
  NOR2_X1   g652(.A1(new_n480), .A2(new_n724), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n840), .A2(KEYINPUT49), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(KEYINPUT49), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n752), .A2(new_n425), .A3(new_n188), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n800), .A2(new_n703), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n841), .A2(new_n706), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n684), .B1(new_n692), .B2(new_n715), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n766), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n691), .A2(new_n423), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n294), .A2(new_n707), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n704), .A3(new_n703), .A4(new_n782), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT109), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT110), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  XNOR2_X1  g671(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n847), .A2(new_n852), .A3(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n731), .A2(new_n738), .A3(new_n680), .A4(new_n762), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n662), .A2(new_n655), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n642), .A3(new_n296), .A4(new_n306), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n740), .A2(new_n741), .B1(new_n863), .B2(new_n640), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n635), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n685), .A2(new_n349), .A3(new_n351), .A4(new_n691), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n868), .A2(new_n704), .A3(new_n809), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n500), .A3(new_n563), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n756), .A2(new_n773), .A3(new_n678), .A4(new_n764), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n794), .A2(new_n779), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT108), .B1(new_n867), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n794), .A2(new_n779), .A3(new_n872), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT108), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n861), .A2(new_n866), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n860), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n847), .A2(new_n852), .A3(KEYINPUT52), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(new_n847), .B2(new_n852), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n501), .A2(new_n490), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n882), .A2(new_n679), .B1(new_n729), .B2(new_n730), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n632), .B(KEYINPUT74), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n864), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n735), .A2(new_n737), .B1(new_n759), .B2(new_n761), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n873), .A2(new_n883), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n876), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n680), .A2(new_n731), .A3(new_n738), .A4(new_n762), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(KEYINPUT108), .A3(new_n885), .A4(new_n873), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n881), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n878), .B(KEYINPUT54), .C1(new_n857), .C2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n859), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n893), .A2(new_n887), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n894), .B(new_n895), .C1(new_n891), .C2(KEYINPUT53), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n892), .A2(KEYINPUT111), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT111), .B1(new_n892), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n805), .A2(new_n415), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n563), .A2(new_n752), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n726), .A2(new_n810), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n899), .A2(new_n683), .A3(new_n726), .A4(new_n759), .ZN(new_n907));
  OR2_X1    g721(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n414), .A2(G952), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n902), .A2(new_n415), .A3(new_n719), .A4(new_n703), .ZN(new_n911));
  INV_X1    g725(.A(new_n655), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n906), .A2(new_n907), .A3(new_n909), .A4(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n914), .A2(KEYINPUT116), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(KEYINPUT116), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n706), .A2(new_n492), .A3(new_n726), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n899), .A2(new_n759), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT114), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT50), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n899), .A2(new_n678), .A3(new_n756), .A4(new_n903), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n911), .A2(new_n685), .A3(new_n653), .A4(new_n798), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT50), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT51), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n839), .A2(new_n424), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n833), .A2(new_n834), .A3(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n899), .A2(new_n759), .A3(new_n810), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI22_X1  g747(.A1(new_n915), .A2(new_n916), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n930), .B(KEYINPUT112), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n833), .A2(new_n834), .A3(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n936), .A2(KEYINPUT113), .A3(new_n932), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT113), .B1(new_n936), .B2(new_n932), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n927), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n934), .B1(new_n939), .B2(KEYINPUT51), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n897), .A2(new_n898), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(G952), .A2(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n845), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT117), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT117), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n945), .B(new_n845), .C1(new_n941), .C2(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(G75));
  NOR2_X1   g761(.A1(new_n414), .A2(G952), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT120), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n286), .A2(new_n289), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(new_n287), .ZN(new_n952));
  XNOR2_X1  g766(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n894), .B1(new_n891), .B2(KEYINPUT53), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(G210), .A3(G902), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT56), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT119), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n955), .A2(new_n959), .A3(G902), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n955), .B2(G902), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n297), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n954), .A2(new_n957), .ZN(new_n964));
  AOI211_X1 g778(.A(new_n950), .B(new_n958), .C1(new_n963), .C2(new_n964), .ZN(G51));
  INV_X1    g779(.A(new_n948), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n960), .A2(new_n961), .A3(new_n822), .ZN(new_n967));
  INV_X1    g781(.A(new_n478), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n955), .A2(KEYINPUT54), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n896), .ZN(new_n970));
  XNOR2_X1  g784(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n770), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n968), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n966), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT122), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT122), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n976), .B(new_n966), .C1(new_n967), .C2(new_n973), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(G54));
  NAND3_X1  g792(.A1(new_n962), .A2(KEYINPUT58), .A3(G475), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(new_n394), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n394), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n980), .A2(new_n981), .A3(new_n948), .ZN(G60));
  INV_X1    g796(.A(KEYINPUT124), .ZN(new_n983));
  INV_X1    g797(.A(new_n649), .ZN(new_n984));
  INV_X1    g798(.A(new_n650), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(G478), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT59), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n969), .B2(new_n896), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n991), .A2(KEYINPUT123), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT123), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n993), .B(new_n990), .C1(new_n969), .C2(new_n896), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n949), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n892), .A2(new_n896), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT111), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n892), .A2(KEYINPUT111), .A3(new_n896), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n987), .B1(new_n1000), .B2(new_n989), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n983), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n991), .B(KEYINPUT123), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n989), .B1(new_n897), .B2(new_n898), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n986), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1003), .A2(new_n1005), .A3(KEYINPUT124), .A4(new_n949), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1002), .A2(new_n1006), .ZN(G63));
  NAND2_X1  g821(.A1(G217), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT60), .Z(new_n1009));
  AND2_X1   g823(.A1(new_n955), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1010), .A2(new_n676), .A3(new_n675), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1011), .B(new_n949), .C1(new_n611), .C2(new_n1010), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g827(.A(G953), .B1(new_n419), .B2(new_n218), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1014), .B1(new_n867), .B2(G953), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n951), .B1(G898), .B2(new_n414), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G69));
  OR2_X1    g831(.A1(new_n846), .A2(new_n766), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n900), .A2(new_n294), .A3(new_n707), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1018), .B1(new_n828), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n794), .A2(new_n779), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT127), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n830), .A2(new_n837), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n686), .B1(new_n1023), .B2(new_n414), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n363), .A2(new_n364), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n538), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(KEYINPUT126), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n414), .B1(G227), .B2(G900), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n713), .A2(new_n1018), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT62), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n862), .B(KEYINPUT125), .Z(new_n1033));
  INV_X1    g847(.A(new_n710), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n884), .A2(new_n1033), .A3(new_n1034), .A4(new_n810), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n830), .A2(new_n1032), .A3(new_n837), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n414), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(new_n1026), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1038), .B1(new_n1026), .B2(new_n1024), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1030), .B(new_n1039), .ZN(G72));
  OAI21_X1  g854(.A(new_n878), .B1(new_n891), .B2(new_n857), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n695), .A2(new_n525), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  NAND2_X1  g858(.A1(new_n696), .A2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g859(.A1(new_n1041), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n867), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1044), .B1(new_n1023), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(new_n1042), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n966), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1044), .B1(new_n1036), .B2(new_n1047), .ZN(new_n1051));
  AOI211_X1 g865(.A(new_n1046), .B(new_n1050), .C1(new_n697), .C2(new_n1051), .ZN(G57));
endmodule


