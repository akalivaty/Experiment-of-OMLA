//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n193), .A2(new_n189), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT24), .B(G110), .Z(new_n197));
  OAI22_X1  g011(.A1(new_n195), .A2(G110), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n199), .A2(KEYINPUT16), .A3(G140), .ZN(new_n200));
  XNOR2_X1  g014(.A(G125), .B(G140), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(KEYINPUT16), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G137), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G221), .ZN(new_n211));
  INV_X1    g025(.A(G234), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n211), .A2(new_n212), .A3(G953), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n213), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n202), .A2(G146), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n203), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT70), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n195), .A2(G110), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n196), .A2(new_n197), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n202), .A2(G146), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n221), .B(new_n222), .C1(new_n224), .C2(new_n217), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT70), .ZN(new_n226));
  AOI211_X1 g040(.A(new_n207), .B(new_n216), .C1(new_n223), .C2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n216), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n226), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n206), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n187), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT25), .ZN(new_n232));
  INV_X1    g046(.A(G217), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(G234), .B2(new_n187), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(new_n187), .C1(new_n227), .C2(new_n230), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n231), .A2(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT2), .B(G113), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(KEYINPUT66), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n245), .B2(new_n241), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  XNOR2_X1  g065(.A(G143), .B(G146), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT0), .B(G128), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n204), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n188), .A2(KEYINPUT0), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT0), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n262), .A3(KEYINPUT64), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(G137), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT11), .A3(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n267), .A2(new_n270), .A3(new_n273), .A4(new_n268), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n252), .A2(KEYINPUT0), .A3(G128), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n264), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n258), .A2(new_n188), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n256), .A2(KEYINPUT1), .A3(G146), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n255), .A3(new_n257), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n268), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n266), .A2(G137), .ZN(new_n284));
  OAI21_X1  g098(.A(G131), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n274), .A3(new_n285), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n249), .B(new_n250), .C1(new_n277), .C2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n277), .A2(new_n247), .A3(new_n248), .A4(new_n286), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n246), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT67), .ZN(new_n291));
  INV_X1    g105(.A(new_n243), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n244), .B2(new_n240), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n277), .A3(new_n286), .ZN(new_n294));
  NOR2_X1   g108(.A1(G237), .A2(G953), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G210), .ZN(new_n296));
  INV_X1    g110(.A(G101), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n299));
  XOR2_X1   g113(.A(new_n298), .B(new_n299), .Z(new_n300));
  NOR3_X1   g114(.A1(new_n252), .A2(new_n253), .A3(new_n251), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT64), .B1(new_n258), .B2(new_n262), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n276), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n272), .A2(new_n274), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n286), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n249), .ZN(new_n306));
  INV_X1    g120(.A(new_n250), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n288), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(new_n246), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n291), .A2(new_n294), .A3(new_n300), .A4(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT31), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n310), .B1(new_n309), .B2(new_n246), .ZN(new_n315));
  AOI211_X1 g129(.A(KEYINPUT67), .B(new_n293), .C1(new_n308), .C2(new_n288), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n317), .A2(KEYINPUT31), .A3(new_n294), .A4(new_n300), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n294), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n305), .A2(new_n246), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n322), .A2(new_n294), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n321), .B1(new_n323), .B2(new_n320), .ZN(new_n324));
  INV_X1    g138(.A(new_n300), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT32), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n314), .A2(new_n318), .B1(new_n324), .B2(new_n325), .ZN(new_n331));
  INV_X1    g145(.A(new_n329), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT32), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n291), .A2(new_n294), .A3(new_n325), .A4(new_n311), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n324), .A2(new_n300), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT29), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT68), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n322), .A2(new_n338), .A3(new_n294), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n338), .B2(new_n322), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n321), .B1(new_n340), .B2(new_n320), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n300), .A2(KEYINPUT29), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n187), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G472), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT69), .B(G472), .C1(new_n337), .C2(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n239), .B1(new_n334), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT9), .B(G234), .Z(new_n351));
  AOI21_X1  g165(.A(new_n211), .B1(new_n351), .B2(new_n187), .ZN(new_n352));
  INV_X1    g166(.A(G104), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT75), .B1(new_n353), .B2(G107), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(G107), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n353), .A2(KEYINPUT75), .A3(G107), .ZN(new_n357));
  OAI21_X1  g171(.A(G101), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT73), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(G104), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n353), .A2(KEYINPUT73), .A3(G107), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OR3_X1    g177(.A1(new_n353), .A2(KEYINPUT3), .A3(G107), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(new_n353), .B2(G107), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n363), .A2(new_n297), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT76), .ZN(new_n368));
  INV_X1    g182(.A(new_n282), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n367), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n282), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n275), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT12), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n304), .B1(new_n372), .B2(new_n374), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT12), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT78), .B1(new_n380), .B2(KEYINPUT12), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT77), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n358), .A2(new_n366), .A3(new_n370), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n370), .B1(new_n358), .B2(new_n366), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n368), .A2(KEYINPUT77), .A3(new_n371), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT10), .A3(new_n282), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n374), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n363), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n364), .A2(new_n365), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n395), .A2(KEYINPUT74), .A3(KEYINPUT4), .A4(new_n366), .ZN(new_n396));
  INV_X1    g210(.A(new_n276), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n254), .B2(new_n263), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT74), .A2(KEYINPUT4), .ZN(new_n399));
  OAI211_X1 g213(.A(G101), .B(new_n399), .C1(new_n394), .C2(new_n393), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n390), .A2(new_n403), .A3(new_n304), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n383), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G140), .ZN(new_n406));
  INV_X1    g220(.A(G953), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n407), .A2(G227), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n406), .B(new_n408), .Z(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n369), .B1(new_n387), .B2(new_n388), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n402), .B1(new_n412), .B2(KEYINPUT10), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n410), .B1(new_n413), .B2(new_n304), .ZN(new_n414));
  AOI211_X1 g228(.A(new_n391), .B(new_n369), .C1(new_n387), .C2(new_n388), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n275), .B1(new_n415), .B2(new_n402), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(KEYINPUT79), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT79), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n409), .B1(new_n383), .B2(new_n404), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n415), .A2(new_n275), .A3(new_n402), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n304), .B1(new_n390), .B2(new_n403), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n421), .A2(new_n422), .A3(new_n410), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n419), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G469), .ZN(new_n426));
  INV_X1    g240(.A(G469), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(new_n187), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n410), .B1(new_n421), .B2(new_n422), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n414), .A2(new_n383), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n428), .B1(new_n431), .B2(new_n427), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n352), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n434));
  NOR2_X1   g248(.A1(G475), .A2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n295), .A2(G143), .A3(G214), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(G143), .B1(new_n295), .B2(G214), .ZN(new_n439));
  OAI21_X1  g253(.A(G131), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT17), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n439), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n273), .A3(new_n437), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n442), .A2(new_n218), .A3(new_n445), .A4(new_n203), .ZN(new_n446));
  XNOR2_X1  g260(.A(G113), .B(G122), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(new_n353), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n201), .B(new_n204), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT18), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n443), .B(new_n437), .C1(new_n450), .C2(new_n273), .ZN(new_n451));
  OAI211_X1 g265(.A(KEYINPUT18), .B(G131), .C1(new_n438), .C2(new_n439), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n446), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n448), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n199), .A2(KEYINPUT19), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT19), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(G125), .A2(G140), .ZN(new_n461));
  NOR2_X1   g275(.A1(G125), .A2(G140), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT84), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n459), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(KEYINPUT84), .B2(new_n201), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n204), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n224), .B1(new_n467), .B2(KEYINPUT85), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n460), .A2(new_n463), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n201), .A2(new_n465), .A3(KEYINPUT84), .ZN(new_n470));
  AOI21_X1  g284(.A(G146), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n471), .A2(new_n472), .B1(new_n440), .B2(new_n444), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n457), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n456), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n440), .A2(new_n444), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n467), .B2(KEYINPUT85), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n203), .B1(new_n471), .B2(new_n472), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n475), .B(new_n453), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n455), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n453), .B1(new_n478), .B2(new_n479), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT86), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n456), .A3(new_n480), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(KEYINPUT87), .A3(new_n455), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n436), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT20), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n434), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n448), .B1(new_n485), .B2(KEYINPUT86), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n483), .B(new_n454), .C1(new_n492), .C2(new_n480), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT87), .B1(new_n487), .B2(new_n455), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n435), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n482), .A2(new_n490), .A3(new_n435), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n448), .B1(new_n446), .B2(new_n453), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n187), .B1(new_n454), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G475), .ZN(new_n501));
  INV_X1    g315(.A(G478), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G116), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT89), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n505), .B2(G122), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(new_n360), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT14), .ZN(new_n510));
  INV_X1    g324(.A(G122), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(G116), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G128), .B(G143), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n266), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n513), .A2(new_n266), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n509), .A2(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n508), .B(new_n360), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n510), .B(new_n507), .C1(G116), .C2(new_n511), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n508), .B(G107), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n266), .B1(new_n513), .B2(KEYINPUT13), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n256), .A2(G128), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(KEYINPUT13), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n514), .B(KEYINPUT91), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n520), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n351), .A2(G217), .A3(new_n407), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n519), .A2(new_n531), .A3(new_n527), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n504), .B1(new_n533), .B2(KEYINPUT92), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n535));
  INV_X1    g349(.A(new_n532), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n531), .B1(new_n519), .B2(new_n527), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n535), .B(new_n187), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n540), .B2(new_n503), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n498), .A2(new_n501), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G214), .B1(G237), .B2(G902), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT80), .Z(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G952), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(G953), .ZN(new_n548));
  NAND2_X1  g362(.A1(G234), .A2(G237), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT21), .B(G898), .Z(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(G902), .A3(G953), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n398), .A2(G125), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n282), .A2(new_n199), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n407), .A2(G224), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n556), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(G224), .A3(new_n407), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT5), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n244), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n192), .A2(G116), .ZN(new_n566));
  OAI21_X1  g380(.A(G113), .B1(new_n566), .B2(KEYINPUT5), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n243), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n389), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n246), .A2(new_n400), .A3(new_n396), .ZN(new_n571));
  XOR2_X1   g385(.A(G110), .B(G122), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n572), .B(KEYINPUT81), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n568), .B1(new_n388), .B2(new_n387), .ZN(new_n576));
  INV_X1    g390(.A(new_n571), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n563), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n570), .A2(new_n571), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT6), .B1(new_n580), .B2(new_n575), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n562), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT82), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n567), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n292), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT83), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n385), .A2(new_n386), .ZN(new_n590));
  OAI22_X1  g404(.A1(new_n589), .A2(new_n590), .B1(new_n373), .B2(new_n569), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n572), .B(KEYINPUT8), .Z(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n558), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n559), .A2(new_n561), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n557), .A2(new_n594), .A3(new_n558), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n593), .A2(new_n598), .A3(new_n574), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n582), .A2(new_n599), .A3(new_n187), .ZN(new_n600));
  OAI21_X1  g414(.A(G210), .B1(G237), .B2(G902), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n582), .A2(new_n599), .A3(new_n187), .A4(new_n601), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n546), .B(new_n554), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n433), .A2(new_n543), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n350), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n297), .ZN(G3));
  NAND2_X1  g422(.A1(new_n498), .A2(new_n501), .ZN(new_n609));
  OR3_X1    g423(.A1(new_n536), .A2(KEYINPUT33), .A3(new_n537), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT33), .B1(new_n536), .B2(new_n537), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(G478), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n533), .A2(new_n502), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n502), .A2(new_n187), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n609), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n603), .A2(new_n604), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n544), .A3(new_n553), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n352), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n427), .B1(new_n418), .B2(new_n424), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n429), .A2(new_n430), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n427), .A3(new_n187), .ZN(new_n625));
  INV_X1    g439(.A(new_n428), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n622), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(G472), .B1(new_n331), .B2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n327), .A2(new_n329), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n628), .A2(new_n631), .A3(new_n239), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n621), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NAND2_X1  g449(.A1(new_n489), .A2(new_n490), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n491), .A2(new_n496), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n538), .A2(new_n539), .A3(new_n504), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n534), .B2(new_n540), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n501), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n620), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND2_X1  g458(.A1(new_n229), .A2(new_n206), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n228), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n647), .B(new_n187), .C1(new_n233), .C2(G234), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n237), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n631), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n606), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G110), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT94), .B(KEYINPUT37), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  AOI22_X1  g470(.A1(new_n330), .A2(new_n333), .B1(new_n346), .B2(new_n347), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n657), .A2(new_n628), .A3(new_n650), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n637), .A2(new_n501), .A3(new_n639), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n660));
  INV_X1    g474(.A(new_n544), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n603), .B2(new_n604), .ZN(new_n662));
  OR3_X1    g476(.A1(new_n552), .A2(KEYINPUT95), .A3(G900), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT95), .B1(new_n552), .B2(G900), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n550), .A3(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n659), .A2(new_n660), .A3(new_n662), .A4(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n637), .A2(new_n639), .A3(new_n501), .A4(new_n665), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n619), .A2(new_n544), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT96), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n658), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  XOR2_X1   g485(.A(new_n665), .B(KEYINPUT39), .Z(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n433), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT40), .Z(new_n675));
  NOR2_X1   g489(.A1(new_n340), .A2(new_n300), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT97), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(KEYINPUT97), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(new_n312), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n679), .A2(KEYINPUT98), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n187), .B1(new_n679), .B2(KEYINPUT98), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n334), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT38), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n619), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n609), .A2(new_n544), .A3(new_n639), .A4(new_n650), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT99), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n675), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  INV_X1    g505(.A(new_n665), .ZN(new_n692));
  AOI211_X1 g506(.A(new_n692), .B(new_n616), .C1(new_n498), .C2(new_n501), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n658), .A2(new_n662), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NAND2_X1  g509(.A1(new_n416), .A2(new_n404), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n696), .A2(new_n410), .B1(new_n414), .B2(new_n383), .ZN(new_n697));
  OAI21_X1  g511(.A(G469), .B1(new_n697), .B2(G902), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n698), .A2(new_n625), .A3(new_n622), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n657), .A2(new_n700), .A3(new_n239), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n621), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND3_X1  g518(.A1(new_n641), .A2(new_n349), .A3(new_n699), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  AND3_X1   g520(.A1(new_n662), .A2(new_n699), .A3(new_n649), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n334), .A2(new_n348), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n553), .A4(new_n543), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  AND4_X1   g524(.A1(new_n544), .A2(new_n609), .A3(new_n619), .A4(new_n639), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n239), .A2(KEYINPUT101), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n237), .A2(new_n713), .A3(new_n238), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n341), .A2(new_n325), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n332), .B1(new_n319), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT100), .B(G472), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n331), .B2(G902), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n699), .A2(new_n715), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n711), .A2(new_n553), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n616), .B1(new_n498), .B2(new_n501), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n327), .A2(new_n187), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n717), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(new_n727), .A3(new_n665), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n662), .A2(new_n699), .A3(new_n649), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n707), .A2(new_n693), .A3(KEYINPUT102), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  NOR2_X1   g547(.A1(new_n420), .A2(new_n423), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(G469), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n352), .B1(new_n432), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n603), .A2(new_n544), .A3(new_n604), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n349), .A2(new_n693), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n725), .A2(new_n665), .A3(new_n737), .A4(new_n736), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n715), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n657), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n273), .ZN(G33));
  INV_X1    g560(.A(new_n667), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n349), .A2(new_n747), .A3(new_n736), .A4(new_n737), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  AND2_X1   g563(.A1(new_n629), .A2(new_n630), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n498), .A2(new_n617), .A3(new_n501), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT43), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n750), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT44), .A3(new_n649), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n737), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT44), .B1(new_n756), .B2(new_n649), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n418), .A2(new_n424), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n734), .A2(KEYINPUT45), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(G469), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n626), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT104), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n626), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n765), .A2(new_n770), .A3(new_n766), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n768), .A2(new_n625), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n622), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT105), .B1(new_n773), .B2(new_n672), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(new_n775), .A3(new_n622), .A4(new_n673), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n760), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  INV_X1    g592(.A(KEYINPUT47), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n772), .A2(KEYINPUT47), .A3(new_n622), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n693), .A2(new_n239), .A3(new_n657), .A4(new_n737), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  AOI21_X1  g600(.A(new_n550), .B1(new_n753), .B2(new_n755), .ZN(new_n787));
  INV_X1    g601(.A(new_n727), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n742), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n698), .A2(new_n625), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n352), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n737), .B(new_n790), .C1(new_n782), .C2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n737), .A2(new_n699), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n787), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n650), .A3(new_n788), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT113), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n239), .A2(new_n550), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n684), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n609), .A3(new_n617), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n686), .A2(new_n661), .A3(new_n699), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n801), .A2(KEYINPUT112), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(KEYINPUT112), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n790), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n790), .A2(new_n802), .A3(KEYINPUT50), .A4(new_n803), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n800), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n793), .A2(new_n797), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n657), .A2(new_n742), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n787), .A2(new_n812), .A3(new_n794), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT48), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n790), .A2(new_n662), .A3(new_n699), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n814), .A2(new_n548), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n809), .A2(new_n810), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n799), .A2(new_n618), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n637), .A2(new_n501), .A3(new_n542), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n708), .A2(new_n433), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n725), .A2(new_n727), .A3(new_n736), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n649), .A3(new_n665), .A4(new_n737), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT106), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n498), .A2(new_n501), .A3(new_n639), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n618), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n826), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n632), .B(new_n605), .C1(new_n828), .C2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n628), .A2(new_n609), .A3(new_n639), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n832), .B(new_n605), .C1(new_n349), .C2(new_n651), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n825), .A2(new_n748), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n739), .B1(new_n350), .B2(new_n740), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n741), .A2(new_n744), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n705), .A2(new_n709), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n553), .A2(new_n727), .A3(new_n699), .A4(new_n715), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n711), .A2(new_n839), .B1(new_n701), .B2(new_n621), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT107), .B1(new_n834), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n666), .A2(new_n669), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n843), .A2(new_n658), .B1(new_n730), .B2(new_n731), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n650), .A2(new_n665), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT108), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n711), .A2(new_n846), .A3(new_n683), .A4(new_n736), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n844), .A2(KEYINPUT52), .A3(new_n694), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n732), .A2(new_n670), .A3(new_n694), .A4(new_n847), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n702), .A2(new_n722), .A3(new_n705), .A4(new_n709), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n745), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT107), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n831), .A2(new_n748), .A3(new_n833), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n825), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n842), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n842), .A2(new_n857), .ZN(new_n860));
  XOR2_X1   g674(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n861));
  NAND2_X1  g675(.A1(new_n849), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n848), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n859), .B(KEYINPUT54), .C1(new_n860), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n858), .A2(new_n864), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  INV_X1    g682(.A(new_n825), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n831), .A2(new_n748), .A3(new_n833), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT110), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n239), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n433), .A2(new_n750), .A3(new_n605), .A4(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n827), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT106), .B1(new_n874), .B2(new_n725), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n875), .B2(new_n829), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n606), .B1(new_n350), .B2(new_n652), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT110), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n879), .A3(new_n748), .A4(new_n825), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n871), .A2(KEYINPUT53), .A3(new_n880), .A4(new_n854), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n848), .A2(new_n862), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n868), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n880), .A2(new_n854), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n864), .B1(new_n834), .B2(KEYINPUT110), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(KEYINPUT111), .A3(new_n863), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n867), .A2(new_n883), .A3(new_n884), .A4(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n819), .A2(new_n820), .A3(new_n866), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n547), .A2(new_n407), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n791), .B(KEYINPUT49), .Z(new_n892));
  NOR3_X1   g706(.A1(new_n892), .A2(new_n546), .A3(new_n742), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n686), .A2(new_n752), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n622), .A3(new_n684), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n895), .ZN(G75));
  NAND3_X1  g710(.A1(new_n867), .A2(new_n883), .A3(new_n887), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(G210), .A3(G902), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n579), .A2(new_n581), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n562), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT55), .Z(new_n902));
  AND3_X1   g716(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n898), .B2(new_n899), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n407), .A2(G952), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(G51));
  NAND2_X1  g720(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n888), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n428), .B(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n624), .ZN(new_n911));
  INV_X1    g725(.A(new_n764), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n897), .A2(G902), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n905), .B1(new_n911), .B2(new_n913), .ZN(G54));
  NAND2_X1  g728(.A1(KEYINPUT58), .A2(G475), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT114), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n897), .A2(G902), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n493), .A2(new_n494), .ZN(new_n918));
  OR3_X1    g732(.A1(new_n917), .A2(KEYINPUT115), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n905), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT115), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G60));
  INV_X1    g736(.A(new_n905), .ZN(new_n923));
  XNOR2_X1  g737(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n615), .B(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n866), .B2(new_n888), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n610), .A2(new_n611), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n926), .B1(new_n610), .B2(new_n611), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n908), .B2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT118), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT117), .B(KEYINPUT60), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n897), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n227), .A2(new_n230), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n647), .B(KEYINPUT119), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n897), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n923), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n938), .A2(KEYINPUT61), .A3(new_n923), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(G66));
  INV_X1    g759(.A(new_n878), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n946), .A2(new_n853), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n853), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT120), .B1(new_n949), .B2(new_n878), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n407), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n551), .A2(G224), .A3(G953), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(G898), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n900), .B1(new_n957), .B2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n956), .B(new_n958), .ZN(G69));
  NAND2_X1  g773(.A1(new_n469), .A2(new_n470), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n309), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n875), .A2(new_n829), .ZN(new_n962));
  INV_X1    g776(.A(new_n674), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(new_n349), .A3(new_n963), .A4(new_n737), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n777), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT124), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n777), .A2(new_n967), .A3(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n844), .A2(new_n970), .A3(new_n694), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n732), .A2(new_n670), .A3(new_n694), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n971), .A2(new_n973), .A3(new_n690), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n971), .A2(new_n973), .A3(KEYINPUT62), .A4(new_n690), .ZN(new_n977));
  AOI22_X1  g791(.A1(new_n976), .A2(new_n977), .B1(new_n782), .B2(new_n784), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n969), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n961), .B1(new_n979), .B2(new_n407), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n837), .A2(new_n971), .A3(new_n973), .A4(new_n748), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n711), .A2(new_n812), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n774), .B(new_n776), .C1(new_n760), .C2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n981), .A2(new_n983), .A3(new_n407), .A4(new_n785), .ZN(new_n984));
  NAND2_X1  g798(.A1(G900), .A2(G953), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n984), .A2(new_n961), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT125), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n407), .B1(G227), .B2(G900), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n980), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n988), .B1(new_n980), .B2(new_n987), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G72));
  NAND4_X1  g805(.A1(new_n951), .A2(new_n981), .A3(new_n785), .A4(new_n983), .ZN(new_n992));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n335), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n992), .A2(KEYINPUT127), .A3(new_n994), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n860), .A2(new_n865), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(KEYINPUT53), .B2(new_n858), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n325), .B1(new_n317), .B2(new_n294), .ZN(new_n1003));
  INV_X1    g817(.A(new_n994), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1003), .A2(new_n998), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n905), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n969), .A2(new_n951), .A3(new_n978), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1003), .B1(new_n1008), .B2(new_n1004), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(KEYINPUT126), .B(new_n1003), .C1(new_n1008), .C2(new_n1004), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1007), .B1(new_n1011), .B2(new_n1012), .ZN(G57));
endmodule


